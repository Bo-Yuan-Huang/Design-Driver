
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire [7:0] ACC_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] PCON_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [7:0] ie_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [6:0] \oc8051_golden_model_1.n0988 ;
  wire \oc8051_golden_model_1.n0989 ;
  wire \oc8051_golden_model_1.n0990 ;
  wire \oc8051_golden_model_1.n0991 ;
  wire \oc8051_golden_model_1.n0992 ;
  wire \oc8051_golden_model_1.n0993 ;
  wire \oc8051_golden_model_1.n0994 ;
  wire \oc8051_golden_model_1.n0995 ;
  wire \oc8051_golden_model_1.n0996 ;
  wire \oc8051_golden_model_1.n1003 ;
  wire [7:0] \oc8051_golden_model_1.n1004 ;
  wire [7:0] \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1017 ;
  wire \oc8051_golden_model_1.n1018 ;
  wire \oc8051_golden_model_1.n1019 ;
  wire \oc8051_golden_model_1.n1026 ;
  wire [7:0] \oc8051_golden_model_1.n1027 ;
  wire \oc8051_golden_model_1.n1043 ;
  wire [7:0] \oc8051_golden_model_1.n1044 ;
  wire [3:0] \oc8051_golden_model_1.n1156 ;
  wire [3:0] \oc8051_golden_model_1.n1158 ;
  wire [3:0] \oc8051_golden_model_1.n1160 ;
  wire [3:0] \oc8051_golden_model_1.n1161 ;
  wire [3:0] \oc8051_golden_model_1.n1162 ;
  wire [3:0] \oc8051_golden_model_1.n1163 ;
  wire [3:0] \oc8051_golden_model_1.n1164 ;
  wire [3:0] \oc8051_golden_model_1.n1165 ;
  wire [3:0] \oc8051_golden_model_1.n1166 ;
  wire \oc8051_golden_model_1.n1213 ;
  wire \oc8051_golden_model_1.n1258 ;
  wire [8:0] \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [7:0] \oc8051_golden_model_1.n1261 ;
  wire \oc8051_golden_model_1.n1262 ;
  wire [2:0] \oc8051_golden_model_1.n1263 ;
  wire \oc8051_golden_model_1.n1264 ;
  wire [1:0] \oc8051_golden_model_1.n1265 ;
  wire [7:0] \oc8051_golden_model_1.n1266 ;
  wire [6:0] \oc8051_golden_model_1.n1267 ;
  wire \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1270 ;
  wire \oc8051_golden_model_1.n1271 ;
  wire \oc8051_golden_model_1.n1272 ;
  wire \oc8051_golden_model_1.n1273 ;
  wire \oc8051_golden_model_1.n1274 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire \oc8051_golden_model_1.n1282 ;
  wire [7:0] \oc8051_golden_model_1.n1283 ;
  wire \oc8051_golden_model_1.n1299 ;
  wire [7:0] \oc8051_golden_model_1.n1300 ;
  wire [15:0] \oc8051_golden_model_1.n1343 ;
  wire [7:0] \oc8051_golden_model_1.n1345 ;
  wire \oc8051_golden_model_1.n1346 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1360 ;
  wire [7:0] \oc8051_golden_model_1.n1361 ;
  wire [8:0] \oc8051_golden_model_1.n1363 ;
  wire [8:0] \oc8051_golden_model_1.n1367 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [3:0] \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1370 ;
  wire [4:0] \oc8051_golden_model_1.n1374 ;
  wire \oc8051_golden_model_1.n1375 ;
  wire [8:0] \oc8051_golden_model_1.n1376 ;
  wire \oc8051_golden_model_1.n1384 ;
  wire [7:0] \oc8051_golden_model_1.n1385 ;
  wire [6:0] \oc8051_golden_model_1.n1386 ;
  wire \oc8051_golden_model_1.n1401 ;
  wire [7:0] \oc8051_golden_model_1.n1402 ;
  wire [8:0] \oc8051_golden_model_1.n1406 ;
  wire \oc8051_golden_model_1.n1407 ;
  wire [4:0] \oc8051_golden_model_1.n1412 ;
  wire \oc8051_golden_model_1.n1413 ;
  wire \oc8051_golden_model_1.n1421 ;
  wire [7:0] \oc8051_golden_model_1.n1422 ;
  wire [6:0] \oc8051_golden_model_1.n1423 ;
  wire \oc8051_golden_model_1.n1438 ;
  wire [7:0] \oc8051_golden_model_1.n1439 ;
  wire [8:0] \oc8051_golden_model_1.n1441 ;
  wire [8:0] \oc8051_golden_model_1.n1443 ;
  wire \oc8051_golden_model_1.n1444 ;
  wire [3:0] \oc8051_golden_model_1.n1445 ;
  wire [4:0] \oc8051_golden_model_1.n1446 ;
  wire [4:0] \oc8051_golden_model_1.n1448 ;
  wire \oc8051_golden_model_1.n1449 ;
  wire [8:0] \oc8051_golden_model_1.n1450 ;
  wire \oc8051_golden_model_1.n1457 ;
  wire [7:0] \oc8051_golden_model_1.n1458 ;
  wire [6:0] \oc8051_golden_model_1.n1459 ;
  wire \oc8051_golden_model_1.n1474 ;
  wire [7:0] \oc8051_golden_model_1.n1475 ;
  wire [8:0] \oc8051_golden_model_1.n1478 ;
  wire \oc8051_golden_model_1.n1479 ;
  wire \oc8051_golden_model_1.n1486 ;
  wire [7:0] \oc8051_golden_model_1.n1487 ;
  wire [6:0] \oc8051_golden_model_1.n1488 ;
  wire [7:0] \oc8051_golden_model_1.n1489 ;
  wire [8:0] \oc8051_golden_model_1.n1491 ;
  wire [8:0] \oc8051_golden_model_1.n1493 ;
  wire \oc8051_golden_model_1.n1494 ;
  wire [4:0] \oc8051_golden_model_1.n1495 ;
  wire [4:0] \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1498 ;
  wire [8:0] \oc8051_golden_model_1.n1499 ;
  wire \oc8051_golden_model_1.n1506 ;
  wire [7:0] \oc8051_golden_model_1.n1507 ;
  wire [6:0] \oc8051_golden_model_1.n1508 ;
  wire \oc8051_golden_model_1.n1523 ;
  wire [7:0] \oc8051_golden_model_1.n1524 ;
  wire [4:0] \oc8051_golden_model_1.n1526 ;
  wire \oc8051_golden_model_1.n1527 ;
  wire [7:0] \oc8051_golden_model_1.n1528 ;
  wire [6:0] \oc8051_golden_model_1.n1529 ;
  wire [7:0] \oc8051_golden_model_1.n1530 ;
  wire [8:0] \oc8051_golden_model_1.n1532 ;
  wire \oc8051_golden_model_1.n1533 ;
  wire \oc8051_golden_model_1.n1540 ;
  wire [7:0] \oc8051_golden_model_1.n1541 ;
  wire [6:0] \oc8051_golden_model_1.n1542 ;
  wire [7:0] \oc8051_golden_model_1.n1543 ;
  wire [7:0] \oc8051_golden_model_1.n1544 ;
  wire [6:0] \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [8:0] \oc8051_golden_model_1.n1549 ;
  wire [8:0] \oc8051_golden_model_1.n1550 ;
  wire [7:0] \oc8051_golden_model_1.n1551 ;
  wire [7:0] \oc8051_golden_model_1.n1552 ;
  wire [6:0] \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire \oc8051_golden_model_1.n1555 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire \oc8051_golden_model_1.n1557 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1559 ;
  wire \oc8051_golden_model_1.n1560 ;
  wire \oc8051_golden_model_1.n1561 ;
  wire \oc8051_golden_model_1.n1568 ;
  wire [7:0] \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [8:0] \oc8051_golden_model_1.n1573 ;
  wire [8:0] \oc8051_golden_model_1.n1575 ;
  wire \oc8051_golden_model_1.n1576 ;
  wire [4:0] \oc8051_golden_model_1.n1577 ;
  wire [4:0] \oc8051_golden_model_1.n1579 ;
  wire \oc8051_golden_model_1.n1580 ;
  wire \oc8051_golden_model_1.n1587 ;
  wire [7:0] \oc8051_golden_model_1.n1588 ;
  wire [6:0] \oc8051_golden_model_1.n1589 ;
  wire \oc8051_golden_model_1.n1604 ;
  wire [7:0] \oc8051_golden_model_1.n1605 ;
  wire [8:0] \oc8051_golden_model_1.n1609 ;
  wire \oc8051_golden_model_1.n1610 ;
  wire [4:0] \oc8051_golden_model_1.n1612 ;
  wire \oc8051_golden_model_1.n1613 ;
  wire \oc8051_golden_model_1.n1620 ;
  wire [7:0] \oc8051_golden_model_1.n1621 ;
  wire [6:0] \oc8051_golden_model_1.n1622 ;
  wire \oc8051_golden_model_1.n1637 ;
  wire [7:0] \oc8051_golden_model_1.n1638 ;
  wire [8:0] \oc8051_golden_model_1.n1642 ;
  wire \oc8051_golden_model_1.n1643 ;
  wire [4:0] \oc8051_golden_model_1.n1645 ;
  wire \oc8051_golden_model_1.n1646 ;
  wire \oc8051_golden_model_1.n1653 ;
  wire [7:0] \oc8051_golden_model_1.n1654 ;
  wire [6:0] \oc8051_golden_model_1.n1655 ;
  wire \oc8051_golden_model_1.n1670 ;
  wire [7:0] \oc8051_golden_model_1.n1671 ;
  wire [8:0] \oc8051_golden_model_1.n1675 ;
  wire \oc8051_golden_model_1.n1676 ;
  wire [4:0] \oc8051_golden_model_1.n1678 ;
  wire \oc8051_golden_model_1.n1679 ;
  wire \oc8051_golden_model_1.n1686 ;
  wire [7:0] \oc8051_golden_model_1.n1687 ;
  wire [6:0] \oc8051_golden_model_1.n1688 ;
  wire \oc8051_golden_model_1.n1703 ;
  wire [7:0] \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1730 ;
  wire [6:0] \oc8051_golden_model_1.n1731 ;
  wire [7:0] \oc8051_golden_model_1.n1732 ;
  wire \oc8051_golden_model_1.n1788 ;
  wire [7:0] \oc8051_golden_model_1.n1789 ;
  wire \oc8051_golden_model_1.n1805 ;
  wire [7:0] \oc8051_golden_model_1.n1806 ;
  wire \oc8051_golden_model_1.n1822 ;
  wire [7:0] \oc8051_golden_model_1.n1823 ;
  wire \oc8051_golden_model_1.n1839 ;
  wire [7:0] \oc8051_golden_model_1.n1840 ;
  wire [7:0] \oc8051_golden_model_1.n1864 ;
  wire [6:0] \oc8051_golden_model_1.n1865 ;
  wire [7:0] \oc8051_golden_model_1.n1866 ;
  wire \oc8051_golden_model_1.n1922 ;
  wire [7:0] \oc8051_golden_model_1.n1923 ;
  wire \oc8051_golden_model_1.n1939 ;
  wire [7:0] \oc8051_golden_model_1.n1940 ;
  wire \oc8051_golden_model_1.n1956 ;
  wire [7:0] \oc8051_golden_model_1.n1957 ;
  wire \oc8051_golden_model_1.n1973 ;
  wire [7:0] \oc8051_golden_model_1.n1974 ;
  wire \oc8051_golden_model_1.n2073 ;
  wire [7:0] \oc8051_golden_model_1.n2074 ;
  wire \oc8051_golden_model_1.n2090 ;
  wire [7:0] \oc8051_golden_model_1.n2091 ;
  wire \oc8051_golden_model_1.n2107 ;
  wire [7:0] \oc8051_golden_model_1.n2108 ;
  wire \oc8051_golden_model_1.n2124 ;
  wire [7:0] \oc8051_golden_model_1.n2125 ;
  wire \oc8051_golden_model_1.n2128 ;
  wire [6:0] \oc8051_golden_model_1.n2129 ;
  wire [7:0] \oc8051_golden_model_1.n2130 ;
  wire [6:0] \oc8051_golden_model_1.n2131 ;
  wire [7:0] \oc8051_golden_model_1.n2132 ;
  wire \oc8051_golden_model_1.n2147 ;
  wire [7:0] \oc8051_golden_model_1.n2148 ;
  wire \oc8051_golden_model_1.n2187 ;
  wire [7:0] \oc8051_golden_model_1.n2188 ;
  wire [6:0] \oc8051_golden_model_1.n2189 ;
  wire [7:0] \oc8051_golden_model_1.n2190 ;
  wire [3:0] \oc8051_golden_model_1.n2197 ;
  wire \oc8051_golden_model_1.n2198 ;
  wire [7:0] \oc8051_golden_model_1.n2199 ;
  wire [6:0] \oc8051_golden_model_1.n2200 ;
  wire \oc8051_golden_model_1.n2215 ;
  wire [7:0] \oc8051_golden_model_1.n2216 ;
  wire [7:0] \oc8051_golden_model_1.n2428 ;
  wire \oc8051_golden_model_1.n2431 ;
  wire \oc8051_golden_model_1.n2433 ;
  wire \oc8051_golden_model_1.n2439 ;
  wire [7:0] \oc8051_golden_model_1.n2440 ;
  wire [6:0] \oc8051_golden_model_1.n2441 ;
  wire \oc8051_golden_model_1.n2456 ;
  wire [7:0] \oc8051_golden_model_1.n2457 ;
  wire \oc8051_golden_model_1.n2461 ;
  wire \oc8051_golden_model_1.n2463 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire [6:0] \oc8051_golden_model_1.n2471 ;
  wire \oc8051_golden_model_1.n2486 ;
  wire [7:0] \oc8051_golden_model_1.n2487 ;
  wire \oc8051_golden_model_1.n2491 ;
  wire \oc8051_golden_model_1.n2493 ;
  wire \oc8051_golden_model_1.n2499 ;
  wire [7:0] \oc8051_golden_model_1.n2500 ;
  wire [6:0] \oc8051_golden_model_1.n2501 ;
  wire \oc8051_golden_model_1.n2516 ;
  wire [7:0] \oc8051_golden_model_1.n2517 ;
  wire \oc8051_golden_model_1.n2521 ;
  wire \oc8051_golden_model_1.n2523 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire [7:0] \oc8051_golden_model_1.n2530 ;
  wire [6:0] \oc8051_golden_model_1.n2531 ;
  wire \oc8051_golden_model_1.n2546 ;
  wire [7:0] \oc8051_golden_model_1.n2547 ;
  wire \oc8051_golden_model_1.n2549 ;
  wire [7:0] \oc8051_golden_model_1.n2550 ;
  wire [6:0] \oc8051_golden_model_1.n2551 ;
  wire [7:0] \oc8051_golden_model_1.n2552 ;
  wire [7:0] \oc8051_golden_model_1.n2553 ;
  wire [6:0] \oc8051_golden_model_1.n2554 ;
  wire [7:0] \oc8051_golden_model_1.n2555 ;
  wire [15:0] \oc8051_golden_model_1.n2559 ;
  wire \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [6:0] \oc8051_golden_model_1.n2567 ;
  wire \oc8051_golden_model_1.n2582 ;
  wire [7:0] \oc8051_golden_model_1.n2583 ;
  wire \oc8051_golden_model_1.n2586 ;
  wire [7:0] \oc8051_golden_model_1.n2587 ;
  wire [6:0] \oc8051_golden_model_1.n2588 ;
  wire [7:0] \oc8051_golden_model_1.n2589 ;
  wire \oc8051_golden_model_1.n2626 ;
  wire [7:0] \oc8051_golden_model_1.n2627 ;
  wire [6:0] \oc8051_golden_model_1.n2628 ;
  wire [7:0] \oc8051_golden_model_1.n2629 ;
  wire \oc8051_golden_model_1.n2634 ;
  wire [7:0] \oc8051_golden_model_1.n2635 ;
  wire [6:0] \oc8051_golden_model_1.n2636 ;
  wire [7:0] \oc8051_golden_model_1.n2637 ;
  wire \oc8051_golden_model_1.n2642 ;
  wire [7:0] \oc8051_golden_model_1.n2643 ;
  wire [6:0] \oc8051_golden_model_1.n2644 ;
  wire [7:0] \oc8051_golden_model_1.n2645 ;
  wire \oc8051_golden_model_1.n2650 ;
  wire [7:0] \oc8051_golden_model_1.n2651 ;
  wire [6:0] \oc8051_golden_model_1.n2652 ;
  wire [7:0] \oc8051_golden_model_1.n2653 ;
  wire \oc8051_golden_model_1.n2658 ;
  wire [7:0] \oc8051_golden_model_1.n2659 ;
  wire [6:0] \oc8051_golden_model_1.n2660 ;
  wire [7:0] \oc8051_golden_model_1.n2661 ;
  wire [7:0] \oc8051_golden_model_1.n2662 ;
  wire [6:0] \oc8051_golden_model_1.n2663 ;
  wire [7:0] \oc8051_golden_model_1.n2664 ;
  wire [3:0] \oc8051_golden_model_1.n2665 ;
  wire [7:0] \oc8051_golden_model_1.n2666 ;
  wire \oc8051_golden_model_1.n2667 ;
  wire \oc8051_golden_model_1.n2668 ;
  wire \oc8051_golden_model_1.n2669 ;
  wire \oc8051_golden_model_1.n2670 ;
  wire \oc8051_golden_model_1.n2671 ;
  wire \oc8051_golden_model_1.n2672 ;
  wire \oc8051_golden_model_1.n2673 ;
  wire \oc8051_golden_model_1.n2674 ;
  wire \oc8051_golden_model_1.n2681 ;
  wire [7:0] \oc8051_golden_model_1.n2682 ;
  wire [7:0] \oc8051_golden_model_1.n2702 ;
  wire [6:0] \oc8051_golden_model_1.n2703 ;
  wire [7:0] \oc8051_golden_model_1.n2719 ;
  wire \oc8051_golden_model_1.n2720 ;
  wire \oc8051_golden_model_1.n2721 ;
  wire \oc8051_golden_model_1.n2722 ;
  wire \oc8051_golden_model_1.n2723 ;
  wire \oc8051_golden_model_1.n2724 ;
  wire \oc8051_golden_model_1.n2725 ;
  wire \oc8051_golden_model_1.n2726 ;
  wire \oc8051_golden_model_1.n2727 ;
  wire \oc8051_golden_model_1.n2734 ;
  wire [7:0] \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2736 ;
  wire \oc8051_golden_model_1.n2737 ;
  wire \oc8051_golden_model_1.n2738 ;
  wire \oc8051_golden_model_1.n2739 ;
  wire \oc8051_golden_model_1.n2740 ;
  wire \oc8051_golden_model_1.n2741 ;
  wire \oc8051_golden_model_1.n2742 ;
  wire \oc8051_golden_model_1.n2743 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire [7:0] \oc8051_golden_model_1.n2751 ;
  wire [7:0] \oc8051_golden_model_1.n2784 ;
  wire [6:0] \oc8051_golden_model_1.n2785 ;
  wire [7:0] \oc8051_golden_model_1.n2786 ;
  wire \oc8051_golden_model_1.n2805 ;
  wire [7:0] \oc8051_golden_model_1.n2806 ;
  wire [6:0] \oc8051_golden_model_1.n2807 ;
  wire \oc8051_golden_model_1.n2822 ;
  wire [7:0] \oc8051_golden_model_1.n2823 ;
  wire [7:0] \oc8051_golden_model_1.n2827 ;
  wire [3:0] \oc8051_golden_model_1.n2828 ;
  wire [7:0] \oc8051_golden_model_1.n2829 ;
  wire \oc8051_golden_model_1.n2830 ;
  wire \oc8051_golden_model_1.n2831 ;
  wire \oc8051_golden_model_1.n2832 ;
  wire \oc8051_golden_model_1.n2833 ;
  wire \oc8051_golden_model_1.n2834 ;
  wire \oc8051_golden_model_1.n2835 ;
  wire \oc8051_golden_model_1.n2836 ;
  wire \oc8051_golden_model_1.n2837 ;
  wire \oc8051_golden_model_1.n2844 ;
  wire [7:0] \oc8051_golden_model_1.n2845 ;
  wire \oc8051_golden_model_1.n2863 ;
  wire [7:0] \oc8051_golden_model_1.n2864 ;
  wire \oc8051_golden_model_1.n2880 ;
  wire [7:0] \oc8051_golden_model_1.n2881 ;
  wire [7:0] \oc8051_golden_model_1.n2882 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff0 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff1 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff2 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff3 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_41654_, rst);
  not (_16087_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_16098_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_16109_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _16098_);
  and (_16120_, _16109_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_16131_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _16098_);
  and (_16142_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _16098_);
  nor (_16153_, _16142_, _16131_);
  and (_16164_, _16153_, _16120_);
  nor (_16175_, _16164_, _16087_);
  and (_16186_, _16087_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_16197_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_16208_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _16197_);
  nor (_16219_, _16208_, _16186_);
  not (_16230_, _16219_);
  and (_16241_, _16230_, _16164_);
  or (_16252_, _16241_, _16175_);
  and (_22329_, _16252_, _41654_);
  nor (_16273_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_16284_, _16273_);
  and (_16295_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_16306_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_16317_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_16328_, _16317_);
  not (_16339_, _16208_);
  nor (_16350_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_16361_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_16372_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _16361_);
  nor (_16383_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_16394_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_16405_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _16394_);
  nor (_16415_, _16405_, _16383_);
  nor (_16426_, _16415_, _16372_);
  not (_16437_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_16459_, _16372_, _16437_);
  nor (_16460_, _16459_, _16426_);
  and (_16471_, _16460_, _16350_);
  not (_16482_, _16471_);
  and (_16493_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16504_, _16493_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_16515_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16526_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _16515_);
  and (_16537_, _16526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_16548_, _16537_, _16504_);
  and (_16559_, _16548_, _16482_);
  nor (_16570_, _16559_, _16339_);
  not (_16581_, _16186_);
  nor (_16592_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_16603_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _16394_);
  nor (_16614_, _16603_, _16592_);
  nor (_16625_, _16614_, _16372_);
  not (_16636_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_16647_, _16372_, _16636_);
  nor (_16658_, _16647_, _16625_);
  and (_16669_, _16658_, _16350_);
  not (_16680_, _16669_);
  and (_16691_, _16493_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_16702_, _16526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_16713_, _16702_, _16691_);
  and (_16724_, _16713_, _16680_);
  nor (_16734_, _16724_, _16581_);
  nor (_16745_, _16734_, _16570_);
  nor (_16756_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_16767_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _16394_);
  nor (_16778_, _16767_, _16756_);
  nor (_16789_, _16778_, _16372_);
  not (_16800_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_16811_, _16372_, _16800_);
  nor (_16822_, _16811_, _16789_);
  and (_16833_, _16822_, _16350_);
  not (_16844_, _16833_);
  and (_16855_, _16493_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_16866_, _16526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_16877_, _16866_, _16855_);
  and (_16888_, _16877_, _16844_);
  nor (_16899_, _16888_, _16230_);
  nor (_16910_, _16899_, _16273_);
  and (_16921_, _16910_, _16745_);
  nor (_16932_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_16943_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _16394_);
  nor (_16954_, _16943_, _16932_);
  nor (_16965_, _16954_, _16372_);
  not (_16976_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_16987_, _16372_, _16976_);
  nor (_16998_, _16987_, _16965_);
  and (_17009_, _16998_, _16350_);
  not (_17020_, _17009_);
  and (_17031_, _16493_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_17042_, _16526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_17053_, _17042_, _17031_);
  and (_17064_, _17053_, _17020_);
  and (_17074_, _17064_, _16273_);
  nor (_17085_, _17074_, _16921_);
  not (_17096_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_17107_, _17096_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_17118_, _17107_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17129_, _17118_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_17140_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_17150_, _17140_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17161_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_17182_, _17161_, _17129_);
  not (_17183_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17204_, _17107_, _17183_);
  and (_17205_, _17204_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_17216_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17227_, _17216_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_17237_, _17227_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_17248_, _17237_, _17205_);
  and (_17259_, _17248_, _17182_);
  and (_17270_, _17140_, _17183_);
  and (_17281_, _17270_, _16998_);
  and (_17292_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_17303_, _17292_, _17183_);
  and (_17314_, _17303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_17324_, _17292_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17335_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_17346_, _17335_, _17314_);
  not (_17357_, _17346_);
  nor (_17368_, _17357_, _17281_);
  and (_17379_, _17368_, _17259_);
  not (_17390_, _17379_);
  and (_17401_, _17390_, _17085_);
  not (_17411_, _17401_);
  nor (_17422_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_17433_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _16394_);
  nor (_17444_, _17433_, _17422_);
  nor (_17455_, _17444_, _16372_);
  not (_17466_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_17477_, _16372_, _17466_);
  nor (_17488_, _17477_, _17455_);
  and (_17498_, _17488_, _16350_);
  not (_17509_, _17498_);
  and (_17520_, _16493_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_17531_, _16526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_17542_, _17531_, _17520_);
  and (_17553_, _17542_, _17509_);
  nor (_17564_, _17553_, _16339_);
  nor (_17575_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_17585_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _16394_);
  nor (_17596_, _17585_, _17575_);
  nor (_17607_, _17596_, _16372_);
  not (_17618_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_17629_, _16372_, _17618_);
  nor (_17640_, _17629_, _17607_);
  and (_17651_, _17640_, _16350_);
  not (_17662_, _17651_);
  and (_17672_, _16493_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_17683_, _16526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17694_, _17683_, _17672_);
  and (_17705_, _17694_, _17662_);
  nor (_17716_, _17705_, _16581_);
  nor (_17727_, _17716_, _17564_);
  nor (_17738_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_17749_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _16394_);
  nor (_17760_, _17749_, _17738_);
  nor (_17771_, _17760_, _16372_);
  not (_17781_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_17792_, _16372_, _17781_);
  nor (_17803_, _17792_, _17771_);
  and (_17814_, _17803_, _16350_);
  not (_17825_, _17814_);
  and (_17836_, _16493_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_17847_, _16526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_17858_, _17847_, _17836_);
  and (_17869_, _17858_, _17825_);
  nor (_17880_, _17869_, _16230_);
  nor (_17890_, _17880_, _16273_);
  and (_17901_, _17890_, _17727_);
  nor (_17912_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_17923_, _16394_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_17934_, _17923_, _17912_);
  nor (_17945_, _17934_, _16372_);
  not (_17956_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_17967_, _16372_, _17956_);
  nor (_17978_, _17967_, _17945_);
  and (_17989_, _17978_, _16350_);
  not (_18000_, _17989_);
  and (_18010_, _16493_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_18021_, _16526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_18032_, _18021_, _18010_);
  and (_18043_, _18032_, _18000_);
  and (_18054_, _18043_, _16273_);
  nor (_18065_, _18054_, _17901_);
  and (_18076_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_18087_, _17118_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_18098_, _18087_, _18076_);
  and (_18109_, _17303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_18119_, _17227_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_18130_, _18119_, _18109_);
  and (_18141_, _18130_, _18098_);
  and (_18152_, _17978_, _17270_);
  and (_18163_, _17204_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_18174_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_18185_, _18174_, _18163_);
  not (_18196_, _18185_);
  nor (_18207_, _18196_, _18152_);
  and (_18218_, _18207_, _18141_);
  not (_18228_, _18218_);
  and (_18239_, _18228_, _18065_);
  and (_18250_, _18239_, _17411_);
  not (_18261_, _18250_);
  and (_18272_, _17118_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_18283_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_18294_, _18283_, _18272_);
  and (_18305_, _17227_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_18316_, _17204_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_18327_, _18316_, _18305_);
  and (_18337_, _18327_, _18294_);
  and (_18348_, _17640_, _17270_);
  and (_18359_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_18370_, _17303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_18381_, _18370_, _18359_);
  not (_18392_, _18381_);
  nor (_18403_, _18392_, _18348_);
  and (_18414_, _18403_, _18337_);
  not (_18425_, _18414_);
  and (_18436_, _18425_, _18065_);
  and (_18446_, _17118_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_18457_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_18468_, _18457_, _18446_);
  and (_18479_, _17227_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_18490_, _17204_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_18501_, _18490_, _18479_);
  and (_18512_, _18501_, _18468_);
  and (_18523_, _17270_, _16658_);
  and (_18533_, _17303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_18544_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_18555_, _18544_, _18533_);
  not (_18566_, _18555_);
  nor (_18577_, _18566_, _18523_);
  and (_18588_, _18577_, _18512_);
  not (_18599_, _18588_);
  and (_18610_, _18599_, _17085_);
  and (_18620_, _18436_, _18610_);
  nor (_18631_, _17401_, _18620_);
  and (_18642_, _17390_, _18620_);
  nor (_18653_, _18642_, _18631_);
  and (_18664_, _18653_, _18436_);
  and (_18675_, _18239_, _17401_);
  and (_18686_, _17390_, _18065_);
  and (_18697_, _18228_, _17085_);
  nor (_18707_, _18697_, _18686_);
  nor (_18718_, _18707_, _18675_);
  and (_18729_, _18718_, _18664_);
  and (_18740_, _18718_, _18642_);
  nor (_18751_, _18740_, _18729_);
  nor (_18762_, _18751_, _18261_);
  and (_18773_, _18065_, _18599_);
  and (_18784_, _17118_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_18794_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_18805_, _18794_, _18784_);
  and (_18816_, _17227_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_18827_, _17204_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_18838_, _18827_, _18816_);
  and (_18849_, _18838_, _18805_);
  and (_18860_, _17488_, _17270_);
  and (_18871_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_18881_, _17303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_18892_, _18881_, _18871_);
  not (_18903_, _18892_);
  nor (_18914_, _18903_, _18860_);
  and (_18925_, _18914_, _18849_);
  not (_18936_, _18925_);
  and (_18947_, _18936_, _17085_);
  and (_18958_, _18947_, _18773_);
  and (_18968_, _18425_, _17085_);
  nor (_18979_, _18968_, _18773_);
  nor (_18990_, _18979_, _18620_);
  and (_19001_, _18990_, _18958_);
  nor (_19012_, _17401_, _18436_);
  nor (_19023_, _19012_, _18664_);
  and (_19034_, _19023_, _19001_);
  nor (_19045_, _18718_, _18664_);
  nor (_19055_, _19045_, _18729_);
  nor (_19066_, _19055_, _18642_);
  nor (_19077_, _19066_, _18740_);
  and (_19088_, _19077_, _19034_);
  nor (_19099_, _19077_, _19034_);
  nor (_19110_, _19099_, _19088_);
  not (_19121_, _19110_);
  and (_19132_, _17118_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_19143_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_19154_, _19143_, _19132_);
  and (_19164_, _17227_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_19175_, _17204_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_19186_, _19175_, _19164_);
  and (_19197_, _19186_, _19154_);
  and (_19208_, _17803_, _17270_);
  and (_19219_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_19230_, _17303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_19241_, _19230_, _19219_);
  not (_19252_, _19241_);
  nor (_19263_, _19252_, _19208_);
  and (_19273_, _19263_, _19197_);
  not (_19284_, _19273_);
  and (_19295_, _19284_, _18065_);
  and (_19306_, _17118_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_19317_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_19328_, _19317_, _19306_);
  and (_19339_, _17227_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_19350_, _17204_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_19361_, _19350_, _19339_);
  and (_19372_, _19361_, _19328_);
  and (_19383_, _17270_, _16460_);
  and (_19393_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and (_19404_, _17303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_19415_, _19404_, _19393_);
  not (_19426_, _19415_);
  nor (_19437_, _19426_, _19383_);
  and (_19448_, _19437_, _19372_);
  not (_19459_, _19448_);
  and (_19470_, _19459_, _17085_);
  and (_19481_, _19470_, _19295_);
  and (_19492_, _19284_, _17085_);
  not (_19502_, _19492_);
  and (_19513_, _19459_, _18065_);
  and (_19524_, _19513_, _19502_);
  and (_19535_, _19524_, _18947_);
  nor (_19546_, _19535_, _19481_);
  and (_19557_, _18936_, _18065_);
  nor (_19568_, _19557_, _18610_);
  nor (_19579_, _19568_, _18958_);
  not (_19590_, _19579_);
  nor (_19601_, _19590_, _19546_);
  nor (_19611_, _18990_, _18958_);
  nor (_19622_, _19611_, _19001_);
  and (_19633_, _19622_, _19601_);
  nor (_19644_, _19023_, _19001_);
  nor (_19655_, _19644_, _19034_);
  and (_19666_, _19655_, _19633_);
  and (_19677_, _17118_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_19688_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_19699_, _19688_, _19677_);
  and (_19710_, _17227_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_19720_, _17204_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_19731_, _19720_, _19710_);
  and (_19742_, _19731_, _19699_);
  and (_19753_, _17270_, _16822_);
  and (_19764_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_19775_, _17303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_19786_, _19775_, _19764_);
  not (_19797_, _19786_);
  nor (_19808_, _19797_, _19753_);
  and (_19819_, _19808_, _19742_);
  not (_19829_, _19819_);
  and (_19840_, _19829_, _18065_);
  and (_19851_, _19840_, _19492_);
  nor (_19862_, _19470_, _19295_);
  nor (_19873_, _19862_, _19481_);
  and (_19884_, _19873_, _19851_);
  nor (_19895_, _19524_, _18947_);
  nor (_19906_, _19895_, _19535_);
  and (_19916_, _19906_, _19884_);
  and (_19927_, _19590_, _19546_);
  nor (_19938_, _19927_, _19601_);
  and (_19949_, _19938_, _19916_);
  nor (_19960_, _19622_, _19601_);
  nor (_19971_, _19960_, _19633_);
  and (_19982_, _19971_, _19949_);
  nor (_19993_, _19655_, _19633_);
  nor (_20003_, _19993_, _19666_);
  and (_20014_, _20003_, _19982_);
  nor (_20025_, _20014_, _19666_);
  nor (_20036_, _20025_, _19121_);
  nor (_20047_, _20036_, _19088_);
  and (_20058_, _18751_, _18261_);
  nor (_20069_, _20058_, _18762_);
  not (_20080_, _20069_);
  nor (_20090_, _20080_, _20047_);
  or (_20101_, _20090_, _18675_);
  nor (_20112_, _20101_, _18762_);
  nor (_20123_, _20112_, _16328_);
  and (_20134_, _20112_, _16328_);
  nor (_20145_, _20134_, _20123_);
  not (_20156_, _20145_);
  and (_20167_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_20177_, _20080_, _20047_);
  nor (_20188_, _20177_, _20090_);
  and (_20199_, _20188_, _20167_);
  and (_20210_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_20221_, _20025_, _19121_);
  nor (_20232_, _20221_, _20036_);
  and (_20243_, _20232_, _20210_);
  nor (_20254_, _20232_, _20210_);
  nor (_20264_, _20254_, _20243_);
  not (_20275_, _20264_);
  and (_20286_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_20297_, _20003_, _19982_);
  nor (_20308_, _20297_, _20014_);
  and (_20319_, _20308_, _20286_);
  nor (_20330_, _20308_, _20286_);
  nor (_20341_, _20330_, _20319_);
  not (_20351_, _20341_);
  and (_20362_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_20373_, _19971_, _19949_);
  nor (_20384_, _20373_, _19982_);
  and (_20395_, _20384_, _20362_);
  nor (_20406_, _20384_, _20362_);
  nor (_20417_, _20406_, _20395_);
  not (_20428_, _20417_);
  and (_20438_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_20449_, _19938_, _19916_);
  nor (_20460_, _20449_, _19949_);
  and (_20471_, _20460_, _20438_);
  and (_20482_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_20493_, _19906_, _19884_);
  nor (_20504_, _20493_, _19916_);
  and (_20514_, _20504_, _20482_);
  and (_20525_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_20536_, _19873_, _19851_);
  nor (_20547_, _20536_, _19884_);
  and (_20558_, _20547_, _20525_);
  nor (_20569_, _20504_, _20482_);
  nor (_20580_, _20569_, _20514_);
  and (_20591_, _20580_, _20558_);
  nor (_20601_, _20591_, _20514_);
  not (_20612_, _20601_);
  nor (_20623_, _20460_, _20438_);
  nor (_20634_, _20623_, _20471_);
  and (_20645_, _20634_, _20612_);
  nor (_20656_, _20645_, _20471_);
  nor (_20667_, _20656_, _20428_);
  nor (_20678_, _20667_, _20395_);
  nor (_20688_, _20678_, _20351_);
  nor (_20699_, _20688_, _20319_);
  nor (_20710_, _20699_, _20275_);
  nor (_20721_, _20710_, _20243_);
  nor (_20732_, _20188_, _20167_);
  nor (_20743_, _20732_, _20199_);
  not (_20754_, _20743_);
  nor (_20765_, _20754_, _20721_);
  nor (_20775_, _20765_, _20199_);
  nor (_20786_, _20775_, _20156_);
  nor (_20797_, _20786_, _20123_);
  not (_20808_, _20797_);
  and (_20819_, _20808_, _16306_);
  and (_20830_, _20819_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_20841_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_20852_, _20841_, _20830_);
  and (_20862_, _20852_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_20873_, _20862_, _16295_);
  and (_20884_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20895_, _20884_, _20873_);
  and (_20906_, _20873_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20917_, _20906_, _20895_);
  and (_24502_, _20917_, _41654_);
  nor (_20938_, _16164_, _16197_);
  and (_20948_, _16164_, _16197_);
  or (_20959_, _20948_, _20938_);
  and (_02427_, _20959_, _41654_);
  and (_20980_, _19829_, _17085_);
  and (_02622_, _20980_, _41654_);
  nor (_21001_, _19840_, _19492_);
  nor (_21012_, _21001_, _19851_);
  and (_02816_, _21012_, _41654_);
  nor (_21032_, _20547_, _20525_);
  nor (_21043_, _21032_, _20558_);
  and (_03014_, _21043_, _41654_);
  nor (_21064_, _20580_, _20558_);
  nor (_21075_, _21064_, _20591_);
  and (_03222_, _21075_, _41654_);
  nor (_21096_, _20634_, _20612_);
  nor (_21106_, _21096_, _20645_);
  and (_03423_, _21106_, _41654_);
  and (_21127_, _20656_, _20428_);
  nor (_21138_, _21127_, _20667_);
  and (_03624_, _21138_, _41654_);
  and (_21159_, _20678_, _20351_);
  nor (_21170_, _21159_, _20688_);
  and (_03825_, _21170_, _41654_);
  and (_21190_, _20699_, _20275_);
  nor (_21201_, _21190_, _20710_);
  and (_04026_, _21201_, _41654_);
  and (_21222_, _20754_, _20721_);
  nor (_21233_, _21222_, _20765_);
  and (_04127_, _21233_, _41654_);
  and (_21254_, _20775_, _20156_);
  nor (_21265_, _21254_, _20786_);
  and (_04228_, _21265_, _41654_);
  nor (_21285_, _20808_, _16306_);
  nor (_21296_, _21285_, _20819_);
  and (_04329_, _21296_, _41654_);
  and (_21317_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_21328_, _21317_, _20819_);
  nor (_21339_, _21328_, _20830_);
  and (_04430_, _21339_, _41654_);
  nor (_21359_, _20841_, _20830_);
  nor (_21370_, _21359_, _20852_);
  and (_04531_, _21370_, _41654_);
  and (_21403_, _16284_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_21415_, _21403_, _20852_);
  nor (_21427_, _21415_, _20862_);
  and (_04632_, _21427_, _41654_);
  nor (_21449_, _20862_, _16295_);
  nor (_21450_, _21449_, _20873_);
  and (_04733_, _21450_, _41654_);
  and (_21471_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _16098_);
  nor (_21482_, _21471_, _16109_);
  not (_21493_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_21504_, _16131_, _21493_);
  and (_21515_, _21504_, _21482_);
  and (_21526_, _21515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_21536_, _21526_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21547_, _21526_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21558_, _21547_, _21536_);
  and (_00840_, _21558_, _41654_);
  and (_00866_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _41654_);
  not (_21589_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_21600_, _17869_, _21589_);
  and (_21611_, _17553_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21621_, _21611_, _21600_);
  nor (_21632_, _21621_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21643_, _17705_, _21589_);
  and (_21654_, _18043_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_21665_, _21654_, _21643_);
  and (_21676_, _21665_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21687_, _21676_, _21632_);
  nor (_21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_21708_, _21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and (_21719_, _21698_, _18218_);
  nor (_21730_, _21719_, _21708_);
  not (_21741_, _21730_);
  and (_21752_, _16888_, _21589_);
  and (_21763_, _16559_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21774_, _21763_, _21752_);
  nor (_21785_, _21774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21795_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21806_, _16724_, _21589_);
  and (_21817_, _17064_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21828_, _21817_, _21806_);
  nor (_21839_, _21828_, _21795_);
  nor (_21850_, _21839_, _21785_);
  nor (_21861_, _21850_, _21741_);
  and (_21872_, _21850_, _21741_);
  nor (_21882_, _21872_, _21861_);
  and (_21893_, _21698_, _17379_);
  nor (_21904_, _21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor (_21915_, _21904_, _21893_);
  not (_21926_, _21915_);
  nor (_21937_, _17869_, _21589_);
  nor (_21958_, _21937_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21959_, _17553_, _21589_);
  and (_21969_, _17705_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21980_, _21969_, _21959_);
  nor (_21991_, _21980_, _21795_);
  nor (_22002_, _21991_, _21958_);
  nor (_22013_, _22002_, _21926_);
  and (_22024_, _22002_, _21926_);
  nor (_22035_, _22024_, _22013_);
  not (_22046_, _22035_);
  nor (_22056_, _21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_22067_, _21698_, _18414_);
  nor (_22078_, _22067_, _22056_);
  not (_22089_, _22078_);
  nor (_22100_, _16888_, _21589_);
  nor (_22111_, _22100_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_22122_, _16559_, _21589_);
  and (_22133_, _16724_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_22143_, _22133_, _22122_);
  nor (_22154_, _22143_, _21795_);
  nor (_22165_, _22154_, _22111_);
  nor (_22176_, _22165_, _22089_);
  and (_22187_, _22165_, _22089_);
  and (_22198_, _21621_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22220_, _22198_);
  and (_22221_, _21698_, _18588_);
  nor (_22231_, _21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  nor (_22242_, _22231_, _22221_);
  and (_22253_, _22242_, _22220_);
  and (_22264_, _21774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22275_, _22264_);
  nor (_22286_, _21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  and (_22297_, _21698_, _18925_);
  nor (_22308_, _22297_, _22286_);
  and (_22318_, _22308_, _22275_);
  nor (_22330_, _22308_, _22275_);
  nor (_22341_, _22330_, _22318_);
  not (_22352_, _22341_);
  and (_22363_, _21937_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22374_, _22363_);
  and (_22385_, _21698_, _19448_);
  nor (_22396_, _21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_22406_, _22396_, _22385_);
  and (_22417_, _22406_, _22374_);
  and (_22428_, _22100_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22439_, _22428_);
  and (_22450_, _21698_, _19273_);
  nor (_22461_, _21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  nor (_22472_, _22461_, _22450_);
  nor (_22483_, _22472_, _22439_);
  not (_22493_, _22483_);
  nor (_22504_, _22406_, _22374_);
  nor (_22515_, _22504_, _22417_);
  and (_22526_, _22515_, _22493_);
  nor (_22537_, _22526_, _22417_);
  nor (_22548_, _22537_, _22352_);
  nor (_22559_, _22548_, _22318_);
  nor (_22569_, _22242_, _22220_);
  nor (_22580_, _22569_, _22253_);
  not (_22591_, _22580_);
  nor (_22602_, _22591_, _22559_);
  nor (_22613_, _22602_, _22253_);
  nor (_22624_, _22613_, _22187_);
  nor (_22635_, _22624_, _22176_);
  nor (_22646_, _22635_, _22046_);
  nor (_22657_, _22646_, _22013_);
  not (_22667_, _22657_);
  and (_22678_, _22667_, _21882_);
  or (_22689_, _22678_, _21861_);
  and (_22700_, _18043_, _17064_);
  or (_22711_, _22700_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_22722_, _21828_);
  and (_22733_, _21665_, _22722_);
  nor (_22744_, _22143_, _21980_);
  and (_22754_, _22744_, _22733_);
  or (_22765_, _22754_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_22776_, _22765_, _22711_);
  and (_22787_, _22776_, _22689_);
  and (_22798_, _22787_, _21687_);
  nor (_22809_, _22667_, _21882_);
  or (_22820_, _22809_, _22678_);
  and (_22831_, _22820_, _22798_);
  nor (_22841_, _22798_, _21730_);
  nor (_22852_, _22841_, _22831_);
  not (_22863_, _22852_);
  and (_22874_, _22852_, _21687_);
  not (_22895_, _21850_);
  nor (_22896_, _22798_, _21926_);
  and (_22907_, _22635_, _22046_);
  nor (_22928_, _22907_, _22646_);
  and (_22929_, _22928_, _22798_);
  or (_22940_, _22929_, _22896_);
  and (_22960_, _22940_, _22895_);
  nor (_22961_, _22940_, _22895_);
  nor (_22972_, _22961_, _22960_);
  not (_22993_, _22972_);
  not (_22994_, _22002_);
  nor (_23005_, _22798_, _22089_);
  nor (_23026_, _22187_, _22176_);
  nor (_23027_, _23026_, _22613_);
  and (_23038_, _23026_, _22613_);
  or (_23058_, _23038_, _23027_);
  and (_23059_, _23058_, _22798_);
  or (_23070_, _23059_, _23005_);
  and (_23091_, _23070_, _22994_);
  nor (_23092_, _23070_, _22994_);
  not (_23103_, _22165_);
  and (_23114_, _22591_, _22559_);
  or (_23125_, _23114_, _22602_);
  and (_23136_, _23125_, _22798_);
  nor (_23147_, _22798_, _22242_);
  nor (_23158_, _23147_, _23136_);
  and (_23168_, _23158_, _23103_);
  and (_23179_, _22537_, _22352_);
  nor (_23190_, _23179_, _22548_);
  not (_23201_, _23190_);
  and (_23212_, _23201_, _22798_);
  nor (_23223_, _22798_, _22308_);
  nor (_23234_, _23223_, _23212_);
  and (_23245_, _23234_, _22220_);
  nor (_23256_, _23234_, _22220_);
  nor (_23267_, _23256_, _23245_);
  not (_23278_, _23267_);
  nor (_23288_, _22515_, _22493_);
  nor (_23299_, _23288_, _22526_);
  not (_23310_, _23299_);
  and (_23321_, _23310_, _22798_);
  nor (_23332_, _22798_, _22406_);
  nor (_23343_, _23332_, _23321_);
  and (_23354_, _23343_, _22275_);
  not (_23365_, _22472_);
  and (_23376_, _22798_, _22428_);
  or (_23387_, _23376_, _23365_);
  nand (_23397_, _22798_, _22428_);
  or (_23408_, _23397_, _22472_);
  and (_23419_, _23408_, _23387_);
  nor (_23430_, _23419_, _22363_);
  and (_23441_, _23419_, _22363_);
  nor (_23452_, _23441_, _23430_);
  and (_23463_, _21698_, _19819_);
  nor (_23474_, _21698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_23485_, _23474_, _23463_);
  nor (_23496_, _23485_, _22439_);
  not (_23506_, _23496_);
  and (_23517_, _23506_, _23452_);
  nor (_23528_, _23517_, _23430_);
  nor (_23539_, _23343_, _22275_);
  nor (_23550_, _23539_, _23354_);
  not (_23561_, _23550_);
  nor (_23572_, _23561_, _23528_);
  nor (_23583_, _23572_, _23354_);
  nor (_23594_, _23583_, _23278_);
  nor (_23605_, _23594_, _23245_);
  nor (_23615_, _23158_, _23103_);
  nor (_23626_, _23615_, _23168_);
  not (_23637_, _23626_);
  nor (_23648_, _23637_, _23605_);
  nor (_23659_, _23648_, _23168_);
  nor (_23670_, _23659_, _23092_);
  nor (_23681_, _23670_, _23091_);
  nor (_23692_, _23681_, _22993_);
  or (_23703_, _23692_, _22960_);
  or (_23714_, _23703_, _22874_);
  and (_23724_, _23714_, _22776_);
  nor (_23735_, _23724_, _22863_);
  and (_23746_, _22874_, _22776_);
  and (_23757_, _23746_, _23703_);
  or (_23768_, _23757_, _23735_);
  and (_00884_, _23768_, _41654_);
  or (_23789_, _22852_, _21687_);
  and (_23800_, _23789_, _23724_);
  and (_02972_, _23800_, _41654_);
  and (_02983_, _22798_, _41654_);
  and (_03003_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _41654_);
  and (_03025_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _41654_);
  and (_03045_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _41654_);
  or (_23860_, _21515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23871_, _21526_, rst);
  and (_03056_, _23871_, _23860_);
  and (_23892_, _23800_, _22428_);
  or (_23903_, _23892_, _23485_);
  nand (_23914_, _23892_, _23485_);
  and (_23925_, _23914_, _23903_);
  and (_03066_, _23925_, _41654_);
  nor (_23945_, _23800_, _23419_);
  nor (_23956_, _23506_, _23452_);
  nor (_23967_, _23956_, _23517_);
  and (_23978_, _23967_, _23800_);
  or (_23989_, _23978_, _23945_);
  and (_03077_, _23989_, _41654_);
  and (_24010_, _23561_, _23528_);
  or (_24021_, _24010_, _23572_);
  nand (_24032_, _24021_, _23800_);
  or (_24043_, _23800_, _23343_);
  and (_24053_, _24043_, _24032_);
  and (_03088_, _24053_, _41654_);
  and (_24086_, _23583_, _23278_);
  or (_24098_, _24086_, _23594_);
  nand (_24110_, _24098_, _23800_);
  or (_24122_, _23800_, _23234_);
  and (_24134_, _24122_, _24110_);
  and (_03098_, _24134_, _41654_);
  and (_24146_, _23637_, _23605_);
  or (_24157_, _24146_, _23648_);
  nand (_24167_, _24157_, _23800_);
  or (_24178_, _23800_, _23158_);
  and (_24189_, _24178_, _24167_);
  and (_03109_, _24189_, _41654_);
  or (_24210_, _23092_, _23091_);
  and (_24221_, _24210_, _23659_);
  nor (_24232_, _24210_, _23659_);
  or (_24243_, _24232_, _24221_);
  nand (_24254_, _24243_, _23800_);
  or (_24265_, _23800_, _23070_);
  and (_24275_, _24265_, _24254_);
  and (_03120_, _24275_, _41654_);
  and (_24296_, _23681_, _22993_);
  or (_24307_, _24296_, _23692_);
  nand (_24318_, _24307_, _23800_);
  or (_24329_, _23800_, _22940_);
  and (_24340_, _24329_, _24318_);
  and (_03131_, _24340_, _41654_);
  not (_24361_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_24372_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _16098_);
  and (_24382_, _24372_, _24361_);
  and (_24393_, _24382_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24404_, _24393_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  not (_24415_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24426_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _16098_);
  and (_24437_, _24426_, _24415_);
  and (_24448_, _24437_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_24459_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24469_, _24459_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24480_, _24459_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24491_, _24480_, _24469_);
  and (_24503_, _24491_, _24448_);
  nor (_24514_, _24503_, _24404_);
  not (_24525_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_24536_, _24437_, _24525_);
  and (_24547_, _24536_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  or (_24558_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24568_, _24558_, _16098_);
  nor (_24579_, _24568_, _24372_);
  and (_24590_, _24579_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  and (_24601_, _24382_, _24415_);
  and (_24612_, _24601_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_24623_, _24612_, _24590_);
  nor (_24634_, _24623_, _24547_);
  and (_24645_, _24634_, _24514_);
  and (_24655_, _24393_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_24666_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24677_, _24666_, _24459_);
  and (_24688_, _24677_, _24448_);
  nor (_24699_, _24688_, _24655_);
  and (_24710_, _24536_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_24721_, _24579_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_24732_, _24601_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_24743_, _24732_, _24721_);
  nor (_24753_, _24743_, _24710_);
  and (_24764_, _24753_, _24699_);
  and (_24775_, _24393_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_24786_, _24579_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_24797_, _24786_, _24775_);
  not (_24808_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24819_, _24448_, _24808_);
  not (_24830_, _24819_);
  and (_24840_, _24601_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_24851_, _24536_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_24862_, _24851_, _24840_);
  and (_24873_, _24862_, _24830_);
  and (_24884_, _24873_, _24797_);
  and (_24895_, _24884_, _24764_);
  and (_24906_, _24895_, _24645_);
  and (_24917_, _24469_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_24928_, _24917_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_24938_, _24928_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_24949_, _24938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_24960_, _24949_);
  not (_24971_, _24448_);
  nor (_24992_, _24938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_24993_, _24992_, _24971_);
  and (_25004_, _24993_, _24960_);
  not (_25015_, _25004_);
  and (_25035_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_25036_, _25035_, _24426_);
  and (_25047_, _24601_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_25068_, _25047_, _25036_);
  and (_25069_, _24536_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_25080_, _24393_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_25091_, _25080_, _25069_);
  and (_25102_, _25091_, _25068_);
  and (_25122_, _25102_, _25015_);
  nor (_25123_, _24928_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_25134_, _25123_);
  nor (_25145_, _24938_, _24971_);
  and (_25156_, _25145_, _25134_);
  not (_25167_, _25156_);
  and (_25178_, _24601_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_25189_, _25178_, _25036_);
  and (_25200_, _24536_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_25210_, _24393_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_25221_, _25210_, _25200_);
  and (_25232_, _25221_, _25189_);
  and (_25253_, _25232_, _25167_);
  nor (_25254_, _25253_, _25122_);
  not (_25265_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_25276_, _24949_, _25265_);
  and (_25287_, _24949_, _25265_);
  nor (_25297_, _25287_, _25276_);
  nor (_25308_, _25297_, _24971_);
  not (_25319_, _25308_);
  and (_25330_, _24601_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_25341_, _25330_, _25036_);
  and (_25352_, _24536_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_25363_, _24393_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_25374_, _25363_, _25352_);
  and (_25385_, _25374_, _25341_);
  and (_25395_, _25385_, _25319_);
  not (_25406_, _25395_);
  and (_25427_, _24393_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_25428_, _24601_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_25439_, _25428_, _25427_);
  not (_25450_, _24917_);
  nor (_25461_, _24469_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_25472_, _25461_, _24971_);
  and (_25483_, _25472_, _25450_);
  and (_25493_, _24579_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_25504_, _24536_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_25515_, _25504_, _25493_);
  not (_25526_, _25515_);
  nor (_25537_, _25526_, _25483_);
  and (_25548_, _25537_, _25439_);
  nor (_25559_, _24917_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_25570_, _25559_, _24971_);
  nor (_25580_, _25570_, _24928_);
  and (_25591_, _24393_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_25602_, _25591_, _25580_);
  and (_25623_, _24601_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and (_25624_, _24579_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_25635_, _25624_, _25623_);
  and (_25646_, _24536_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_25657_, _25646_, _25036_);
  and (_25668_, _25657_, _25635_);
  and (_25678_, _25668_, _25602_);
  not (_25689_, _25678_);
  and (_25700_, _25689_, _25548_);
  and (_25711_, _25700_, _25406_);
  and (_25722_, _25711_, _25254_);
  nand (_25733_, _25722_, _24906_);
  and (_25744_, _23768_, _21515_);
  not (_25755_, _25744_);
  and (_25766_, _20917_, _16164_);
  not (_25777_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_25788_, _16109_, _25777_);
  and (_25799_, _25788_, _16153_);
  not (_25810_, _25799_);
  nor (_25821_, _18218_, _18043_);
  and (_25832_, _18218_, _18043_);
  nor (_25843_, _25832_, _25821_);
  not (_25854_, _17064_);
  nor (_25865_, _17379_, _25854_);
  nor (_25876_, _17379_, _17064_);
  and (_25887_, _17379_, _17064_);
  nor (_25898_, _25887_, _25876_);
  not (_25909_, _17705_);
  nor (_25920_, _18414_, _25909_);
  nor (_25931_, _18414_, _17705_);
  and (_25941_, _18414_, _17705_);
  nor (_25952_, _25941_, _25931_);
  not (_25973_, _16724_);
  and (_25974_, _18588_, _25973_);
  nor (_25985_, _25974_, _25952_);
  nor (_25996_, _25985_, _25920_);
  nor (_26007_, _25996_, _25898_);
  nor (_26018_, _26007_, _25865_);
  and (_26029_, _25996_, _25898_);
  nor (_26040_, _26029_, _26007_);
  not (_26051_, _26040_);
  and (_26062_, _25974_, _25952_);
  nor (_26083_, _26062_, _25985_);
  not (_26084_, _26083_);
  nor (_26095_, _18588_, _16724_);
  and (_26106_, _18588_, _16724_);
  nor (_26117_, _26106_, _26095_);
  not (_26128_, _26117_);
  and (_26139_, _18925_, _17553_);
  nor (_26150_, _18925_, _17553_);
  nor (_26161_, _26150_, _26139_);
  nor (_26172_, _19448_, _16559_);
  and (_26183_, _19448_, _16559_);
  nor (_26194_, _26183_, _26172_);
  nor (_26205_, _19273_, _17869_);
  and (_26216_, _19273_, _17869_);
  nor (_26227_, _26216_, _26205_);
  not (_26238_, _16888_);
  and (_26249_, _19819_, _26238_);
  nor (_26260_, _26249_, _26227_);
  not (_26271_, _17869_);
  nor (_26282_, _19273_, _26271_);
  nor (_26293_, _26282_, _26260_);
  nor (_26304_, _26293_, _26194_);
  not (_26315_, _16559_);
  nor (_26326_, _19448_, _26315_);
  nor (_26337_, _26326_, _26304_);
  nor (_26347_, _26337_, _26161_);
  and (_26358_, _26337_, _26161_);
  nor (_26369_, _26358_, _26347_);
  not (_26380_, _26369_);
  and (_26391_, _26293_, _26194_);
  nor (_26402_, _26391_, _26304_);
  not (_26413_, _26402_);
  and (_26424_, _26249_, _26227_);
  nor (_26435_, _26424_, _26260_);
  not (_26446_, _26435_);
  nor (_26457_, _19819_, _16888_);
  and (_26468_, _19819_, _16888_);
  nor (_26479_, _26468_, _26457_);
  not (_26490_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_26501_, _16372_, _26490_);
  not (_26512_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26533_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26534_, _26533_, _17934_);
  nor (_26545_, _26534_, _26512_);
  nor (_26556_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26567_, _26556_, _16614_);
  not (_26578_, _26567_);
  not (_26589_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_26600_, _26589_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26611_, _26600_, _16954_);
  not (_26622_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26633_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _26622_);
  and (_26644_, _26633_, _17596_);
  nor (_26655_, _26644_, _26611_);
  and (_26666_, _26655_, _26578_);
  and (_26677_, _26666_, _26545_);
  and (_26688_, _26533_, _17444_);
  nor (_26699_, _26688_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26709_, _26633_, _17760_);
  not (_26720_, _26709_);
  and (_26731_, _26600_, _16415_);
  and (_26742_, _26556_, _16778_);
  nor (_26753_, _26742_, _26731_);
  and (_26764_, _26753_, _26720_);
  and (_26775_, _26764_, _26699_);
  nor (_26786_, _26775_, _26677_);
  nor (_26797_, _26786_, _16372_);
  nor (_26808_, _26797_, _26501_);
  and (_26829_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_26830_, _26829_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_26841_, _26830_);
  and (_26852_, _26841_, _26808_);
  and (_26863_, _26841_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_26874_, _26863_, _26852_);
  nor (_26885_, _26874_, _26479_);
  and (_26896_, _26885_, _26446_);
  and (_26907_, _26896_, _26413_);
  and (_26918_, _26907_, _26380_);
  not (_26939_, _17553_);
  or (_26940_, _18925_, _26939_);
  and (_26951_, _18925_, _26939_);
  or (_26962_, _26337_, _26951_);
  and (_26973_, _26962_, _26940_);
  or (_26984_, _26973_, _26918_);
  and (_26995_, _26984_, _26128_);
  and (_27006_, _26995_, _26084_);
  and (_27017_, _27006_, _26051_);
  nor (_27028_, _27017_, _26018_);
  nor (_27039_, _27028_, _25843_);
  and (_27050_, _27028_, _25843_);
  nor (_27060_, _27050_, _27039_);
  nor (_27071_, _27060_, _25810_);
  not (_27082_, _27071_);
  not (_27093_, _25843_);
  not (_27104_, _25898_);
  and (_27115_, _26095_, _25952_);
  nor (_27126_, _27115_, _25931_);
  nor (_27137_, _27126_, _27104_);
  not (_27158_, _26194_);
  and (_27159_, _26457_, _26227_);
  nor (_27170_, _27159_, _26205_);
  nor (_27181_, _27170_, _27158_);
  nor (_27192_, _27181_, _26172_);
  nor (_27203_, _27192_, _26161_);
  and (_27214_, _27192_, _26161_);
  nor (_27225_, _27214_, _27203_);
  not (_27236_, _26479_);
  nor (_27247_, _26874_, _27236_);
  and (_27258_, _27247_, _26227_);
  and (_27269_, _27170_, _27158_);
  nor (_27280_, _27269_, _27181_);
  and (_27291_, _27280_, _27258_);
  not (_27302_, _27291_);
  nor (_27313_, _27302_, _27225_);
  nor (_27324_, _27192_, _26139_);
  or (_27335_, _27324_, _26150_);
  or (_27346_, _27335_, _27313_);
  and (_27357_, _27346_, _26117_);
  and (_27368_, _27357_, _25952_);
  and (_27379_, _27126_, _27104_);
  nor (_27390_, _27379_, _27137_);
  and (_27401_, _27390_, _27368_);
  or (_27421_, _27401_, _27137_);
  nor (_27422_, _27421_, _25876_);
  and (_27433_, _27422_, _27093_);
  nor (_27444_, _27422_, _27093_);
  not (_27455_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_27466_, _21471_, _27455_);
  and (_27477_, _27466_, _16153_);
  not (_27488_, _27477_);
  or (_27499_, _27488_, _27444_);
  nor (_27510_, _27499_, _27433_);
  and (_27521_, _16142_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27532_, _27521_, _25788_);
  nor (_27543_, _19819_, _19273_);
  and (_27554_, _27543_, _19459_);
  and (_27565_, _27554_, _18936_);
  and (_27576_, _27565_, _18599_);
  and (_27587_, _27576_, _18425_);
  and (_27598_, _27587_, _17390_);
  and (_27609_, _27598_, _26874_);
  not (_27620_, _26874_);
  and (_27631_, _17379_, _18414_);
  and (_27642_, _19819_, _19273_);
  and (_27653_, _27642_, _19448_);
  and (_27664_, _27653_, _18925_);
  and (_27675_, _27664_, _18588_);
  and (_27686_, _27675_, _27631_);
  and (_27707_, _27686_, _27620_);
  nor (_27708_, _27707_, _27609_);
  and (_27719_, _27708_, _18218_);
  nor (_27730_, _27708_, _18218_);
  nor (_27741_, _27730_, _27719_);
  and (_27752_, _27741_, _27532_);
  not (_27763_, _18043_);
  nor (_27773_, _26874_, _27763_);
  not (_27784_, _27773_);
  and (_27795_, _26874_, _18218_);
  and (_27806_, _27521_, _16120_);
  not (_27817_, _27806_);
  nor (_27828_, _27817_, _27795_);
  and (_27839_, _27828_, _27784_);
  nor (_27850_, _27839_, _27752_);
  and (_27861_, _27466_, _21504_);
  and (_27872_, _19448_, _19273_);
  nor (_27883_, _27872_, _18925_);
  and (_27894_, _27883_, _27861_);
  and (_27905_, _27894_, _18599_);
  nor (_27916_, _27905_, _18425_);
  and (_27927_, _27916_, _17379_);
  nor (_27938_, _27631_, _18218_);
  nor (_27949_, _27938_, _27894_);
  and (_27960_, _27949_, _26874_);
  nor (_27971_, _27960_, _27927_);
  nor (_27982_, _27971_, _18228_);
  and (_27993_, _27971_, _18228_);
  nor (_28004_, _27993_, _27982_);
  and (_28015_, _28004_, _27861_);
  and (_28026_, _27521_, _27466_);
  not (_28037_, _28026_);
  nor (_28048_, _28037_, _26874_);
  not (_28059_, _28048_);
  not (_28070_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_28081_, _16142_, _28070_);
  and (_28092_, _28081_, _27466_);
  not (_28103_, _28092_);
  nor (_28114_, _28103_, _25832_);
  and (_28124_, _28081_, _21482_);
  and (_28145_, _28124_, _25843_);
  nor (_28146_, _28145_, _28114_);
  and (_28157_, _21504_, _16120_);
  and (_28168_, _28157_, _25821_);
  and (_28179_, _25788_, _21504_);
  and (_28190_, _28179_, _18218_);
  nor (_28201_, _28190_, _28168_);
  and (_28212_, _21482_, _16153_);
  not (_28223_, _28212_);
  nor (_28234_, _28223_, _18218_);
  not (_28245_, _28234_);
  and (_28256_, _27521_, _21482_);
  not (_28267_, _28256_);
  nor (_28278_, _28267_, _19819_);
  and (_28289_, _28081_, _16109_);
  not (_28300_, _28289_);
  nor (_28311_, _28300_, _17379_);
  nor (_28332_, _28311_, _28278_);
  and (_28333_, _28332_, _28245_);
  and (_28344_, _28333_, _28201_);
  and (_28355_, _28344_, _28146_);
  and (_28366_, _28355_, _28059_);
  not (_28377_, _28366_);
  nor (_28388_, _28377_, _28015_);
  and (_28399_, _28388_, _27850_);
  not (_28410_, _28399_);
  nor (_28421_, _28410_, _27510_);
  and (_28432_, _28421_, _27082_);
  not (_28443_, _28432_);
  nor (_28454_, _28443_, _25766_);
  and (_28465_, _28454_, _25755_);
  not (_28475_, _28465_);
  or (_28486_, _28475_, _25733_);
  not (_28497_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_28508_, \oc8051_top_1.oc8051_decoder1.wr , _16098_);
  not (_28519_, _28508_);
  nor (_28530_, _28519_, _24437_);
  and (_28541_, _28530_, _28497_);
  not (_28552_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_28563_, _25733_, _28552_);
  and (_28574_, _28563_, _28541_);
  and (_28585_, _28574_, _28486_);
  nor (_28596_, _28530_, _28552_);
  nor (_28607_, _27444_, _25821_);
  nor (_28618_, _28607_, _27488_);
  not (_28629_, _28618_);
  and (_28640_, _18218_, _27763_);
  nor (_28651_, _28640_, _27039_);
  nor (_28662_, _28651_, _25810_);
  and (_28673_, _28081_, _16120_);
  not (_28684_, _28673_);
  nor (_28695_, _28684_, _18218_);
  not (_28706_, _28695_);
  or (_28717_, _28223_, _26874_);
  nor (_28728_, _28037_, _19819_);
  nor (_28739_, _28728_, _27894_);
  and (_28750_, _28739_, _28717_);
  and (_28761_, _28750_, _28706_);
  nor (_28772_, _26863_, _26808_);
  not (_28783_, _28124_);
  nor (_28793_, _28783_, _26852_);
  nor (_28804_, _28793_, _28092_);
  or (_28815_, _28804_, _28772_);
  and (_28826_, _26874_, _17379_);
  and (_28837_, _28826_, _27916_);
  nor (_28848_, _28837_, _27795_);
  not (_28869_, _27861_);
  nor (_28870_, _26874_, _18218_);
  not (_28881_, _28870_);
  nor (_28892_, _28881_, _27927_);
  nor (_28903_, _28892_, _28869_);
  and (_28914_, _28903_, _28848_);
  and (_28925_, _26830_, _26808_);
  and (_28936_, _28081_, _25788_);
  and (_28947_, _28157_, _26808_);
  nor (_28958_, _28947_, _28936_);
  nor (_28969_, _28958_, _28925_);
  nor (_28980_, _28267_, _26808_);
  and (_28991_, _28980_, _27620_);
  and (_29002_, _28179_, _26874_);
  or (_29013_, _29002_, _28991_);
  or (_29024_, _29013_, _28969_);
  nor (_29035_, _29024_, _28914_);
  and (_29046_, _29035_, _28815_);
  and (_29057_, _29046_, _28761_);
  not (_29068_, _29057_);
  nor (_29079_, _29068_, _28662_);
  and (_29090_, _29079_, _28629_);
  not (_29101_, _24645_);
  nor (_29112_, _24884_, _24764_);
  and (_29122_, _29112_, _29101_);
  and (_29133_, _29122_, _25722_);
  nand (_29144_, _29133_, _29090_);
  or (_29155_, _29133_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_29166_, _28530_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_29177_, _29166_, _29155_);
  and (_29188_, _29177_, _29144_);
  or (_29199_, _29188_, _28596_);
  or (_29210_, _29199_, _28585_);
  and (_06649_, _29210_, _41654_);
  and (_29231_, _23925_, _21515_);
  not (_29242_, _29231_);
  and (_29253_, _21233_, _16164_);
  nor (_29264_, _28783_, _26457_);
  nor (_29275_, _29264_, _28092_);
  or (_29286_, _29275_, _26468_);
  and (_29297_, _27521_, _27455_);
  not (_29308_, _29297_);
  nor (_29319_, _29308_, _19273_);
  and (_29330_, _28936_, _18228_);
  nor (_29341_, _29330_, _29319_);
  and (_29352_, _29341_, _29286_);
  nor (_29363_, _28684_, _26874_);
  nor (_29374_, _27817_, _16888_);
  and (_29385_, _27532_, _19819_);
  nor (_29396_, _29385_, _29374_);
  nor (_29417_, _28212_, _27861_);
  nor (_29418_, _29417_, _19819_);
  not (_29429_, _29418_);
  nand (_29439_, _29429_, _29396_);
  nor (_29450_, _29439_, _29363_);
  and (_29461_, _29450_, _29352_);
  and (_29472_, _26874_, _27236_);
  nor (_29483_, _29472_, _27247_);
  not (_29494_, _29483_);
  nor (_29505_, _27477_, _25799_);
  nor (_29516_, _29505_, _29494_);
  not (_29527_, _29516_);
  and (_29538_, _28157_, _26457_);
  and (_29549_, _28179_, _19819_);
  nor (_29560_, _29549_, _29538_);
  and (_29571_, _29560_, _29527_);
  and (_29582_, _29571_, _29461_);
  not (_29593_, _29582_);
  nor (_29604_, _29593_, _29253_);
  and (_29615_, _29604_, _29242_);
  not (_29626_, _29615_);
  or (_29637_, _29626_, _25733_);
  not (_29648_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_29659_, _25733_, _29648_);
  and (_29680_, _29659_, _28541_);
  and (_29681_, _29680_, _29637_);
  nor (_29692_, _28530_, _29648_);
  not (_29703_, _29090_);
  or (_29714_, _29703_, _25733_);
  and (_29725_, _29659_, _29166_);
  and (_29736_, _29725_, _29714_);
  or (_29746_, _29736_, _29692_);
  or (_29757_, _29746_, _29681_);
  and (_08887_, _29757_, _41654_);
  and (_29778_, _21265_, _16164_);
  not (_29789_, _29778_);
  and (_29800_, _23989_, _21515_);
  nor (_29811_, _27817_, _17869_);
  nor (_29822_, _27642_, _27543_);
  not (_29833_, _29822_);
  nor (_29844_, _29833_, _26874_);
  and (_29855_, _29833_, _26874_);
  nor (_29866_, _29855_, _29844_);
  and (_29877_, _29866_, _27532_);
  nor (_29888_, _29877_, _29811_);
  nor (_29899_, _27883_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_29910_, _29899_, _19284_);
  nor (_29921_, _29899_, _19284_);
  nor (_29932_, _29921_, _29910_);
  nor (_29943_, _29932_, _28869_);
  not (_29954_, _29943_);
  nor (_29965_, _28223_, _19273_);
  not (_29986_, _29965_);
  nor (_29987_, _29308_, _19448_);
  nor (_29998_, _28300_, _19819_);
  nor (_30009_, _29998_, _29987_);
  and (_30020_, _30009_, _29986_);
  and (_30031_, _28124_, _26227_);
  nor (_30042_, _28103_, _26216_);
  not (_30053_, _30042_);
  and (_30063_, _28157_, _26205_);
  and (_30074_, _28179_, _19273_);
  nor (_30085_, _30074_, _30063_);
  nand (_30096_, _30085_, _30053_);
  nor (_30107_, _30096_, _30031_);
  and (_30118_, _30107_, _30020_);
  and (_30129_, _30118_, _29954_);
  nor (_30140_, _26457_, _26227_);
  or (_30151_, _30140_, _27159_);
  and (_30162_, _30151_, _27247_);
  nor (_30173_, _30151_, _27247_);
  or (_30184_, _30173_, _30162_);
  and (_30195_, _30184_, _27477_);
  nor (_30206_, _26885_, _26446_);
  nor (_30217_, _30206_, _26896_);
  nor (_30228_, _30217_, _25810_);
  nor (_30239_, _30228_, _30195_);
  and (_30250_, _30239_, _30129_);
  and (_30261_, _30250_, _29888_);
  not (_30272_, _30261_);
  nor (_30283_, _30272_, _29800_);
  and (_30294_, _30283_, _29789_);
  not (_30315_, _30294_);
  or (_30316_, _30315_, _25733_);
  not (_30327_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_30338_, _25733_, _30327_);
  and (_30349_, _30338_, _28541_);
  and (_30359_, _30349_, _30316_);
  nor (_30370_, _28530_, _30327_);
  nand (_30382_, _25722_, _24645_);
  not (_30403_, _24884_);
  and (_30414_, _30403_, _24764_);
  not (_30425_, _30414_);
  nor (_30436_, _30425_, _30382_);
  nand (_30447_, _30436_, _29090_);
  or (_30458_, _30436_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_30469_, _30458_, _29166_);
  and (_30480_, _30469_, _30447_);
  or (_30491_, _30480_, _30370_);
  or (_30502_, _30491_, _30359_);
  and (_08898_, _30502_, _41654_);
  and (_30523_, _24053_, _21515_);
  not (_30534_, _30523_);
  and (_30545_, _21296_, _16164_);
  nor (_30556_, _27817_, _16559_);
  and (_30567_, _27642_, _27620_);
  and (_30578_, _27543_, _26874_);
  nor (_30589_, _30578_, _30567_);
  nor (_30600_, _30589_, _19448_);
  not (_30611_, _27532_);
  and (_30622_, _30589_, _19448_);
  or (_30633_, _30622_, _30611_);
  nor (_30644_, _30633_, _30600_);
  nor (_30655_, _30644_, _30556_);
  nor (_30666_, _26896_, _26413_);
  nor (_30676_, _30666_, _26907_);
  nor (_30687_, _30676_, _25810_);
  nor (_30698_, _29308_, _18925_);
  and (_30709_, _28157_, _26172_);
  and (_30720_, _28179_, _19448_);
  nor (_30731_, _30720_, _30709_);
  nor (_30742_, _28103_, _26183_);
  and (_30753_, _28124_, _26194_);
  nor (_30764_, _30753_, _30742_);
  nor (_30775_, _28300_, _19273_);
  nor (_30786_, _28223_, _19448_);
  nor (_30807_, _30786_, _30775_);
  and (_30808_, _30807_, _30764_);
  nand (_30818_, _30808_, _30731_);
  nor (_30829_, _30818_, _30698_);
  not (_30840_, _30829_);
  nor (_30851_, _30840_, _30687_);
  nor (_30862_, _27280_, _27258_);
  nor (_30873_, _30862_, _27488_);
  and (_30884_, _30873_, _27302_);
  nor (_30895_, _29921_, _19448_);
  and (_30906_, _27872_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_30917_, _30906_, _30895_);
  nor (_30928_, _30917_, _28869_);
  nor (_30939_, _30928_, _30884_);
  and (_30950_, _30939_, _30851_);
  and (_30960_, _30950_, _30655_);
  not (_30971_, _30960_);
  nor (_30982_, _30971_, _30545_);
  and (_30993_, _30982_, _30534_);
  not (_31004_, _30993_);
  or (_31015_, _31004_, _25733_);
  not (_31036_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_31037_, _25733_, _31036_);
  and (_31048_, _31037_, _28541_);
  and (_31059_, _31048_, _31015_);
  nor (_31070_, _28530_, _31036_);
  or (_31081_, _29112_, _30382_);
  and (_31092_, _31081_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_31103_, _24764_);
  and (_31113_, _24645_, _24884_);
  and (_31124_, _31113_, _31103_);
  not (_31135_, _31124_);
  nor (_31146_, _31135_, _29090_);
  and (_31157_, _24645_, _24764_);
  and (_31168_, _31157_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_31179_, _31168_, _31146_);
  and (_31190_, _31179_, _25722_);
  or (_31201_, _31190_, _31092_);
  and (_31212_, _31201_, _29166_);
  or (_31223_, _31212_, _31070_);
  or (_31234_, _31223_, _31059_);
  and (_08908_, _31234_, _41654_);
  and (_31254_, _21339_, _16164_);
  not (_31265_, _31254_);
  and (_31276_, _24134_, _21515_);
  nor (_31287_, _26907_, _26380_);
  nor (_31298_, _31287_, _26918_);
  nor (_31309_, _31298_, _25810_);
  not (_31320_, _31309_);
  and (_31331_, _28157_, _26150_);
  and (_31342_, _28179_, _18925_);
  nor (_31353_, _31342_, _31331_);
  nor (_31364_, _29308_, _18588_);
  nor (_31375_, _28300_, _19448_);
  nor (_31386_, _28223_, _18925_);
  or (_31397_, _31386_, _31375_);
  nor (_31407_, _31397_, _31364_);
  and (_31418_, _31407_, _31353_);
  and (_31429_, _27302_, _27225_);
  or (_31440_, _31429_, _27488_);
  nor (_31451_, _31440_, _27313_);
  nor (_31462_, _27817_, _17553_);
  and (_31473_, _27554_, _26874_);
  and (_31484_, _27653_, _27620_);
  nor (_31495_, _31484_, _31473_);
  nor (_31506_, _31495_, _18925_);
  and (_31517_, _31495_, _18925_);
  or (_31528_, _31517_, _30611_);
  nor (_31539_, _31528_, _31506_);
  nor (_31550_, _31539_, _31462_);
  nor (_31560_, _28103_, _26139_);
  and (_31571_, _28124_, _26161_);
  nor (_31582_, _31571_, _31560_);
  not (_31593_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_31614_, _27872_, _31593_);
  nor (_31615_, _31614_, _18936_);
  or (_31626_, _31615_, _28869_);
  or (_31637_, _31626_, _27883_);
  and (_31648_, _31637_, _31582_);
  nand (_31659_, _31648_, _31550_);
  nor (_31670_, _31659_, _31451_);
  and (_31681_, _31670_, _31418_);
  and (_31692_, _31681_, _31320_);
  not (_31703_, _31692_);
  nor (_31713_, _31703_, _31276_);
  and (_31724_, _31713_, _31265_);
  not (_31735_, _31724_);
  or (_31746_, _31735_, _25733_);
  not (_31757_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_31768_, _25733_, _31757_);
  and (_31779_, _31768_, _28541_);
  and (_31790_, _31779_, _31746_);
  nor (_31801_, _28530_, _31757_);
  and (_31812_, _30382_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_31822_, _29112_, _24645_);
  not (_31833_, _31822_);
  nor (_31844_, _31833_, _29090_);
  nor (_31855_, _31157_, _31113_);
  nor (_31866_, _31855_, _31757_);
  or (_31877_, _31866_, _31844_);
  and (_31888_, _31877_, _25722_);
  or (_31899_, _31888_, _31812_);
  and (_31910_, _31899_, _29166_);
  or (_31921_, _31910_, _31801_);
  or (_31931_, _31921_, _31790_);
  and (_08919_, _31931_, _41654_);
  and (_31952_, _24189_, _21515_);
  not (_31963_, _31952_);
  and (_31974_, _21370_, _16164_);
  nor (_31985_, _26984_, _26117_);
  and (_31996_, _26984_, _26117_);
  nor (_32007_, _31996_, _31985_);
  and (_32018_, _32007_, _25799_);
  not (_32029_, _32018_);
  nor (_32039_, _27346_, _26117_);
  not (_32050_, _32039_);
  nor (_32061_, _27488_, _27357_);
  and (_32072_, _32061_, _32050_);
  nor (_32083_, _26874_, _16724_);
  and (_32094_, _26874_, _18599_);
  nor (_32105_, _32094_, _32083_);
  nor (_32116_, _32105_, _27817_);
  and (_32127_, _27565_, _26874_);
  and (_32138_, _27664_, _27620_);
  nor (_32148_, _32138_, _32127_);
  and (_32159_, _32148_, _18588_);
  nor (_32170_, _32148_, _18588_);
  nor (_32181_, _32170_, _32159_);
  and (_32192_, _32181_, _27532_);
  nor (_32203_, _32192_, _32116_);
  nor (_32214_, _27894_, _18599_);
  not (_32225_, _32214_);
  nor (_32246_, _27905_, _28869_);
  and (_32247_, _32246_, _32225_);
  not (_32257_, _32247_);
  and (_32268_, _28124_, _26117_);
  and (_32279_, _28157_, _26095_);
  nor (_32290_, _28103_, _26106_);
  and (_32301_, _28179_, _18588_);
  or (_32312_, _32301_, _32290_);
  or (_32323_, _32312_, _32279_);
  nor (_32334_, _32323_, _32268_);
  nor (_32345_, _28223_, _18588_);
  nor (_32356_, _28300_, _18925_);
  nor (_32366_, _29308_, _18414_);
  or (_32377_, _32366_, _32356_);
  nor (_32388_, _32377_, _32345_);
  and (_32399_, _32388_, _32334_);
  and (_32410_, _32399_, _32257_);
  and (_32421_, _32410_, _32203_);
  not (_32432_, _32421_);
  nor (_32443_, _32432_, _32072_);
  and (_32454_, _32443_, _32029_);
  not (_32465_, _32454_);
  nor (_32475_, _32465_, _31974_);
  and (_32486_, _32475_, _31963_);
  not (_32497_, _32486_);
  or (_32508_, _32497_, _25733_);
  not (_32519_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_32530_, _25733_, _32519_);
  and (_32551_, _32530_, _28541_);
  and (_32552_, _32551_, _32508_);
  nor (_32563_, _28530_, _32519_);
  not (_32574_, _25722_);
  and (_32584_, _24895_, _29101_);
  nor (_32595_, _24895_, _29101_);
  nor (_32606_, _32595_, _32584_);
  or (_32617_, _32606_, _32574_);
  and (_32628_, _32617_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_32639_, _32584_, _29703_);
  and (_32650_, _32595_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_32661_, _32650_, _32639_);
  and (_32672_, _32661_, _25722_);
  or (_32683_, _32672_, _32628_);
  and (_32693_, _32683_, _29166_);
  or (_32704_, _32693_, _32563_);
  or (_32715_, _32704_, _32552_);
  and (_08930_, _32715_, _41654_);
  and (_32736_, _24275_, _21515_);
  not (_32747_, _32736_);
  and (_32758_, _21427_, _16164_);
  nor (_32769_, _26095_, _25952_);
  nor (_32780_, _32769_, _27115_);
  nor (_32791_, _32780_, _27357_);
  nor (_32801_, _32791_, _27368_);
  and (_32812_, _32801_, _27477_);
  not (_32823_, _32812_);
  nor (_32834_, _26995_, _26084_);
  nor (_32845_, _32834_, _27006_);
  nor (_32856_, _32845_, _25810_);
  nor (_32867_, _26874_, _17705_);
  and (_32878_, _26874_, _18425_);
  nor (_32899_, _32878_, _32867_);
  nor (_32900_, _32899_, _27817_);
  and (_32910_, _27576_, _26874_);
  and (_32921_, _27675_, _27620_);
  nor (_32932_, _32921_, _32910_);
  and (_32943_, _32932_, _18414_);
  nor (_32954_, _32932_, _18414_);
  or (_32965_, _32954_, _30611_);
  nor (_32976_, _32965_, _32943_);
  nor (_32987_, _32976_, _32900_);
  nor (_32998_, _27960_, _27905_);
  and (_33009_, _32998_, _18414_);
  nor (_33019_, _32998_, _18414_);
  nor (_33030_, _33019_, _33009_);
  nor (_33041_, _33030_, _28869_);
  and (_33052_, _28124_, _25952_);
  not (_33063_, _33052_);
  nor (_33074_, _28103_, _25941_);
  not (_33085_, _33074_);
  and (_33096_, _28157_, _25931_);
  and (_33107_, _28179_, _18414_);
  nor (_33118_, _33107_, _33096_);
  and (_33128_, _33118_, _33085_);
  and (_33139_, _33128_, _33063_);
  nor (_33150_, _29308_, _17379_);
  not (_33161_, _33150_);
  nor (_33172_, _28223_, _18414_);
  nor (_33183_, _28300_, _18588_);
  nor (_33194_, _33183_, _33172_);
  and (_33205_, _33194_, _33161_);
  and (_33216_, _33205_, _33139_);
  not (_33227_, _33216_);
  nor (_33238_, _33227_, _33041_);
  and (_33248_, _33238_, _32987_);
  not (_33269_, _33248_);
  nor (_33270_, _33269_, _32856_);
  and (_33281_, _33270_, _32823_);
  not (_33292_, _33281_);
  nor (_33303_, _33292_, _32758_);
  and (_33314_, _33303_, _32747_);
  not (_33325_, _33314_);
  or (_33336_, _33325_, _25733_);
  not (_33346_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_33357_, _25733_, _33346_);
  and (_33368_, _33357_, _28541_);
  and (_33379_, _33368_, _33336_);
  nor (_33390_, _28530_, _33346_);
  and (_33401_, _30414_, _29101_);
  and (_33412_, _33401_, _25722_);
  nand (_33423_, _33412_, _29090_);
  or (_33434_, _33412_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_33445_, _33434_, _29166_);
  and (_33455_, _33445_, _33423_);
  or (_33466_, _33455_, _33390_);
  or (_33477_, _33466_, _33379_);
  and (_08941_, _33477_, _41654_);
  and (_33498_, _24340_, _21515_);
  not (_33509_, _33498_);
  and (_33520_, _21450_, _16164_);
  nor (_33531_, _27006_, _26051_);
  nor (_33542_, _33531_, _27017_);
  nor (_33553_, _33542_, _25810_);
  not (_33563_, _33553_);
  nor (_33574_, _27390_, _27368_);
  not (_33585_, _33574_);
  nor (_33596_, _27488_, _27401_);
  and (_33607_, _33596_, _33585_);
  nor (_33618_, _26874_, _25854_);
  or (_33629_, _33618_, _27817_);
  nor (_33640_, _33629_, _28826_);
  or (_33651_, _26874_, _18414_);
  or (_33662_, _32921_, _27587_);
  and (_33672_, _33662_, _33651_);
  nor (_33683_, _33672_, _17390_);
  not (_33694_, _33683_);
  and (_33705_, _33672_, _17390_);
  nor (_33716_, _33705_, _30611_);
  and (_33727_, _33716_, _33694_);
  nor (_33738_, _33727_, _33640_);
  nor (_33749_, _33009_, _17379_);
  and (_33760_, _33009_, _17379_);
  nor (_33771_, _33760_, _33749_);
  nor (_33791_, _33771_, _28869_);
  nor (_33792_, _28103_, _25887_);
  and (_33803_, _28124_, _25898_);
  nor (_33814_, _33803_, _33792_);
  and (_33825_, _28157_, _25876_);
  and (_33836_, _28179_, _17379_);
  nor (_33847_, _33836_, _33825_);
  nor (_33858_, _28223_, _17379_);
  not (_33869_, _33858_);
  nor (_33880_, _29308_, _18218_);
  nor (_33891_, _28300_, _18414_);
  nor (_33901_, _33891_, _33880_);
  and (_33912_, _33901_, _33869_);
  and (_33923_, _33912_, _33847_);
  and (_33934_, _33923_, _33814_);
  not (_33945_, _33934_);
  nor (_33956_, _33945_, _33791_);
  and (_33967_, _33956_, _33738_);
  not (_33978_, _33967_);
  nor (_33989_, _33978_, _33607_);
  and (_34000_, _33989_, _33563_);
  not (_34010_, _34000_);
  nor (_34021_, _34010_, _33520_);
  and (_34032_, _34021_, _33509_);
  not (_34043_, _34032_);
  or (_34064_, _34043_, _25733_);
  not (_34065_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_34076_, _25733_, _34065_);
  and (_34086_, _34076_, _28541_);
  and (_34097_, _34086_, _34064_);
  nor (_34108_, _28530_, _34065_);
  nor (_34119_, _24645_, _24764_);
  and (_34130_, _34119_, _24884_);
  and (_34141_, _34130_, _25722_);
  nand (_34152_, _34141_, _29090_);
  or (_34163_, _34141_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_34174_, _34163_, _29166_);
  and (_34185_, _34174_, _34152_);
  or (_34196_, _34185_, _34108_);
  or (_34206_, _34196_, _34097_);
  and (_08952_, _34206_, _41654_);
  and (_34227_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_34238_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_34249_, _34238_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_34260_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_34271_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_34282_, _34271_, _34260_);
  and (_34293_, _34238_, _16098_);
  and (_34304_, _34293_, _34282_);
  not (_34314_, _34304_);
  and (_34325_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_34336_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_34347_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_34358_, _34347_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_34369_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_34380_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_34391_, _34380_, _34369_);
  and (_34402_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not (_34413_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_34424_, _34413_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34434_, _34424_, _34369_);
  and (_34445_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_34456_, _34445_, _34402_);
  and (_34467_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34478_, _34467_, _34369_);
  and (_34489_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not (_34500_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34511_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _34500_);
  and (_34522_, _34511_, _34369_);
  and (_34533_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_34544_, _34533_, _34489_);
  and (_34555_, _34380_, _34369_);
  and (_34565_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_34576_, _34380_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_34587_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_34598_, _34587_, _34565_);
  and (_34609_, _34598_, _34544_);
  and (_34620_, _34609_, _34456_);
  nor (_34631_, _34620_, _34358_);
  nor (_34642_, _34631_, _34336_);
  nor (_34653_, _34642_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34664_, _34653_, _34325_);
  nor (_34685_, _34664_, _34314_);
  and (_34686_, _34282_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_34696_, _34686_, _34314_);
  nor (_34707_, _34696_, _34685_);
  and (_34718_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34729_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_34740_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34751_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_34762_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_34773_, _34762_, _34751_);
  and (_34784_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34795_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_34806_, _34795_, _34784_);
  and (_34816_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_34827_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_34838_, _34827_, _34816_);
  and (_34849_, _34838_, _34806_);
  and (_34860_, _34849_, _34773_);
  nor (_34871_, _34860_, _34347_);
  and (_34882_, _34871_, _34740_);
  nor (_34893_, _34882_, _34729_);
  nor (_34904_, _34893_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34915_, _34904_, _34718_);
  nor (_34926_, _34915_, _34314_);
  and (_34937_, _34282_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_34948_, _34937_, _34314_);
  nor (_34959_, _34948_, _34926_);
  not (_34970_, _34959_);
  and (_34981_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34992_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35003_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_35014_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_35025_, _35014_, _35003_);
  and (_35036_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_35047_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_35058_, _35047_, _35036_);
  and (_35069_, _35058_, _35025_);
  and (_35080_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_35091_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_35102_, _35091_, _35080_);
  and (_35113_, _35102_, _35069_);
  nor (_35124_, _35113_, _34358_);
  nor (_35135_, _35124_, _34992_);
  nor (_35146_, _35135_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35157_, _35146_, _34981_);
  nor (_35168_, _35157_, _34314_);
  and (_35179_, _34282_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_35190_, _35179_, _34314_);
  nor (_35201_, _35190_, _35168_);
  nor (_35212_, _35201_, _34970_);
  and (_35223_, _35212_, _34707_);
  and (_35234_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not (_35245_, _35234_);
  and (_35256_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_35267_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_35278_, _35267_, _35256_);
  and (_35289_, _35278_, _35245_);
  and (_35300_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_35311_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_35322_, _35311_, _35300_);
  and (_35333_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_35344_, _34347_, _35333_);
  and (_35355_, _35344_, _35322_);
  and (_35366_, _35355_, _35289_);
  and (_35377_, _35366_, _34740_);
  nor (_35399_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _34740_);
  nor (_35400_, _35399_, _35377_);
  nor (_35422_, _35400_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_35423_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35445_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _35423_);
  nor (_35446_, _35445_, _35422_);
  and (_35468_, _35446_, _34304_);
  and (_35469_, _34282_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_35480_, _35469_, _34314_);
  nor (_35491_, _35480_, _35468_);
  and (_35502_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35513_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35524_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_35535_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_35546_, _35535_, _35524_);
  and (_35557_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_35568_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_35579_, _35568_, _35557_);
  and (_35590_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_35601_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_35612_, _35601_, _35590_);
  and (_35623_, _35612_, _35579_);
  and (_35634_, _35623_, _35546_);
  nor (_35645_, _34358_, _35634_);
  nor (_35656_, _35645_, _35513_);
  nor (_35667_, _35656_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35678_, _35667_, _35502_);
  nor (_35689_, _35678_, _34314_);
  and (_35700_, _34282_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_35711_, _35700_, _34314_);
  nor (_35722_, _35711_, _35689_);
  nor (_35733_, _35722_, _35491_);
  and (_35744_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35755_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35766_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_35777_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_35788_, _35777_, _35766_);
  and (_35799_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_35810_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_35821_, _35810_, _35799_);
  and (_35832_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_35843_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_35854_, _35843_, _35832_);
  and (_35865_, _35854_, _35821_);
  and (_35876_, _35865_, _35788_);
  nor (_35887_, _35876_, _34347_);
  and (_35898_, _35887_, _34740_);
  or (_35909_, _35898_, _35755_);
  and (_35920_, _35909_, _35423_);
  nor (_35931_, _35920_, _35744_);
  nor (_35942_, _35931_, _34314_);
  and (_35953_, _34282_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_35964_, _35953_, _34314_);
  nor (_35975_, _35964_, _35942_);
  and (_35986_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_35997_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_36008_, _35997_, _35986_);
  and (_36019_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_36030_, _36019_, _34347_);
  and (_36041_, _36030_, _36008_);
  and (_36052_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_36063_, _36052_);
  and (_36074_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_36085_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_36096_, _36085_, _36074_);
  and (_36107_, _36096_, _36063_);
  and (_36118_, _36107_, _36041_);
  and (_36129_, _36118_, _34740_);
  nor (_36140_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _34740_);
  or (_36151_, _36140_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_36162_, _36151_, _36129_);
  and (_36173_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_36184_, _36173_, _36162_);
  and (_36195_, _36184_, _34304_);
  and (_36206_, _34282_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_36217_, _36206_, _34314_);
  nor (_36228_, _36217_, _36195_);
  not (_36239_, _36228_);
  and (_36250_, _36239_, _35975_);
  and (_36261_, _36250_, _35733_);
  and (_36272_, _36261_, _35223_);
  and (_36283_, _35733_, _35975_);
  and (_36294_, _35201_, _34707_);
  and (_36305_, _36294_, _34970_);
  and (_36316_, _36305_, _36283_);
  or (_36326_, _36316_, _36272_);
  not (_36337_, _36326_);
  and (_36348_, _36294_, _34959_);
  and (_36359_, _36348_, _36283_);
  not (_36370_, _34707_);
  and (_36381_, _35201_, _36370_);
  and (_36392_, _36381_, _34970_);
  and (_36403_, _36392_, _36261_);
  nor (_36414_, _36403_, _36359_);
  not (_36425_, _36414_);
  and (_36436_, _36381_, _34959_);
  and (_36446_, _36436_, _36228_);
  and (_36457_, _36446_, _36283_);
  nor (_36468_, _36457_, _36425_);
  and (_36479_, _35975_, _35722_);
  and (_36490_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_36501_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_36512_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_36523_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_36534_, _36523_, _36512_);
  and (_36545_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_36556_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_36567_, _36556_, _36545_);
  and (_36578_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_36589_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_36600_, _36589_, _36578_);
  and (_36611_, _36600_, _36567_);
  and (_36622_, _36611_, _36534_);
  nor (_36633_, _36622_, _34347_);
  and (_36644_, _36633_, _34740_);
  nor (_36655_, _36644_, _36501_);
  nor (_36666_, _36655_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_36677_, _36666_, _36490_);
  nor (_36687_, _36677_, _34314_);
  and (_36698_, _34282_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_36709_, _36698_, _34314_);
  nor (_36720_, _36709_, _36687_);
  and (_36731_, _36720_, _35491_);
  and (_36742_, _36731_, _36479_);
  and (_36753_, _35212_, _36370_);
  and (_36764_, _36753_, _36239_);
  and (_36775_, _36764_, _36742_);
  not (_36786_, _35491_);
  and (_36796_, _36479_, _36786_);
  and (_36807_, _36796_, _36720_);
  and (_36818_, _36807_, _36305_);
  nor (_36829_, _36818_, _36775_);
  and (_36840_, _36829_, _36468_);
  and (_36851_, _36840_, _36337_);
  not (_36862_, _36720_);
  and (_36873_, _36796_, _36862_);
  and (_36884_, _36392_, _36228_);
  and (_36895_, _36884_, _36873_);
  not (_36905_, _36895_);
  and (_36916_, _36436_, _36239_);
  and (_36927_, _36916_, _36873_);
  nor (_36938_, _35201_, _34959_);
  and (_36949_, _36938_, _34707_);
  and (_36960_, _36949_, _36239_);
  and (_36971_, _36960_, _36873_);
  nor (_36982_, _36971_, _36927_);
  and (_36993_, _36982_, _36905_);
  and (_37004_, _36949_, _36228_);
  and (_37014_, _37004_, _36283_);
  not (_37025_, _37014_);
  and (_37036_, _36228_, _36283_);
  and (_37047_, _37036_, _35223_);
  and (_37058_, _36938_, _36370_);
  and (_37069_, _37058_, _37036_);
  or (_37080_, _37069_, _37047_);
  and (_37091_, _36753_, _36283_);
  and (_37102_, _36916_, _36283_);
  nor (_37113_, _37102_, _37091_);
  not (_37124_, _37113_);
  nor (_37135_, _37124_, _37080_);
  and (_37146_, _37135_, _37025_);
  and (_37157_, _37146_, _36993_);
  and (_37168_, _37157_, _36851_);
  nor (_37179_, _37168_, _34249_);
  not (_37189_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_37197_, _16098_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_37205_, _37197_, _37189_);
  and (_37212_, _37205_, _36949_);
  and (_37220_, _37212_, _36742_);
  and (_37228_, _36818_, _37197_);
  and (_37235_, _37228_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_37243_, _37235_, _37220_);
  nor (_37251_, _37243_, _37179_);
  nor (_37254_, _37251_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37255_, _37254_, _34227_);
  and (_37256_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_37265_, _36392_, _37036_);
  not (_37276_, _37265_);
  not (_37287_, _35722_);
  and (_37298_, _35975_, _37287_);
  nor (_37309_, _36720_, _36786_);
  and (_37320_, _37309_, _37298_);
  and (_37331_, _37058_, _36228_);
  and (_37342_, _37331_, _37320_);
  and (_37353_, _36381_, _36239_);
  and (_37364_, _37353_, _37320_);
  nor (_37375_, _37364_, _37342_);
  and (_37386_, _37375_, _37276_);
  and (_37397_, _35223_, _36239_);
  nor (_37408_, _37397_, _36305_);
  not (_37419_, _37320_);
  nor (_37429_, _37419_, _37408_);
  not (_37436_, _37429_);
  not (_37447_, _36818_);
  nor (_37458_, _36239_, _35975_);
  and (_37469_, _37458_, _36392_);
  and (_37480_, _36348_, _36228_);
  and (_37491_, _37480_, _37320_);
  nor (_37502_, _37491_, _37469_);
  and (_37513_, _37502_, _37447_);
  and (_37524_, _37513_, _37436_);
  and (_37535_, _37320_, _37004_);
  and (_37546_, _36753_, _36228_);
  and (_37557_, _37546_, _37320_);
  nor (_37568_, _37557_, _37535_);
  and (_37579_, _36884_, _36807_);
  and (_37590_, _36807_, _36764_);
  nor (_37601_, _37590_, _37579_);
  and (_37612_, _37601_, _37568_);
  and (_37623_, _37612_, _37524_);
  and (_37634_, _37623_, _37386_);
  and (_37645_, _36884_, _36742_);
  and (_37656_, _35223_, _36228_);
  and (_37667_, _37656_, _37320_);
  nor (_37678_, _37667_, _37645_);
  and (_37689_, _37656_, _36873_);
  and (_37700_, _37656_, _36807_);
  nor (_37711_, _37700_, _37689_);
  and (_37722_, _37711_, _37678_);
  and (_37733_, _36392_, _36239_);
  and (_37744_, _36807_, _37733_);
  and (_37755_, _37546_, _36807_);
  nor (_37766_, _37755_, _37744_);
  and (_37777_, _36348_, _36239_);
  and (_37788_, _37320_, _37777_);
  and (_37799_, _37320_, _36764_);
  nor (_37810_, _37799_, _37788_);
  and (_37821_, _37810_, _37766_);
  and (_37832_, _36742_, _37733_);
  and (_37843_, _36960_, _36807_);
  nor (_37854_, _37843_, _37832_);
  and (_37865_, _37854_, _37821_);
  and (_37876_, _37865_, _37722_);
  and (_37887_, _36807_, _36446_);
  and (_37898_, _36796_, _37397_);
  nor (_37909_, _37898_, _37887_);
  and (_37920_, _36916_, _36807_);
  and (_37931_, _37320_, _36446_);
  nor (_37942_, _37931_, _37920_);
  and (_37953_, _37942_, _37909_);
  and (_37964_, _36742_, _36305_);
  and (_37975_, _37964_, _36228_);
  not (_37986_, _36742_);
  and (_37997_, _36239_, _36305_);
  nor (_38008_, _37997_, _37777_);
  nor (_38019_, _38008_, _37986_);
  nor (_38030_, _38019_, _37975_);
  and (_38041_, _36753_, _36742_);
  and (_38052_, _37004_, _36796_);
  nor (_38063_, _38052_, _38041_);
  and (_38074_, _38063_, _38030_);
  and (_38084_, _38074_, _37953_);
  and (_38095_, _38084_, _37876_);
  and (_38106_, _38095_, _37634_);
  nor (_38116_, _38106_, _34249_);
  and (_38127_, _37197_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_38138_, _38127_, _36818_);
  not (_38149_, _38138_);
  nor (_38160_, _35201_, _36370_);
  and (_38171_, _36742_, _38160_);
  and (_38182_, _38171_, _37205_);
  not (_38186_, _37205_);
  and (_38187_, _36228_, _36305_);
  and (_38188_, _38187_, _36742_);
  and (_38189_, _36742_, _37777_);
  nor (_38190_, _38189_, _38188_);
  nor (_38191_, _38190_, _38186_);
  nor (_38192_, _38191_, _38182_);
  and (_38193_, _38192_, _38149_);
  not (_38194_, _38193_);
  nor (_38195_, _38194_, _38116_);
  nor (_38196_, _38195_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38197_, _38196_, _37256_);
  nor (_38198_, _38197_, _37255_);
  and (_38199_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38200_, _36731_, _37298_);
  and (_38201_, _38200_, _36446_);
  and (_38202_, _38200_, _36884_);
  nor (_38203_, _38202_, _38201_);
  and (_38204_, _38203_, _36993_);
  nor (_38205_, _38204_, _34249_);
  nor (_38206_, _38205_, _38182_);
  not (_38207_, _34249_);
  nor (_38208_, _38203_, _38207_);
  not (_38209_, _38208_);
  and (_38210_, _38209_, _38206_);
  nor (_38211_, _38210_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38212_, _38211_, _38199_);
  and (_38213_, _38212_, _41654_);
  and (_09497_, _38213_, _38198_);
  and (_38214_, _25253_, _25122_);
  nor (_38215_, _25689_, _25395_);
  and (_38216_, _38215_, _38214_);
  and (_38217_, _30414_, _24645_);
  and (_38218_, _38217_, _25548_);
  and (_38219_, _38218_, _38216_);
  and (_38220_, _38219_, _28530_);
  and (_38221_, _38220_, _28497_);
  not (_38222_, _38221_);
  and (_38223_, _38222_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_38224_, _38216_, _25548_);
  and (_38225_, _38224_, _24645_);
  and (_38226_, _38225_, _30414_);
  and (_38227_, _38226_, _28541_);
  not (_38228_, _38227_);
  nor (_38229_, _21515_, _16164_);
  and (_38230_, _27466_, _21493_);
  nor (_38231_, _28289_, _38230_);
  and (_38232_, _38231_, _28223_);
  and (_38233_, _38232_, _38229_);
  and (_38234_, _38233_, _29308_);
  nor (_38235_, _38234_, _17379_);
  not (_38236_, _38235_);
  and (_38237_, _38236_, _33847_);
  and (_38238_, _38237_, _33814_);
  and (_38239_, _38238_, _33738_);
  nor (_38240_, _38239_, _38228_);
  nor (_38241_, _38240_, _38223_);
  and (_38242_, _38222_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38243_, _38234_, _18414_);
  not (_38244_, _38243_);
  and (_38245_, _38244_, _33139_);
  and (_38246_, _38245_, _32987_);
  nor (_38247_, _38246_, _38228_);
  nor (_38248_, _38247_, _38242_);
  and (_38249_, _38222_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38250_, _38234_, _18588_);
  not (_38251_, _38250_);
  and (_38252_, _38251_, _32334_);
  and (_38253_, _38252_, _32203_);
  nor (_38254_, _38253_, _38228_);
  nor (_38255_, _38254_, _38249_);
  and (_38256_, _38222_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38257_, _38234_, _18925_);
  not (_38258_, _38257_);
  and (_38259_, _38258_, _31353_);
  and (_38260_, _38259_, _31582_);
  and (_38261_, _38260_, _31550_);
  nor (_38262_, _38261_, _38228_);
  nor (_38263_, _38262_, _38256_);
  and (_38264_, _38222_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38265_, _38234_, _19448_);
  not (_38266_, _38265_);
  and (_38267_, _38266_, _30731_);
  and (_38268_, _38267_, _30764_);
  and (_38269_, _38268_, _30655_);
  nor (_38270_, _38269_, _38228_);
  nor (_38271_, _38270_, _38264_);
  and (_38272_, _38222_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38273_, _38234_, _19273_);
  not (_38274_, _38273_);
  and (_38275_, _38274_, _30107_);
  and (_38276_, _38275_, _29888_);
  not (_38277_, _38276_);
  and (_38278_, _38277_, _38227_);
  nor (_38279_, _38278_, _38272_);
  nor (_38280_, _38221_, _24808_);
  nor (_38281_, _38234_, _19819_);
  not (_38282_, _38281_);
  and (_38283_, _38282_, _29396_);
  and (_38284_, _38283_, _29560_);
  and (_38285_, _38284_, _29286_);
  not (_38286_, _38285_);
  and (_38287_, _38286_, _38227_);
  nor (_38288_, _38287_, _38280_);
  and (_38289_, _38288_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38290_, _38289_, _38279_);
  and (_38291_, _38290_, _38271_);
  and (_38292_, _38291_, _38263_);
  and (_38293_, _38292_, _38255_);
  and (_38294_, _38293_, _38248_);
  and (_38295_, _38294_, _38241_);
  nor (_38296_, _38221_, _25265_);
  nand (_38297_, _38296_, _38295_);
  or (_38298_, _38296_, _38295_);
  and (_38299_, _38298_, _24971_);
  and (_38300_, _38299_, _38297_);
  or (_38301_, _38221_, _25308_);
  or (_38302_, _38301_, _38300_);
  nor (_38303_, _38234_, _18218_);
  not (_38304_, _38303_);
  and (_38305_, _38304_, _28201_);
  and (_38306_, _38305_, _28146_);
  and (_38307_, _38306_, _27850_);
  nand (_38308_, _38307_, _38221_);
  and (_38309_, _38308_, _38302_);
  and (_09517_, _38309_, _41654_);
  not (_38310_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38311_, _38288_, _38310_);
  nor (_38312_, _38288_, _38310_);
  nor (_38313_, _38312_, _38311_);
  and (_38314_, _38313_, _24971_);
  nor (_38315_, _38314_, _24819_);
  nor (_38316_, _38315_, _38227_);
  nor (_38317_, _38316_, _38287_);
  nand (_10643_, _38317_, _41654_);
  nor (_38318_, _38289_, _38279_);
  nor (_38319_, _38318_, _38290_);
  nor (_38320_, _38319_, _24448_);
  nor (_38321_, _38320_, _24688_);
  nor (_38322_, _38321_, _38227_);
  nor (_38323_, _38322_, _38278_);
  nand (_10654_, _38323_, _41654_);
  nor (_38324_, _38290_, _38271_);
  nor (_38325_, _38324_, _38291_);
  nor (_38326_, _38325_, _24448_);
  nor (_38327_, _38326_, _24503_);
  nor (_38328_, _38327_, _38227_);
  nor (_38329_, _38328_, _38270_);
  nand (_10665_, _38329_, _41654_);
  nor (_38330_, _38291_, _38263_);
  nor (_38331_, _38330_, _38292_);
  nor (_38332_, _38331_, _24448_);
  nor (_38333_, _38332_, _25483_);
  nor (_38334_, _38333_, _38227_);
  nor (_38335_, _38334_, _38262_);
  nor (_10676_, _38335_, rst);
  nor (_38336_, _38292_, _38255_);
  or (_38337_, _38336_, _38293_);
  and (_38338_, _38337_, _24971_);
  or (_38339_, _38338_, _25580_);
  and (_38340_, _38339_, _38228_);
  or (_38341_, _38340_, _38254_);
  and (_10687_, _38341_, _41654_);
  nor (_38342_, _38293_, _38248_);
  nor (_38343_, _38342_, _38294_);
  nor (_38344_, _38343_, _24448_);
  nor (_38345_, _38344_, _25156_);
  nor (_38346_, _38345_, _38227_);
  nor (_38347_, _38346_, _38247_);
  nor (_10698_, _38347_, rst);
  nor (_38348_, _38294_, _38241_);
  nor (_38349_, _38348_, _38295_);
  nor (_38350_, _38349_, _24448_);
  nor (_38351_, _38350_, _25004_);
  nor (_38352_, _38351_, _38227_);
  nor (_38353_, _38352_, _38240_);
  nor (_10709_, _38353_, rst);
  and (_38354_, _28541_, _25548_);
  and (_38355_, _38354_, _31822_);
  nand (_38356_, _38355_, _38216_);
  nor (_38357_, _38356_, _28465_);
  and (_38358_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _16098_);
  and (_38359_, _38358_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38360_, _38356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38361_, _38360_, _38359_);
  or (_38362_, _38361_, _38357_);
  nor (_38363_, _28223_, _18043_);
  nor (_38364_, _28684_, _18925_);
  and (_38365_, _27598_, _18228_);
  and (_38366_, _38365_, _26238_);
  and (_38367_, _38366_, _26271_);
  and (_38368_, _38367_, _26315_);
  and (_38369_, _38368_, _26939_);
  nor (_38370_, _38369_, _27620_);
  and (_38371_, _26874_, _16724_);
  nor (_38372_, _38371_, _38370_);
  and (_38373_, _27686_, _18218_);
  and (_38374_, _17553_, _16559_);
  and (_38375_, _17869_, _16888_);
  and (_38376_, _38375_, _38374_);
  and (_38377_, _38376_, _38373_);
  and (_38378_, _17705_, _16724_);
  and (_38379_, _38378_, _38377_);
  nor (_38380_, _38379_, _26874_);
  and (_38381_, _26874_, _17705_);
  nor (_38382_, _38381_, _38380_);
  and (_38383_, _38382_, _38372_);
  nor (_38384_, _26874_, _17064_);
  and (_38385_, _26874_, _17064_);
  nor (_38386_, _38385_, _38384_);
  and (_38387_, _38386_, _38383_);
  and (_38388_, _38387_, _27763_);
  nor (_38389_, _38387_, _27763_);
  nor (_38390_, _38389_, _38388_);
  and (_38391_, _38390_, _27532_);
  and (_38392_, _26874_, _27763_);
  nor (_38393_, _38392_, _28870_);
  nor (_38394_, _38393_, _27817_);
  or (_38395_, _38394_, _38391_);
  or (_38396_, _38395_, _38364_);
  and (_38397_, _21515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_38398_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38399_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38400_, _38399_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38401_, _38400_, _38398_);
  nor (_38402_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38403_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38404_, _38403_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38405_, _38404_, _38402_);
  nor (_38406_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38407_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38408_, _38407_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38409_, _38408_, _38406_);
  not (_38410_, _38409_);
  nor (_38411_, _38410_, _28607_);
  nor (_38412_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38413_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38414_, _38413_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38415_, _38414_, _38412_);
  and (_38416_, _38415_, _38411_);
  nor (_38417_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38418_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38419_, _38418_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38420_, _38419_, _38417_);
  and (_38421_, _38420_, _38416_);
  and (_38422_, _38421_, _38405_);
  nor (_38423_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38424_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38425_, _38424_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38426_, _38425_, _38423_);
  and (_38427_, _38426_, _38422_);
  and (_38428_, _38427_, _38401_);
  nor (_38429_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38430_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38431_, _38430_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38432_, _38431_, _38429_);
  and (_38433_, _38432_, _38428_);
  nor (_38434_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38435_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38436_, _38435_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38437_, _38436_, _38434_);
  nand (_38438_, _38437_, _38433_);
  or (_38439_, _38437_, _38433_);
  and (_38440_, _38439_, _27477_);
  and (_38441_, _38440_, _38438_);
  and (_38442_, _21201_, _16164_);
  or (_38443_, _38442_, _38441_);
  or (_38444_, _38443_, _38397_);
  or (_38445_, _38444_, _38396_);
  nor (_38446_, _38445_, _38363_);
  nand (_38447_, _38446_, _38359_);
  and (_38448_, _38447_, _41654_);
  and (_12656_, _38448_, _38362_);
  and (_38449_, _38354_, _31124_);
  and (_38450_, _38449_, _38216_);
  nor (_38451_, _38450_, _38359_);
  not (_38452_, _38451_);
  nand (_38453_, _38452_, _28465_);
  or (_38454_, _38452_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38455_, _38454_, _41654_);
  and (_12677_, _38455_, _38453_);
  nor (_38456_, _38356_, _29615_);
  and (_38457_, _38356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38458_, _38457_, _38359_);
  or (_38459_, _38458_, _38456_);
  nor (_38460_, _28223_, _16888_);
  nor (_38461_, _28684_, _18588_);
  nor (_38462_, _28870_, _27795_);
  not (_38463_, _38462_);
  nor (_38464_, _38463_, _27708_);
  nor (_38465_, _38464_, _26238_);
  and (_38466_, _38464_, _26238_);
  or (_38467_, _38466_, _30611_);
  nor (_38468_, _38467_, _38465_);
  nor (_38469_, _27817_, _19819_);
  or (_38470_, _38469_, _38468_);
  or (_38471_, _38470_, _38461_);
  and (_38472_, _23800_, _21515_);
  and (_38473_, _38410_, _28607_);
  nor (_38474_, _38473_, _38411_);
  and (_38475_, _38474_, _27477_);
  and (_38476_, _20980_, _16164_);
  or (_38477_, _38476_, _38475_);
  or (_38478_, _38477_, _38472_);
  or (_38479_, _38478_, _38471_);
  nor (_38480_, _38479_, _38460_);
  nand (_38481_, _38480_, _38359_);
  and (_38482_, _38481_, _41654_);
  and (_13571_, _38482_, _38459_);
  nor (_38483_, _38356_, _30294_);
  and (_38484_, _38356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38485_, _38484_, _38359_);
  or (_38486_, _38485_, _38483_);
  nor (_38487_, _28223_, _17869_);
  nor (_38488_, _28684_, _18414_);
  nor (_38489_, _38366_, _27620_);
  and (_38490_, _38373_, _16888_);
  nor (_38491_, _38490_, _26874_);
  or (_38492_, _38491_, _38489_);
  nor (_38493_, _38492_, _26271_);
  and (_38494_, _38492_, _26271_);
  nor (_38495_, _38494_, _38493_);
  nor (_38496_, _38495_, _30611_);
  nor (_38497_, _27817_, _19273_);
  or (_38498_, _38497_, _38496_);
  or (_38499_, _38498_, _38488_);
  and (_38500_, _22798_, _21515_);
  nor (_38501_, _38415_, _38411_);
  not (_38502_, _38501_);
  nor (_38503_, _38416_, _27488_);
  and (_38504_, _38503_, _38502_);
  and (_38505_, _21012_, _16164_);
  or (_38506_, _38505_, _38504_);
  or (_38507_, _38506_, _38500_);
  or (_38508_, _38507_, _38499_);
  nor (_38509_, _38508_, _38487_);
  nand (_38510_, _38509_, _38359_);
  and (_38511_, _38510_, _41654_);
  and (_13580_, _38511_, _38486_);
  nor (_38512_, _38356_, _30993_);
  and (_38513_, _38356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38514_, _38513_, _38359_);
  or (_38515_, _38514_, _38512_);
  nor (_38516_, _28223_, _16559_);
  nor (_38517_, _28684_, _17379_);
  and (_38518_, _38490_, _17869_);
  and (_38519_, _38518_, _27620_);
  and (_38520_, _38367_, _26874_);
  nor (_38521_, _38520_, _38519_);
  and (_38522_, _38521_, _16559_);
  nor (_38523_, _38521_, _16559_);
  nor (_38524_, _38523_, _38522_);
  and (_38525_, _38524_, _27532_);
  nor (_38526_, _27817_, _19448_);
  or (_38527_, _38526_, _38525_);
  or (_38528_, _38527_, _38517_);
  and (_38529_, _21515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38530_, _38420_, _38416_);
  nor (_38531_, _38530_, _38421_);
  and (_38532_, _38531_, _27477_);
  and (_38533_, _21043_, _16164_);
  or (_38534_, _38533_, _38532_);
  or (_38535_, _38534_, _38529_);
  or (_38536_, _38535_, _38528_);
  nor (_38537_, _38536_, _38516_);
  nand (_38538_, _38537_, _38359_);
  and (_38539_, _38538_, _41654_);
  and (_13591_, _38539_, _38515_);
  nor (_38540_, _38356_, _31724_);
  and (_38541_, _38356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38542_, _38541_, _38359_);
  or (_38543_, _38542_, _38540_);
  nor (_38544_, _28223_, _17553_);
  nor (_38545_, _38368_, _26939_);
  not (_38546_, _38545_);
  and (_38547_, _38546_, _38370_);
  and (_38548_, _38518_, _16559_);
  nor (_38549_, _38548_, _17553_);
  nor (_38550_, _38549_, _38377_);
  nor (_38551_, _38550_, _26874_);
  nor (_38552_, _38551_, _38547_);
  nor (_38553_, _38552_, _30611_);
  nor (_38554_, _27817_, _18925_);
  or (_38555_, _38554_, _38553_);
  or (_38556_, _38555_, _28695_);
  and (_38557_, _21515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_38558_, _38421_, _38405_);
  nor (_38559_, _38558_, _38422_);
  and (_38560_, _38559_, _27477_);
  and (_38561_, _21075_, _16164_);
  or (_38562_, _38561_, _38560_);
  or (_38563_, _38562_, _38557_);
  or (_38564_, _38563_, _38556_);
  nor (_38565_, _38564_, _38544_);
  nand (_38566_, _38565_, _38359_);
  and (_38567_, _38566_, _41654_);
  and (_13600_, _38567_, _38543_);
  nor (_38568_, _38356_, _32486_);
  and (_38569_, _38356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38570_, _38569_, _38359_);
  or (_38571_, _38570_, _38568_);
  nor (_38572_, _28223_, _16724_);
  nor (_38573_, _28684_, _19819_);
  nor (_38574_, _38377_, _26874_);
  nor (_38575_, _38574_, _38370_);
  and (_38576_, _38575_, _16724_);
  nor (_38577_, _38575_, _16724_);
  nor (_38578_, _38577_, _38576_);
  nor (_38579_, _38578_, _30611_);
  nor (_38580_, _26874_, _18599_);
  or (_38581_, _38580_, _27817_);
  nor (_38582_, _38581_, _38371_);
  or (_38583_, _38582_, _38579_);
  or (_38584_, _38583_, _38573_);
  and (_38585_, _21515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38586_, _38426_, _38422_);
  not (_38587_, _38586_);
  nor (_38588_, _38427_, _27488_);
  and (_38589_, _38588_, _38587_);
  and (_38590_, _21106_, _16164_);
  or (_38591_, _38590_, _38589_);
  or (_38592_, _38591_, _38585_);
  or (_38593_, _38592_, _38584_);
  nor (_38594_, _38593_, _38572_);
  nand (_38595_, _38594_, _38359_);
  and (_38596_, _38595_, _41654_);
  and (_13610_, _38596_, _38571_);
  nor (_38597_, _38356_, _33314_);
  and (_38598_, _38356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38599_, _38598_, _38359_);
  or (_38600_, _38599_, _38597_);
  nor (_38601_, _28223_, _17705_);
  nor (_38602_, _28684_, _19273_);
  and (_38603_, _38377_, _16724_);
  nor (_38604_, _38603_, _26874_);
  not (_38605_, _38604_);
  and (_38606_, _38605_, _38372_);
  and (_38607_, _38606_, _17705_);
  nor (_38608_, _38606_, _17705_);
  nor (_38609_, _38608_, _38607_);
  nor (_38610_, _38609_, _30611_);
  nor (_38611_, _26874_, _18425_);
  or (_38612_, _38611_, _27817_);
  nor (_38613_, _38612_, _38381_);
  or (_38614_, _38613_, _38610_);
  or (_38615_, _38614_, _38602_);
  and (_38616_, _21515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_38617_, _38427_, _38401_);
  not (_38618_, _38617_);
  nor (_38619_, _38428_, _27488_);
  and (_38620_, _38619_, _38618_);
  and (_38621_, _21138_, _16164_);
  or (_38622_, _38621_, _38620_);
  or (_38623_, _38622_, _38616_);
  or (_38624_, _38623_, _38615_);
  nor (_38626_, _38624_, _38601_);
  nand (_38629_, _38626_, _38359_);
  and (_38630_, _38629_, _41654_);
  and (_13619_, _38630_, _38600_);
  nor (_38631_, _38356_, _34032_);
  and (_38632_, _38356_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38633_, _38632_, _38359_);
  or (_38634_, _38633_, _38631_);
  nor (_38635_, _28223_, _17064_);
  nor (_38636_, _28684_, _19448_);
  and (_38637_, _38383_, _17064_);
  nor (_38638_, _38383_, _17064_);
  nor (_38647_, _38638_, _38637_);
  nor (_38653_, _38647_, _30611_);
  nor (_38659_, _26874_, _17390_);
  or (_38663_, _38659_, _27817_);
  nor (_38664_, _38663_, _38385_);
  or (_38665_, _38664_, _38653_);
  or (_38666_, _38665_, _38636_);
  and (_38667_, _21515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_38668_, _38432_, _38428_);
  nor (_38669_, _38668_, _38433_);
  and (_38670_, _38669_, _27477_);
  and (_38671_, _21170_, _16164_);
  or (_38672_, _38671_, _38670_);
  or (_38673_, _38672_, _38667_);
  or (_38674_, _38673_, _38666_);
  nor (_38675_, _38674_, _38635_);
  nand (_38676_, _38675_, _38359_);
  and (_38677_, _38676_, _41654_);
  and (_13628_, _38677_, _38634_);
  nand (_38678_, _38452_, _29615_);
  or (_38679_, _38452_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_38680_, _38679_, _41654_);
  and (_13638_, _38680_, _38678_);
  nand (_38681_, _38452_, _30294_);
  or (_38682_, _38452_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38683_, _38682_, _41654_);
  and (_13648_, _38683_, _38681_);
  nand (_38684_, _38452_, _30993_);
  or (_38686_, _38452_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38688_, _38686_, _41654_);
  and (_13657_, _38688_, _38684_);
  nand (_38689_, _38452_, _31724_);
  or (_38690_, _38452_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38691_, _38690_, _41654_);
  and (_13667_, _38691_, _38689_);
  nand (_38692_, _38452_, _32486_);
  or (_38693_, _38452_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38694_, _38693_, _41654_);
  and (_13676_, _38694_, _38692_);
  nand (_38695_, _38452_, _33314_);
  or (_38696_, _38452_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38697_, _38696_, _41654_);
  and (_13686_, _38697_, _38695_);
  nand (_38698_, _38452_, _34032_);
  or (_38699_, _38452_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38700_, _38699_, _41654_);
  and (_13696_, _38700_, _38698_);
  and (_38701_, _28541_, _24906_);
  nor (_38702_, _25122_, _25395_);
  and (_38703_, _25700_, _25253_);
  and (_38704_, _38703_, _38702_);
  and (_38705_, _38704_, _38701_);
  nand (_38706_, _38705_, _38307_);
  and (_38707_, _38704_, _29166_);
  not (_38708_, _29122_);
  nor (_38709_, _38708_, _29090_);
  not (_38710_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38711_, _29122_, _38710_);
  or (_38712_, _38711_, _38709_);
  and (_38713_, _38712_, _38707_);
  nor (_38714_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_38715_, _38714_);
  nand (_38716_, _38715_, _29090_);
  and (_38717_, _38714_, _38710_);
  nor (_38718_, _38717_, _38707_);
  and (_38719_, _38718_, _38716_);
  or (_38721_, _38719_, _38705_);
  or (_38724_, _38721_, _38713_);
  and (_38730_, _38724_, _38706_);
  and (_16448_, _38730_, _41654_);
  not (_38741_, _38705_);
  nor (_38748_, _38741_, _38276_);
  not (_38758_, _25122_);
  and (_38759_, _38703_, _38758_);
  not (_38760_, _29166_);
  nor (_38761_, _38760_, _25395_);
  and (_38762_, _38761_, _38759_);
  and (_38763_, _38762_, _38217_);
  or (_38764_, _38763_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_38765_, _38764_, _38741_);
  nand (_38766_, _38763_, _29090_);
  and (_38767_, _38766_, _38765_);
  or (_38768_, _38767_, _38748_);
  and (_21381_, _38768_, _41654_);
  nor (_38769_, _38741_, _38269_);
  or (_38770_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_38771_, _21265_, _21233_);
  or (_38772_, _38771_, _21296_);
  or (_38773_, _38772_, _21339_);
  or (_38774_, _38773_, _21370_);
  or (_38775_, _38774_, _21427_);
  or (_38776_, _38775_, _21450_);
  or (_38777_, _38776_, _20917_);
  and (_38778_, _38777_, _16164_);
  not (_38779_, _25821_);
  nand (_38780_, _27422_, _38779_);
  or (_38781_, _27422_, _25832_);
  and (_38782_, _27477_, _38781_);
  and (_38783_, _38782_, _38780_);
  and (_38784_, _38378_, _22700_);
  and (_38785_, _38376_, _21515_);
  nand (_38786_, _38785_, _38784_);
  nand (_38787_, _38786_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_38788_, _38787_, _38783_);
  or (_38789_, _28651_, _27028_);
  not (_38790_, _28640_);
  nand (_38791_, _38790_, _27028_);
  and (_38792_, _38791_, _25799_);
  and (_38793_, _38792_, _38789_);
  or (_38794_, _38793_, _38788_);
  or (_38798_, _38794_, _38778_);
  and (_38809_, _38798_, _38770_);
  or (_38812_, _38809_, _38707_);
  nand (_38813_, _31135_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand (_38814_, _38813_, _38707_);
  or (_38823_, _38814_, _31146_);
  and (_38831_, _38823_, _38741_);
  and (_38832_, _38831_, _38812_);
  or (_38833_, _38832_, _38769_);
  and (_21392_, _38833_, _41654_);
  not (_38834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_38835_, _38707_, _31822_);
  nand (_38836_, _38835_, _38834_);
  and (_38837_, _38836_, _38741_);
  or (_38838_, _38835_, _29703_);
  and (_38839_, _38838_, _38837_);
  nor (_38840_, _38741_, _38261_);
  or (_38841_, _38840_, _38839_);
  and (_21404_, _38841_, _41654_);
  not (_38842_, _38762_);
  or (_38843_, _38842_, _32606_);
  and (_38844_, _38843_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_38845_, _32595_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_38846_, _38845_, _32639_);
  and (_38847_, _38846_, _38707_);
  or (_38848_, _38847_, _38844_);
  and (_38849_, _38848_, _38741_);
  nor (_38850_, _38741_, _38253_);
  or (_38851_, _38850_, _38849_);
  and (_21416_, _38851_, _41654_);
  nor (_38852_, _38741_, _38246_);
  and (_38853_, _38762_, _33401_);
  or (_38854_, _38853_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_38855_, _38854_, _38741_);
  nand (_38856_, _38853_, _29090_);
  and (_38857_, _38856_, _38855_);
  or (_38858_, _38857_, _38852_);
  and (_21428_, _38858_, _41654_);
  nor (_38859_, _38741_, _38239_);
  and (_38860_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_38861_, _27477_, _27346_);
  and (_38862_, _26984_, _25799_);
  or (_38863_, _38862_, _38861_);
  and (_38864_, _38863_, _38860_);
  nand (_38865_, _38860_, _28223_);
  and (_38866_, _38865_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_38867_, _38866_, _38707_);
  or (_38868_, _38867_, _38864_);
  not (_38869_, _34130_);
  nor (_38870_, _38869_, _29090_);
  nor (_38871_, _34130_, _31593_);
  or (_38872_, _38871_, _38870_);
  or (_38873_, _38872_, _38842_);
  and (_38874_, _38873_, _38868_);
  and (_38875_, _38874_, _38741_);
  or (_38876_, _38875_, _38859_);
  and (_21439_, _38876_, _41654_);
  not (_38877_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38878_, _38358_, _38877_);
  and (_38879_, _38878_, _38446_);
  nor (_38880_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38881_, _38880_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not (_38882_, _25253_);
  and (_38883_, _25678_, _38882_);
  and (_38884_, _38354_, _24906_);
  and (_38885_, _38884_, _38883_);
  and (_38886_, _38885_, _38702_);
  nor (_38887_, _38886_, _38881_);
  nor (_38888_, _38887_, _28465_);
  and (_38889_, _25678_, _25548_);
  and (_38890_, _38889_, _25254_);
  and (_38891_, _38890_, _38761_);
  and (_38892_, _38891_, _29122_);
  and (_38893_, _38892_, _29090_);
  nor (_38894_, _38892_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_38895_, _38878_);
  and (_38896_, _38887_, _38895_);
  not (_38897_, _38896_);
  nor (_38898_, _38897_, _38894_);
  not (_38899_, _38898_);
  nor (_38900_, _38899_, _38893_);
  nor (_38901_, _38900_, _38878_);
  not (_38902_, _38901_);
  nor (_38903_, _38902_, _38888_);
  nor (_38904_, _38903_, _38879_);
  and (_22209_, _38904_, _41654_);
  nor (_38905_, _38887_, _29615_);
  and (_38906_, _38891_, _24906_);
  and (_38907_, _38906_, _29090_);
  nor (_38908_, _38906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38909_, _38908_, _38897_);
  not (_38910_, _38909_);
  nor (_38911_, _38910_, _38907_);
  or (_38912_, _38911_, _38905_);
  and (_38913_, _38912_, _38895_);
  nor (_38914_, _38895_, _38480_);
  or (_38915_, _38914_, _38913_);
  and (_24064_, _38915_, _41654_);
  and (_38916_, _38878_, _38509_);
  nor (_38917_, _38887_, _30294_);
  and (_38918_, _38891_, _38217_);
  and (_38919_, _38918_, _29090_);
  nor (_38920_, _38918_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_38921_, _38920_, _38897_);
  not (_38922_, _38921_);
  nor (_38923_, _38922_, _38919_);
  nor (_38924_, _38923_, _38878_);
  not (_38925_, _38924_);
  nor (_38926_, _38925_, _38917_);
  nor (_38927_, _38926_, _38916_);
  and (_24075_, _38927_, _41654_);
  nor (_38928_, _38887_, _30993_);
  and (_38929_, _38891_, _31124_);
  and (_38930_, _38929_, _29090_);
  nor (_38931_, _38929_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_38932_, _38931_, _38897_);
  not (_38933_, _38932_);
  nor (_38934_, _38933_, _38930_);
  or (_38935_, _38934_, _38928_);
  and (_38936_, _38935_, _38895_);
  nor (_38937_, _38895_, _38537_);
  or (_38938_, _38937_, _38936_);
  and (_24087_, _38938_, _41654_);
  nor (_38939_, _38887_, _31724_);
  not (_38940_, _38891_);
  and (_38941_, _38896_, _38940_);
  and (_38942_, _38941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38943_, _31833_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_38944_, _38943_, _31844_);
  and (_38945_, _38891_, _38895_);
  not (_38946_, _38945_);
  nor (_38947_, _38946_, _38944_);
  and (_38948_, _38947_, _38896_);
  nor (_38949_, _38948_, _38942_);
  and (_38950_, _38949_, _38895_);
  not (_38951_, _38950_);
  nor (_38952_, _38951_, _38939_);
  and (_38953_, _38878_, _38565_);
  or (_38954_, _38953_, _38952_);
  nor (_24099_, _38954_, rst);
  nor (_38955_, _38887_, _32486_);
  and (_38956_, _38891_, _32584_);
  and (_38957_, _38956_, _29090_);
  nor (_38958_, _38956_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_38959_, _38958_, _38897_);
  not (_38960_, _38959_);
  nor (_38961_, _38960_, _38957_);
  or (_38962_, _38961_, _38955_);
  and (_38963_, _38962_, _38895_);
  nor (_38964_, _38895_, _38594_);
  or (_38965_, _38964_, _38963_);
  and (_24111_, _38965_, _41654_);
  nor (_38966_, _38887_, _33314_);
  and (_38967_, _38891_, _33401_);
  and (_38968_, _38967_, _29090_);
  nor (_38969_, _38967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_38970_, _38969_, _38897_);
  not (_38971_, _38970_);
  nor (_38972_, _38971_, _38968_);
  or (_38973_, _38972_, _38966_);
  and (_38974_, _38973_, _38895_);
  nor (_38975_, _38895_, _38626_);
  or (_38976_, _38975_, _38974_);
  and (_24123_, _38976_, _41654_);
  nor (_38977_, _38887_, _34032_);
  and (_38978_, _38891_, _34130_);
  and (_38979_, _38978_, _29090_);
  nor (_38980_, _38978_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_38981_, _38980_, _38897_);
  not (_38982_, _38981_);
  nor (_38983_, _38982_, _38979_);
  or (_38984_, _38983_, _38977_);
  and (_38985_, _38984_, _38895_);
  nor (_38986_, _38895_, _38675_);
  or (_38987_, _38986_, _38985_);
  and (_24135_, _38987_, _41654_);
  and (_38988_, _38224_, _29122_);
  nand (_38989_, _38988_, _29090_);
  or (_38990_, _38988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_38991_, _38990_, _29166_);
  and (_38992_, _38991_, _38989_);
  and (_38993_, _24906_, _25548_);
  and (_38994_, _38216_, _38993_);
  nand (_38995_, _38994_, _38307_);
  or (_38996_, _38994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_38997_, _38996_, _28541_);
  and (_38998_, _38997_, _38995_);
  not (_38999_, _28530_);
  and (_39000_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_39001_, _39000_, rst);
  or (_39002_, _39001_, _38998_);
  or (_35388_, _39002_, _38992_);
  nor (_39003_, _38758_, _25395_);
  and (_39004_, _38703_, _39003_);
  and (_39011_, _39004_, _29122_);
  nand (_39022_, _39011_, _29090_);
  or (_39033_, _39011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39043_, _39033_, _29166_);
  and (_39049_, _39043_, _39022_);
  and (_39059_, _39004_, _24906_);
  not (_39070_, _39059_);
  nor (_39081_, _39070_, _38307_);
  and (_39092_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_39103_, _39092_, _39081_);
  and (_39114_, _39103_, _28541_);
  and (_39125_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_39136_, _39125_, rst);
  or (_39147_, _39136_, _39114_);
  or (_35411_, _39147_, _39049_);
  and (_39168_, _38882_, _25122_);
  and (_39179_, _39168_, _38889_);
  and (_39190_, _39179_, _25406_);
  and (_39201_, _39190_, _29122_);
  nand (_39212_, _39201_, _29090_);
  or (_39218_, _39201_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39219_, _39218_, _29166_);
  and (_39220_, _39219_, _39212_);
  and (_39221_, _38883_, _39003_);
  and (_39222_, _39221_, _38993_);
  not (_39223_, _39222_);
  nor (_39224_, _39223_, _38307_);
  and (_39225_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_39226_, _39225_, _39224_);
  and (_39227_, _39226_, _28541_);
  and (_39228_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_39229_, _39228_, rst);
  or (_39230_, _39229_, _39227_);
  or (_35434_, _39230_, _39220_);
  and (_39231_, _39168_, _25711_);
  and (_39232_, _39231_, _29122_);
  nand (_39233_, _39232_, _29090_);
  or (_39234_, _39232_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_39235_, _39234_, _29166_);
  and (_39236_, _39235_, _39233_);
  nor (_39237_, _25678_, _25253_);
  and (_39238_, _39003_, _39237_);
  and (_39239_, _39238_, _38993_);
  not (_39240_, _39239_);
  nor (_39241_, _39240_, _38307_);
  and (_39242_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_39243_, _39242_, _39241_);
  and (_39244_, _39243_, _28541_);
  and (_39245_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_39246_, _39245_, rst);
  or (_39247_, _39246_, _39244_);
  or (_35457_, _39247_, _39236_);
  not (_39248_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39249_, _38994_, _39248_);
  nand (_39250_, _38224_, _24906_);
  nor (_39251_, _39250_, _29090_);
  or (_39252_, _39251_, _39249_);
  and (_39253_, _39252_, _29166_);
  and (_39254_, _38994_, _38286_);
  or (_39255_, _39254_, _39249_);
  and (_39256_, _39255_, _28541_);
  nor (_39257_, _28530_, _39248_);
  or (_39258_, _39257_, rst);
  or (_39259_, _39258_, _39256_);
  or (_41059_, _39259_, _39253_);
  or (_39260_, _38219_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39261_, _39260_, _29166_);
  nand (_39262_, _38226_, _29090_);
  and (_39263_, _39262_, _39261_);
  nand (_39264_, _38994_, _38276_);
  or (_39265_, _38994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39266_, _39265_, _28541_);
  and (_39267_, _39266_, _39264_);
  and (_39268_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_39269_, _39268_, rst);
  or (_39270_, _39269_, _39267_);
  or (_41061_, _39270_, _39263_);
  not (_39271_, _31855_);
  nand (_39272_, _38224_, _39271_);
  and (_39273_, _39272_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39274_, _31157_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39275_, _39274_, _31146_);
  and (_39276_, _39275_, _38224_);
  or (_39277_, _39276_, _39273_);
  and (_39278_, _39277_, _29166_);
  nand (_39279_, _38994_, _38269_);
  or (_39280_, _38994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39281_, _39280_, _28541_);
  and (_39282_, _39281_, _39279_);
  and (_39283_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39284_, _39283_, rst);
  or (_39285_, _39284_, _39282_);
  or (_41062_, _39285_, _39278_);
  not (_39286_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_39287_, _38225_, _39286_);
  nor (_39288_, _31855_, _39286_);
  or (_39289_, _39288_, _31844_);
  and (_39290_, _39289_, _38224_);
  or (_39291_, _39290_, _39287_);
  and (_39292_, _39291_, _29166_);
  nand (_39293_, _38994_, _38261_);
  or (_39294_, _38994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39295_, _39294_, _28541_);
  and (_39296_, _39295_, _39293_);
  nor (_39297_, _28530_, _39286_);
  or (_39298_, _39297_, rst);
  or (_39299_, _39298_, _39296_);
  or (_41064_, _39299_, _39292_);
  not (_39300_, _38224_);
  or (_39301_, _39300_, _32606_);
  and (_39302_, _39301_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39303_, _32595_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39304_, _39303_, _32639_);
  and (_39305_, _39304_, _38224_);
  or (_39306_, _39305_, _39302_);
  and (_39307_, _39306_, _29166_);
  nand (_39308_, _38994_, _38253_);
  or (_39309_, _38994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39310_, _39309_, _28541_);
  and (_39311_, _39310_, _39308_);
  and (_39312_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39313_, _39312_, rst);
  or (_39314_, _39313_, _39311_);
  or (_41066_, _39314_, _39307_);
  and (_39315_, _38224_, _33401_);
  nand (_39316_, _39315_, _29090_);
  or (_39317_, _39315_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39318_, _39317_, _29166_);
  and (_39319_, _39318_, _39316_);
  nand (_39320_, _38994_, _38246_);
  or (_39321_, _38994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39322_, _39321_, _28541_);
  and (_39323_, _39322_, _39320_);
  and (_39324_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39325_, _39324_, rst);
  or (_39326_, _39325_, _39323_);
  or (_41068_, _39326_, _39319_);
  and (_39327_, _38224_, _34130_);
  nand (_39328_, _39327_, _29090_);
  or (_39329_, _39327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39330_, _39329_, _29166_);
  and (_39331_, _39330_, _39328_);
  nand (_39332_, _38994_, _38239_);
  or (_39333_, _38994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39334_, _39333_, _28541_);
  and (_39335_, _39334_, _39332_);
  and (_39336_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39337_, _39336_, rst);
  or (_39338_, _39337_, _39335_);
  or (_41069_, _39338_, _39331_);
  nand (_39339_, _39059_, _29090_);
  or (_39340_, _39059_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39341_, _39340_, _29166_);
  and (_39342_, _39341_, _39339_);
  and (_39343_, _39059_, _38286_);
  and (_39344_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_39345_, _39344_, _39343_);
  and (_39346_, _39345_, _28541_);
  and (_39347_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_39348_, _39347_, rst);
  or (_39349_, _39348_, _39346_);
  or (_41071_, _39349_, _39342_);
  and (_39350_, _39004_, _38217_);
  nand (_39351_, _39350_, _29090_);
  or (_39352_, _39350_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39353_, _39352_, _29166_);
  and (_39354_, _39353_, _39351_);
  nor (_39355_, _39070_, _38276_);
  and (_39356_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39357_, _39356_, _39355_);
  and (_39358_, _39357_, _28541_);
  and (_39359_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39360_, _39359_, rst);
  or (_39361_, _39360_, _39358_);
  or (_41073_, _39361_, _39354_);
  and (_39362_, _39004_, _31124_);
  nand (_39363_, _39362_, _29090_);
  or (_39364_, _39362_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39365_, _39364_, _29166_);
  and (_39366_, _39365_, _39363_);
  nor (_39367_, _39070_, _38269_);
  and (_39368_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39369_, _39368_, _39367_);
  and (_39370_, _39369_, _28541_);
  and (_39371_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39372_, _39371_, rst);
  or (_39373_, _39372_, _39370_);
  or (_41075_, _39373_, _39366_);
  and (_39374_, _39004_, _31822_);
  nand (_39375_, _39374_, _29090_);
  or (_39376_, _39374_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39377_, _39376_, _29166_);
  and (_39378_, _39377_, _39375_);
  nor (_39379_, _39070_, _38261_);
  and (_39380_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39381_, _39380_, _39379_);
  and (_39382_, _39381_, _28541_);
  and (_39383_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39384_, _39383_, rst);
  or (_39385_, _39384_, _39382_);
  or (_41076_, _39385_, _39378_);
  and (_39386_, _39004_, _32584_);
  nand (_39387_, _39386_, _29090_);
  or (_39388_, _39386_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39389_, _39388_, _29166_);
  and (_39390_, _39389_, _39387_);
  nor (_39391_, _39070_, _38253_);
  and (_39392_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39393_, _39392_, _39391_);
  and (_39394_, _39393_, _28541_);
  and (_39395_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39396_, _39395_, rst);
  or (_39397_, _39396_, _39394_);
  or (_41078_, _39397_, _39390_);
  and (_39398_, _39004_, _33401_);
  nand (_39399_, _39398_, _29090_);
  or (_39400_, _39398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39401_, _39400_, _29166_);
  and (_39402_, _39401_, _39399_);
  nor (_39403_, _39070_, _38246_);
  and (_39404_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39405_, _39404_, _39403_);
  and (_39406_, _39405_, _28541_);
  and (_39407_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39408_, _39407_, rst);
  or (_39409_, _39408_, _39406_);
  or (_41080_, _39409_, _39402_);
  and (_39410_, _39004_, _34130_);
  nand (_39411_, _39410_, _29090_);
  or (_39412_, _39410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39413_, _39412_, _29166_);
  and (_39414_, _39413_, _39411_);
  nor (_39415_, _39070_, _38239_);
  and (_39416_, _39070_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39417_, _39416_, _39415_);
  and (_39418_, _39417_, _28541_);
  and (_39419_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39420_, _39419_, rst);
  or (_39421_, _39420_, _39418_);
  or (_41082_, _39421_, _39414_);
  nand (_39422_, _39222_, _29090_);
  or (_39423_, _39222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39424_, _39423_, _29166_);
  and (_39425_, _39424_, _39422_);
  and (_39426_, _39222_, _38286_);
  and (_39427_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_39428_, _39427_, _39426_);
  and (_39432_, _39428_, _28541_);
  and (_39435_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_39436_, _39435_, rst);
  or (_39437_, _39436_, _39432_);
  or (_41083_, _39437_, _39425_);
  and (_39438_, _39190_, _38217_);
  nand (_39439_, _39438_, _29090_);
  or (_39440_, _39438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39441_, _39440_, _29166_);
  and (_39442_, _39441_, _39439_);
  nor (_39443_, _39223_, _38276_);
  and (_39444_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39445_, _39444_, _39443_);
  and (_39446_, _39445_, _28541_);
  and (_39447_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39448_, _39447_, rst);
  or (_39449_, _39448_, _39446_);
  or (_41085_, _39449_, _39442_);
  and (_39450_, _39190_, _31124_);
  nand (_39451_, _39450_, _29090_);
  or (_39452_, _39450_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39453_, _39452_, _29166_);
  and (_39454_, _39453_, _39451_);
  nor (_39455_, _39223_, _38269_);
  and (_39456_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39457_, _39456_, _39455_);
  and (_39458_, _39457_, _28541_);
  and (_39459_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39460_, _39459_, rst);
  or (_39461_, _39460_, _39458_);
  or (_41087_, _39461_, _39454_);
  and (_39477_, _39190_, _31822_);
  nand (_39488_, _39477_, _29090_);
  or (_39492_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39493_, _39492_, _29166_);
  and (_39494_, _39493_, _39488_);
  nor (_39495_, _39223_, _38261_);
  and (_39496_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39497_, _39496_, _39495_);
  and (_39498_, _39497_, _28541_);
  and (_39499_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39500_, _39499_, rst);
  or (_39501_, _39500_, _39498_);
  or (_41089_, _39501_, _39494_);
  and (_39502_, _39190_, _32584_);
  nand (_39503_, _39502_, _29090_);
  or (_39504_, _39502_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39505_, _39504_, _29166_);
  and (_39506_, _39505_, _39503_);
  nor (_39507_, _39223_, _38253_);
  and (_39508_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39509_, _39508_, _39507_);
  and (_39510_, _39509_, _28541_);
  and (_39511_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39512_, _39511_, rst);
  or (_39513_, _39512_, _39510_);
  or (_41090_, _39513_, _39506_);
  and (_39514_, _39190_, _33401_);
  nand (_39515_, _39514_, _29090_);
  or (_39516_, _39514_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39517_, _39516_, _29166_);
  and (_39518_, _39517_, _39515_);
  nor (_39519_, _39223_, _38246_);
  and (_39520_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39525_, _39520_, _39519_);
  and (_39526_, _39525_, _28541_);
  and (_39527_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39528_, _39527_, rst);
  or (_39529_, _39528_, _39526_);
  or (_41092_, _39529_, _39518_);
  and (_39530_, _39190_, _34130_);
  nand (_39531_, _39530_, _29090_);
  or (_39532_, _39530_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39533_, _39532_, _29166_);
  and (_39534_, _39533_, _39531_);
  nor (_39535_, _39223_, _38239_);
  and (_39536_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39537_, _39536_, _39535_);
  and (_39538_, _39537_, _28541_);
  and (_39539_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39540_, _39539_, rst);
  or (_39541_, _39540_, _39538_);
  or (_41094_, _39541_, _39534_);
  and (_39542_, _39231_, _24906_);
  nand (_39543_, _39542_, _29090_);
  or (_39544_, _39542_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39545_, _39544_, _29166_);
  and (_39546_, _39545_, _39543_);
  and (_39547_, _39239_, _38286_);
  and (_39548_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_39549_, _39548_, _39547_);
  and (_39550_, _39549_, _28541_);
  and (_39551_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_39552_, _39551_, rst);
  or (_39553_, _39552_, _39550_);
  or (_41095_, _39553_, _39546_);
  and (_39554_, _39231_, _38217_);
  nand (_39555_, _39554_, _29090_);
  or (_39556_, _39554_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39557_, _39556_, _29166_);
  and (_39558_, _39557_, _39555_);
  nor (_39559_, _39240_, _38276_);
  and (_39560_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39561_, _39560_, _39559_);
  and (_39562_, _39561_, _28541_);
  and (_39563_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39564_, _39563_, rst);
  or (_39565_, _39564_, _39562_);
  or (_41097_, _39565_, _39558_);
  and (_39566_, _39231_, _31124_);
  nand (_39567_, _39566_, _29090_);
  or (_39568_, _39566_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39569_, _39568_, _29166_);
  and (_39570_, _39569_, _39567_);
  nor (_39571_, _39240_, _38269_);
  and (_39572_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39573_, _39572_, _39571_);
  and (_39574_, _39573_, _28541_);
  and (_39575_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39576_, _39575_, rst);
  or (_39577_, _39576_, _39574_);
  or (_41099_, _39577_, _39570_);
  and (_39578_, _39231_, _31822_);
  nand (_39579_, _39578_, _29090_);
  or (_39580_, _39578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39581_, _39580_, _29166_);
  and (_39582_, _39581_, _39579_);
  nor (_39583_, _39240_, _38261_);
  and (_39584_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39585_, _39584_, _39583_);
  and (_39588_, _39585_, _28541_);
  and (_39594_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39595_, _39594_, rst);
  or (_39596_, _39595_, _39588_);
  or (_41101_, _39596_, _39582_);
  and (_39597_, _39231_, _32584_);
  nand (_39598_, _39597_, _29090_);
  or (_39599_, _39597_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39600_, _39599_, _29166_);
  and (_39601_, _39600_, _39598_);
  nor (_39602_, _39240_, _38253_);
  and (_39603_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39604_, _39603_, _39602_);
  and (_39605_, _39604_, _28541_);
  and (_39606_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39607_, _39606_, rst);
  or (_39608_, _39607_, _39605_);
  or (_41103_, _39608_, _39601_);
  and (_39609_, _39231_, _33401_);
  nand (_39610_, _39609_, _29090_);
  or (_39611_, _39609_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39612_, _39611_, _29166_);
  and (_39613_, _39612_, _39610_);
  nor (_39614_, _39240_, _38246_);
  and (_39615_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39616_, _39615_, _39614_);
  and (_39617_, _39616_, _28541_);
  and (_39618_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39619_, _39618_, rst);
  or (_39620_, _39619_, _39617_);
  or (_41104_, _39620_, _39613_);
  and (_39621_, _39231_, _34130_);
  nand (_39622_, _39621_, _29090_);
  or (_39623_, _39621_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39624_, _39623_, _29166_);
  and (_39625_, _39624_, _39622_);
  nor (_39626_, _39240_, _38239_);
  and (_39627_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39628_, _39627_, _39626_);
  and (_39629_, _39628_, _28541_);
  and (_39630_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39631_, _39630_, rst);
  or (_39632_, _39631_, _39629_);
  or (_41106_, _39632_, _39625_);
  nor (_39633_, _25678_, _25548_);
  and (_39634_, _39633_, _39168_);
  and (_39635_, _39634_, _38761_);
  and (_39637_, _39635_, _29122_);
  nand (_39641_, _39637_, _29090_);
  not (_39642_, _25548_);
  and (_39643_, _38701_, _39642_);
  and (_39644_, _39643_, _39238_);
  not (_39645_, _39644_);
  or (_39646_, _39637_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_39647_, _39646_, _39645_);
  and (_39648_, _39647_, _39641_);
  nor (_39649_, _39645_, _38307_);
  or (_39650_, _39649_, _39648_);
  and (_41597_, _39650_, _41654_);
  and (_39651_, _25678_, _39642_);
  and (_39652_, _39651_, _38761_);
  and (_39653_, _39652_, _39168_);
  and (_39654_, _39653_, _29122_);
  nand (_39658_, _39654_, _29090_);
  and (_39665_, _39643_, _39221_);
  not (_39666_, _39665_);
  or (_39667_, _39654_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_39668_, _39667_, _39666_);
  and (_39669_, _39668_, _39658_);
  nor (_39670_, _39666_, _38307_);
  or (_39671_, _39670_, _39669_);
  and (_41599_, _39671_, _41654_);
  or (_39672_, _24895_, _31113_);
  and (_39673_, _39672_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39674_, _39673_, _38870_);
  and (_39675_, _39652_, _38214_);
  and (_39676_, _39675_, _39674_);
  and (_39677_, _39643_, _38216_);
  nand (_39678_, _39675_, _24884_);
  and (_39679_, _39678_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39680_, _39679_, _39677_);
  or (_39681_, _39680_, _39676_);
  nand (_39682_, _39677_, _38239_);
  and (_39683_, _39682_, _41654_);
  and (_41601_, _39683_, _39681_);
  and (_39684_, _29166_, _29112_);
  nor (_39685_, _24645_, _25548_);
  and (_39686_, _39685_, _38216_);
  and (_39687_, _39686_, _39684_);
  nand (_39688_, _39687_, _29090_);
  not (_39689_, _39677_);
  not (_39690_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_39691_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_39692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_39693_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _39692_);
  and (_39694_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39695_, _39694_, _39693_);
  nor (_39696_, _39695_, _39691_);
  or (_39697_, _39696_, _39690_);
  and (_39698_, _39692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_39699_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_39700_, _39699_, _39698_);
  nor (_39701_, _39700_, _39691_);
  and (_39702_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _39692_);
  and (_39703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39704_, _39703_, _39702_);
  nand (_39705_, _39704_, _39701_);
  or (_39706_, _39705_, _39697_);
  and (_39707_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_39708_, _39707_, _39687_);
  and (_39709_, _39708_, _39689_);
  and (_39710_, _39709_, _39688_);
  nor (_39711_, _39689_, _38307_);
  or (_39712_, _39711_, _39710_);
  and (_41604_, _39712_, _41654_);
  and (_39713_, _29166_, _30414_);
  and (_39714_, _39713_, _39686_);
  nand (_39715_, _39714_, _29090_);
  nor (_39716_, _39704_, _39691_);
  nand (_39717_, _39716_, _39700_);
  or (_39718_, _39717_, _39697_);
  and (_39719_, _39718_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_39720_, _39719_, _39714_);
  and (_39721_, _39720_, _39689_);
  and (_39722_, _39721_, _39715_);
  nor (_39723_, _39689_, _38246_);
  or (_39724_, _39723_, _39722_);
  and (_41606_, _39724_, _41654_);
  nor (_39725_, _29101_, _25548_);
  and (_39726_, _39725_, _38216_);
  and (_39727_, _39726_, _39713_);
  nand (_39728_, _39727_, _29090_);
  not (_39729_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_39730_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _39729_);
  nand (_39731_, _39696_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_39732_, _39716_, _39701_);
  or (_39733_, _39732_, _39731_);
  and (_39734_, _39733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_39735_, _39734_, _39730_);
  or (_39736_, _39735_, _39727_);
  and (_39737_, _39736_, _39689_);
  and (_39738_, _39737_, _39728_);
  nor (_39739_, _39689_, _38276_);
  or (_39740_, _39739_, _39738_);
  and (_41608_, _39740_, _41654_);
  and (_39741_, _39726_, _39684_);
  nand (_39742_, _39741_, _29090_);
  and (_39743_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_39744_, _39731_, _39717_);
  and (_39745_, _39744_, _39743_);
  or (_39746_, _39745_, _39741_);
  and (_39747_, _39746_, _39689_);
  and (_39748_, _39747_, _39742_);
  nor (_39749_, _39689_, _38261_);
  or (_39750_, _39749_, _39748_);
  and (_41610_, _39750_, _41654_);
  and (_39751_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_39752_, _39751_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_39753_, _39752_);
  and (_39754_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_39755_, _39754_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_39756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_39757_, _39756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_39758_, _39757_, _39755_);
  and (_39759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_39760_, _39759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  not (_39761_, _39760_);
  and (_39762_, _39761_, _39758_);
  and (_39763_, _39762_, _39753_);
  not (_39764_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_39765_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_39766_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _39692_);
  or (_39767_, _39766_, _39765_);
  nor (_39768_, _39767_, _39764_);
  nor (_39769_, _39768_, _39691_);
  nor (_39770_, _39769_, _39763_);
  and (_39771_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_39772_, _39771_, _39692_);
  and (_39773_, _39772_, _39770_);
  and (_39774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _39691_);
  not (_39775_, _39774_);
  not (_39776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_39777_, _39754_, _39776_);
  not (_39778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_39779_, _39756_, _39778_);
  nor (_39780_, _39779_, _39777_);
  not (_39781_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_39782_, _39759_, _39781_);
  not (_39783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_39784_, _39751_, _39783_);
  nor (_39785_, _39784_, _39782_);
  and (_39786_, _39785_, _39780_);
  nor (_39787_, _39786_, _39775_);
  nand (_39788_, _39787_, _39772_);
  and (_39789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41654_);
  nand (_39790_, _39789_, _39788_);
  nor (_41641_, _39790_, _39773_);
  nor (_39791_, _39771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_39792_, _39791_);
  nor (_39793_, _39787_, _39770_);
  nor (_39794_, _39793_, _39792_);
  nand (_39795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41654_);
  nor (_41643_, _39795_, _39794_);
  and (_39796_, _39752_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_39797_, _39758_);
  or (_39798_, _39797_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_39799_, _39798_, _39796_);
  or (_39800_, _39762_, _39698_);
  and (_39801_, _39800_, _39799_);
  and (_39802_, _39801_, _39770_);
  or (_39803_, _39802_, _39771_);
  and (_39804_, _39793_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_39805_, _39770_);
  and (_39806_, _39787_, _39805_);
  and (_39807_, _39784_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_39808_, _39807_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_39809_, _39780_);
  and (_39810_, _39782_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39811_, _39810_, _39809_);
  and (_39812_, _39811_, _39808_);
  and (_39813_, _39809_, _39698_);
  or (_39814_, _39813_, _39812_);
  and (_39815_, _39814_, _39806_);
  or (_39816_, _39815_, _39804_);
  or (_39817_, _39816_, _39803_);
  not (_39818_, _39771_);
  or (_39819_, _39818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_39820_, _39819_, _41654_);
  and (_41645_, _39820_, _39817_);
  and (_39821_, _39752_, _39692_);
  or (_39822_, _39797_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_39823_, _39822_, _39821_);
  or (_39824_, _39762_, _39699_);
  and (_39825_, _39824_, _39823_);
  and (_39826_, _39825_, _39770_);
  or (_39827_, _39826_, _39771_);
  and (_39828_, _39793_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_39829_, _39784_, _39692_);
  or (_39830_, _39829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_39831_, _39782_, _39692_);
  nor (_39832_, _39831_, _39809_);
  and (_39833_, _39832_, _39830_);
  and (_39834_, _39809_, _39699_);
  or (_39835_, _39834_, _39833_);
  and (_39836_, _39835_, _39806_);
  or (_39837_, _39836_, _39828_);
  or (_39838_, _39837_, _39827_);
  or (_39839_, _39818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_39840_, _39839_, _41654_);
  and (_41647_, _39840_, _39838_);
  nand (_39841_, _39793_, _39691_);
  nor (_39842_, _39692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_39843_, _39842_, _39771_);
  and (_39844_, _39843_, _41654_);
  and (_41649_, _39844_, _39841_);
  and (_39845_, _39793_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_39846_, _39692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_39847_, _39846_, _39842_);
  nor (_39848_, _39847_, _39805_);
  or (_39849_, _39848_, _39771_);
  or (_39850_, _39849_, _39845_);
  or (_39851_, _39847_, _39818_);
  and (_39852_, _39851_, _41654_);
  and (_41651_, _39852_, _39850_);
  and (_39853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41654_);
  and (_41652_, _39853_, _39771_);
  nor (_39854_, _39793_, _39771_);
  and (_39855_, _39771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_39856_, _39855_, _39854_);
  and (_42571_, _39856_, _41654_);
  and (_39857_, _39771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_39858_, _39857_, _39854_);
  and (_42573_, _39858_, _41654_);
  and (_39859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _41654_);
  and (_42574_, _39859_, _39771_);
  not (_39860_, _39777_);
  nor (_39861_, _39784_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_39862_, _39861_, _39782_);
  or (_39863_, _39862_, _39779_);
  and (_39864_, _39863_, _39860_);
  and (_39865_, _39864_, _39806_);
  not (_39866_, _39755_);
  or (_39867_, _39752_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39868_, _39867_, _39761_);
  or (_39869_, _39868_, _39757_);
  and (_39870_, _39869_, _39866_);
  and (_39871_, _39870_, _39770_);
  or (_39872_, _39871_, _39771_);
  or (_39873_, _39872_, _39865_);
  or (_39874_, _39818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39875_, _39874_, _41654_);
  and (_42576_, _39875_, _39873_);
  nand (_39876_, _39780_, _39774_);
  nor (_39877_, _39876_, _39785_);
  or (_39878_, _39877_, _39770_);
  nand (_39879_, _39770_, _39797_);
  and (_39880_, _39879_, _39878_);
  or (_39881_, _39880_, _39771_);
  or (_39882_, _39818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39883_, _39882_, _41654_);
  and (_42578_, _39883_, _39881_);
  and (_39884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _41654_);
  and (_42580_, _39884_, _39771_);
  and (_39885_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _41654_);
  and (_42582_, _39885_, _39771_);
  nand (_39886_, _39793_, _39791_);
  nor (_39887_, _39771_, _39770_);
  or (_39888_, _39887_, _39692_);
  and (_39889_, _39888_, _41654_);
  and (_42584_, _39889_, _39886_);
  not (_39890_, _39854_);
  and (_39891_, _39890_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_39892_, _39821_);
  and (_39893_, _39892_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_39894_, _39760_, _39692_);
  or (_39895_, _39894_, _39757_);
  or (_39896_, _39895_, _39893_);
  not (_39897_, _39757_);
  or (_39898_, _39897_, _39694_);
  and (_39899_, _39898_, _39896_);
  or (_39900_, _39899_, _39755_);
  or (_39901_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _39692_);
  or (_39902_, _39901_, _39866_);
  and (_39903_, _39902_, _39770_);
  and (_39904_, _39903_, _39900_);
  not (_39905_, _39829_);
  and (_39906_, _39905_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_39907_, _39831_, _39779_);
  or (_39908_, _39907_, _39906_);
  not (_39909_, _39779_);
  or (_39910_, _39909_, _39694_);
  and (_39911_, _39910_, _39860_);
  and (_39912_, _39911_, _39908_);
  and (_39913_, _39901_, _39777_);
  or (_39914_, _39913_, _39912_);
  and (_39915_, _39914_, _39806_);
  or (_39916_, _39915_, _39904_);
  and (_39917_, _39916_, _39818_);
  or (_39918_, _39917_, _39891_);
  and (_42586_, _39918_, _41654_);
  and (_39919_, _39890_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_39920_, _39892_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_39921_, _39920_, _39895_);
  or (_39922_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _39692_);
  or (_39923_, _39922_, _39897_);
  and (_39924_, _39923_, _39866_);
  and (_39925_, _39924_, _39921_);
  and (_39926_, _39755_, _39703_);
  or (_39927_, _39926_, _39925_);
  and (_39928_, _39927_, _39770_);
  and (_39929_, _39905_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_39930_, _39929_, _39907_);
  or (_39931_, _39922_, _39909_);
  and (_39932_, _39931_, _39860_);
  and (_39933_, _39932_, _39930_);
  and (_39934_, _39777_, _39703_);
  or (_39935_, _39934_, _39933_);
  and (_39936_, _39935_, _39806_);
  or (_39937_, _39936_, _39928_);
  and (_39938_, _39937_, _39818_);
  or (_39939_, _39938_, _39919_);
  and (_42587_, _39939_, _41654_);
  and (_39940_, _39890_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_39941_, _39796_);
  and (_39942_, _39941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_39943_, _39760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_39944_, _39943_, _39757_);
  or (_39945_, _39944_, _39942_);
  or (_39946_, _39897_, _39693_);
  and (_39947_, _39946_, _39945_);
  or (_39948_, _39947_, _39755_);
  or (_39949_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_39950_, _39949_, _39866_);
  and (_39951_, _39950_, _39770_);
  and (_39952_, _39951_, _39948_);
  not (_39953_, _39807_);
  and (_39954_, _39953_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_39955_, _39810_, _39779_);
  or (_39956_, _39955_, _39954_);
  or (_39957_, _39909_, _39693_);
  and (_39958_, _39957_, _39860_);
  and (_39959_, _39958_, _39956_);
  and (_39960_, _39949_, _39777_);
  or (_39961_, _39960_, _39959_);
  and (_39962_, _39961_, _39806_);
  or (_39963_, _39962_, _39952_);
  and (_39964_, _39963_, _39818_);
  or (_39965_, _39964_, _39940_);
  and (_42589_, _39965_, _41654_);
  and (_39966_, _39890_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_39967_, _39941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_39968_, _39967_, _39944_);
  or (_39969_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_39970_, _39969_, _39897_);
  and (_39971_, _39970_, _39866_);
  and (_39972_, _39971_, _39968_);
  and (_39973_, _39755_, _39702_);
  or (_39974_, _39973_, _39972_);
  and (_39975_, _39974_, _39770_);
  and (_39976_, _39953_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_39977_, _39976_, _39955_);
  or (_39978_, _39969_, _39909_);
  and (_39979_, _39978_, _39860_);
  and (_39980_, _39979_, _39977_);
  and (_39981_, _39777_, _39702_);
  or (_39982_, _39981_, _39980_);
  and (_39983_, _39982_, _39806_);
  or (_39984_, _39983_, _39975_);
  and (_39985_, _39984_, _39818_);
  or (_39986_, _39985_, _39966_);
  and (_42591_, _39986_, _41654_);
  and (_39987_, _39791_, _39770_);
  nand (_39988_, _39791_, _39787_);
  and (_39989_, _39988_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_39990_, _39989_, _39987_);
  and (_42593_, _39990_, _41654_);
  and (_39991_, _39788_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_39992_, _39991_, _39773_);
  and (_42595_, _39992_, _41654_);
  and (_39993_, _39675_, _24906_);
  or (_39994_, _39993_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_39995_, _39994_, _39689_);
  nand (_39996_, _39993_, _29090_);
  and (_39997_, _39996_, _39995_);
  and (_39998_, _39677_, _38286_);
  or (_39999_, _39998_, _39997_);
  and (_42597_, _39999_, _41654_);
  and (_40000_, _39675_, _31124_);
  nand (_40001_, _40000_, _29090_);
  or (_40002_, _40000_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_40003_, _40002_, _39689_);
  and (_40004_, _40003_, _40001_);
  nor (_40005_, _39689_, _38269_);
  or (_40006_, _40005_, _40004_);
  and (_42599_, _40006_, _41654_);
  and (_40007_, _39675_, _32584_);
  nand (_40008_, _40007_, _29090_);
  or (_40009_, _40007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_40010_, _40009_, _39689_);
  and (_40011_, _40010_, _40008_);
  nor (_40012_, _39689_, _38253_);
  or (_40013_, _40012_, _40011_);
  and (_42601_, _40013_, _41654_);
  and (_40014_, _39653_, _24906_);
  nand (_40015_, _40014_, _29090_);
  or (_40016_, _40014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40017_, _40016_, _39666_);
  and (_40018_, _40017_, _40015_);
  and (_40019_, _39665_, _38286_);
  or (_40020_, _40019_, _40018_);
  and (_42603_, _40020_, _41654_);
  and (_40021_, _39653_, _38217_);
  nand (_40022_, _40021_, _29090_);
  or (_40023_, _40021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40024_, _40023_, _39666_);
  and (_40025_, _40024_, _40022_);
  nor (_40026_, _39666_, _38276_);
  or (_40027_, _40026_, _40025_);
  and (_42604_, _40027_, _41654_);
  and (_40028_, _31157_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40029_, _40028_, _31146_);
  and (_40030_, _40029_, _39653_);
  nand (_40031_, _39653_, _39271_);
  and (_40032_, _40031_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40033_, _40032_, _39665_);
  or (_40034_, _40033_, _40030_);
  nand (_40035_, _39665_, _38269_);
  and (_40036_, _40035_, _41654_);
  and (_42606_, _40036_, _40034_);
  and (_40037_, _39653_, _31822_);
  nand (_40038_, _40037_, _29090_);
  or (_40039_, _40037_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40040_, _40039_, _39666_);
  and (_40041_, _40040_, _40038_);
  nor (_40042_, _39666_, _38261_);
  or (_40043_, _40042_, _40041_);
  and (_42608_, _40043_, _41654_);
  and (_40044_, _39653_, _32584_);
  nand (_40045_, _40044_, _29090_);
  or (_40046_, _40044_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_40047_, _40046_, _39666_);
  and (_40048_, _40047_, _40045_);
  nor (_40049_, _39666_, _38253_);
  or (_40050_, _40049_, _40048_);
  and (_42610_, _40050_, _41654_);
  and (_40051_, _39653_, _33401_);
  nand (_40052_, _40051_, _29090_);
  or (_40053_, _40051_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_40054_, _40053_, _39666_);
  and (_40055_, _40054_, _40052_);
  nor (_40056_, _39666_, _38246_);
  or (_40057_, _40056_, _40055_);
  and (_42612_, _40057_, _41654_);
  and (_40058_, _39653_, _34130_);
  nand (_40059_, _40058_, _29090_);
  or (_40060_, _40058_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_40061_, _40060_, _39666_);
  and (_40062_, _40061_, _40059_);
  nor (_40063_, _39666_, _38239_);
  or (_40064_, _40063_, _40062_);
  and (_42614_, _40064_, _41654_);
  and (_40065_, _39635_, _24906_);
  nand (_40066_, _40065_, _29090_);
  or (_40067_, _40065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40068_, _40067_, _39645_);
  and (_40069_, _40068_, _40066_);
  and (_40070_, _39644_, _38286_);
  or (_40071_, _40070_, _40069_);
  and (_42616_, _40071_, _41654_);
  and (_40072_, _39635_, _38217_);
  nand (_40073_, _40072_, _29090_);
  or (_40074_, _40072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40075_, _40074_, _39645_);
  and (_40076_, _40075_, _40073_);
  nor (_40077_, _39645_, _38276_);
  or (_40078_, _40077_, _40076_);
  and (_42618_, _40078_, _41654_);
  and (_40079_, _31157_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40080_, _40079_, _31146_);
  and (_40081_, _40080_, _39635_);
  nand (_40082_, _39635_, _39271_);
  and (_40083_, _40082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40084_, _40083_, _39644_);
  or (_40085_, _40084_, _40081_);
  nand (_40086_, _39644_, _38269_);
  and (_40087_, _40086_, _41654_);
  and (_42620_, _40087_, _40085_);
  and (_40088_, _39635_, _31822_);
  nand (_40089_, _40088_, _29090_);
  or (_40090_, _40088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40091_, _40090_, _39645_);
  and (_40092_, _40091_, _40089_);
  nor (_40093_, _39645_, _38261_);
  or (_40094_, _40093_, _40092_);
  and (_42622_, _40094_, _41654_);
  and (_40095_, _39635_, _32584_);
  nand (_40096_, _40095_, _29090_);
  or (_40097_, _40095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40098_, _40097_, _39645_);
  and (_40099_, _40098_, _40096_);
  nor (_40100_, _39645_, _38253_);
  or (_40101_, _40100_, _40099_);
  and (_42624_, _40101_, _41654_);
  and (_40102_, _39635_, _33401_);
  nand (_40103_, _40102_, _29090_);
  or (_40104_, _40102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40105_, _40104_, _39645_);
  and (_40106_, _40105_, _40103_);
  nor (_40107_, _39645_, _38246_);
  or (_40108_, _40107_, _40106_);
  and (_42626_, _40108_, _41654_);
  and (_40109_, _39635_, _34130_);
  nand (_40110_, _40109_, _29090_);
  or (_40111_, _40109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_40112_, _40111_, _39645_);
  and (_40113_, _40112_, _40110_);
  nor (_40114_, _39645_, _38239_);
  or (_40115_, _40114_, _40113_);
  and (_42628_, _40115_, _41654_);
  and (_40116_, _38212_, _38198_);
  and (_40117_, _38309_, _40116_);
  not (_40118_, _40117_);
  not (_40119_, _37255_);
  nor (_40120_, _38197_, _40119_);
  not (_40121_, _34293_);
  and (_40122_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_40123_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_40124_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_40125_, _40124_, _40123_);
  and (_40126_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_40127_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_40128_, _40127_, _40126_);
  and (_40129_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_40130_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_40131_, _40130_, _40129_);
  and (_40132_, _40131_, _40128_);
  and (_40133_, _40132_, _40125_);
  nor (_40134_, _34347_, _40121_);
  not (_40135_, _40134_);
  nor (_40136_, _40135_, _40133_);
  nor (_40137_, _40136_, _40122_);
  not (_40138_, _40137_);
  and (_40139_, _40138_, _40120_);
  not (_40140_, _40139_);
  not (_40141_, _38212_);
  and (_40142_, _38197_, _40119_);
  and (_40143_, _36720_, _30403_);
  nor (_40144_, _36720_, _30403_);
  not (_40145_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_40146_, _28508_, _40145_);
  and (_40147_, _40146_, _31157_);
  nand (_40148_, _40147_, _25395_);
  or (_40149_, _40148_, _40144_);
  nor (_40150_, _40149_, _40143_);
  nor (_40151_, _38705_, _38834_);
  nor (_40152_, _40151_, _38840_);
  and (_40153_, _40152_, _39642_);
  nor (_40154_, _40152_, _39642_);
  nor (_40155_, _40154_, _40153_);
  and (_40156_, _40155_, _40150_);
  nor (_40157_, _40152_, _36862_);
  and (_40158_, _40157_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_40159_, _40152_, _36862_);
  and (_40160_, _40159_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_40161_, _40160_, _40158_);
  nor (_40162_, _40152_, _36720_);
  and (_40163_, _40162_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_40164_, _40152_, _36720_);
  and (_40165_, _40164_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_40166_, _40165_, _40163_);
  and (_40167_, _40166_, _40161_);
  nor (_40168_, _40167_, _40156_);
  not (_40169_, _38307_);
  and (_40170_, _40156_, _40169_);
  nor (_40171_, _40170_, _40168_);
  not (_40172_, _40171_);
  and (_40173_, _40172_, _40142_);
  nor (_40174_, _40173_, _40141_);
  and (_40175_, _40174_, _40140_);
  and (_40176_, _40175_, _40118_);
  not (_40177_, _37920_);
  and (_40178_, _40177_, _37601_);
  nor (_40179_, _37645_, _37843_);
  nor (_40180_, _37887_, _37832_);
  and (_40181_, _40180_, _40179_);
  and (_40182_, _38030_, _37766_);
  and (_40183_, _40182_, _40181_);
  and (_40184_, _40183_, _40178_);
  nor (_40185_, _40184_, _34249_);
  and (_40186_, _37997_, _36742_);
  nor (_40187_, _38189_, _40186_);
  nor (_40188_, _40187_, _38186_);
  nor (_40189_, _40188_, _40185_);
  not (_40190_, _40189_);
  and (_40191_, _40190_, _40176_);
  and (_40192_, _40120_, _38212_);
  and (_40193_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_40194_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_40195_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_40196_, _40195_, _40194_);
  and (_40197_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_40198_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_40199_, _40198_, _40197_);
  and (_40200_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_40201_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_40202_, _40201_, _40200_);
  and (_40203_, _40202_, _40199_);
  and (_40204_, _40203_, _40196_);
  nor (_40205_, _40204_, _40135_);
  nor (_40206_, _40205_, _40193_);
  not (_40207_, _40206_);
  and (_40208_, _40207_, _40192_);
  not (_40209_, _40208_);
  and (_40210_, _40141_, _37255_);
  and (_40211_, _40210_, _38197_);
  not (_40212_, _38347_);
  and (_40213_, _40212_, _40116_);
  nor (_40214_, _40213_, _40211_);
  and (_40215_, _40214_, _40209_);
  and (_40216_, _40141_, _38198_);
  and (_40217_, _40142_, _38212_);
  and (_40218_, _40162_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_40219_, _40159_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_40220_, _40219_, _40218_);
  and (_40221_, _40164_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_40222_, _40157_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_40223_, _40222_, _40221_);
  and (_40224_, _40223_, _40220_);
  nor (_40225_, _40224_, _40156_);
  not (_40226_, _38246_);
  and (_40227_, _40156_, _40226_);
  nor (_40228_, _40227_, _40225_);
  not (_40229_, _40228_);
  and (_40230_, _40229_, _40217_);
  nor (_40231_, _40230_, _40216_);
  and (_40232_, _40231_, _40215_);
  not (_40233_, _40232_);
  and (_40234_, _40233_, _40191_);
  and (_40235_, _38212_, _37255_);
  and (_40236_, _40235_, _38197_);
  and (_40237_, _40236_, _37287_);
  and (_40238_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_40239_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_40240_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_40241_, _40240_, _40239_);
  and (_40242_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_40243_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_40244_, _40243_, _40242_);
  and (_40245_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_40246_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_40247_, _40246_, _40245_);
  and (_40248_, _40247_, _40244_);
  and (_40249_, _40248_, _40241_);
  nor (_40250_, _40249_, _40135_);
  nor (_40251_, _40250_, _40238_);
  not (_40252_, _40251_);
  and (_40253_, _40252_, _40192_);
  nor (_40254_, _40253_, _40237_);
  not (_40255_, _38329_);
  and (_40256_, _40255_, _40116_);
  and (_40257_, _40162_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_40258_, _40159_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_40259_, _40258_, _40257_);
  and (_40260_, _40164_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_40261_, _40157_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_40262_, _40261_, _40260_);
  and (_40263_, _40262_, _40259_);
  nor (_40264_, _40263_, _40156_);
  not (_40265_, _40156_);
  nor (_40266_, _40265_, _38269_);
  nor (_40267_, _40266_, _40264_);
  not (_40268_, _40267_);
  and (_40269_, _40268_, _40217_);
  nor (_40270_, _40269_, _40256_);
  and (_40271_, _40270_, _40254_);
  nor (_40272_, _40271_, _40190_);
  nor (_40273_, _40272_, _40234_);
  and (_40274_, _25395_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40275_, _40274_, _38882_);
  nor (_40276_, _24645_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40277_, _40276_, _40275_);
  not (_40278_, _40277_);
  and (_40279_, _40278_, _40273_);
  not (_40280_, _40152_);
  and (_40281_, _40236_, _40280_);
  and (_40282_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_40283_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_40284_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_40285_, _40284_, _40283_);
  and (_40286_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_40287_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_40288_, _40287_, _40286_);
  and (_40289_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_40290_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_40291_, _40290_, _40289_);
  and (_40292_, _40291_, _40288_);
  and (_40293_, _40292_, _40285_);
  nor (_40294_, _40293_, _40135_);
  nor (_40295_, _40294_, _40282_);
  not (_40296_, _40295_);
  and (_40297_, _40296_, _40192_);
  nor (_40298_, _40297_, _40281_);
  not (_40299_, _38335_);
  and (_40300_, _40299_, _40116_);
  not (_40301_, _38261_);
  and (_40302_, _40156_, _40301_);
  and (_40303_, _40162_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_40304_, _40159_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_40305_, _40304_, _40303_);
  and (_40306_, _40164_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_40307_, _40157_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_40308_, _40307_, _40306_);
  and (_40309_, _40308_, _40305_);
  nor (_40310_, _40309_, _40156_);
  nor (_40311_, _40310_, _40302_);
  not (_40312_, _40311_);
  and (_40313_, _40312_, _40217_);
  nor (_40314_, _40313_, _40300_);
  and (_40315_, _40314_, _40298_);
  not (_40316_, _40315_);
  and (_40317_, _40316_, _40191_);
  and (_40318_, _40236_, _36862_);
  and (_40319_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_40320_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_40321_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_40322_, _40321_, _40320_);
  and (_40323_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_40324_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_40325_, _40324_, _40323_);
  and (_40326_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_40327_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_40328_, _40327_, _40326_);
  and (_40329_, _40328_, _40325_);
  and (_40330_, _40329_, _40322_);
  nor (_40331_, _40330_, _40135_);
  nor (_40332_, _40331_, _40319_);
  not (_40333_, _40332_);
  and (_40334_, _40333_, _40192_);
  nor (_40335_, _40334_, _40318_);
  not (_40336_, _38317_);
  and (_40337_, _40336_, _40116_);
  and (_40338_, _40162_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_40339_, _40159_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_40340_, _40339_, _40338_);
  and (_40341_, _40164_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_40342_, _40157_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_40343_, _40342_, _40341_);
  and (_40344_, _40343_, _40340_);
  nor (_40345_, _40344_, _40156_);
  and (_40346_, _40156_, _38286_);
  nor (_40347_, _40346_, _40345_);
  not (_40348_, _40347_);
  and (_40349_, _40348_, _40217_);
  nor (_40350_, _40349_, _40337_);
  and (_40351_, _40350_, _40335_);
  nor (_40352_, _40351_, _40190_);
  nor (_40353_, _40352_, _40317_);
  and (_40354_, _40274_, _39642_);
  nor (_40355_, _24884_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40356_, _40355_, _40354_);
  not (_40357_, _40356_);
  nor (_40358_, _40357_, _40353_);
  nor (_40359_, _40358_, _40279_);
  nor (_40360_, _40278_, _40273_);
  not (_40361_, _40360_);
  and (_40362_, _40157_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_40363_, _40159_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_40364_, _40363_, _40362_);
  and (_40365_, _40162_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_40366_, _40164_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_40367_, _40366_, _40365_);
  and (_40368_, _40367_, _40364_);
  nor (_40369_, _40368_, _40156_);
  not (_40370_, _38239_);
  and (_40371_, _40156_, _40370_);
  nor (_40372_, _40371_, _40369_);
  not (_40373_, _40372_);
  and (_40374_, _40373_, _40217_);
  and (_40375_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_40376_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_40377_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_40378_, _40377_, _40376_);
  and (_40379_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_40380_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_40381_, _40380_, _40379_);
  and (_40382_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_40383_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_40384_, _40383_, _40382_);
  and (_40385_, _40384_, _40381_);
  and (_40386_, _40385_, _40378_);
  nor (_40387_, _40386_, _40135_);
  nor (_40388_, _40387_, _40375_);
  not (_40389_, _40388_);
  and (_40390_, _40389_, _40120_);
  or (_40391_, _40390_, _40210_);
  nor (_40392_, _40391_, _40374_);
  not (_40393_, _38353_);
  and (_40394_, _40393_, _40116_);
  nor (_40395_, _40394_, _40216_);
  and (_40396_, _40395_, _40392_);
  and (_40397_, _40396_, _40191_);
  nor (_40398_, _40316_, _40191_);
  nor (_40399_, _40398_, _40397_);
  nor (_40400_, _40274_, _39642_);
  and (_40401_, _40274_, _25122_);
  nor (_40402_, _40401_, _40400_);
  not (_40403_, _40402_);
  and (_40404_, _40403_, _40399_);
  nor (_40405_, _40403_, _40399_);
  nor (_40406_, _40405_, _40404_);
  and (_40407_, _40406_, _40361_);
  and (_40408_, _38341_, _40116_);
  or (_40409_, _40408_, _40210_);
  and (_40410_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_40411_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_40412_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_40413_, _40412_, _40411_);
  and (_40414_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_40415_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_40416_, _40415_, _40414_);
  and (_40417_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_40418_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_40419_, _40418_, _40417_);
  and (_40420_, _40419_, _40416_);
  and (_40421_, _40420_, _40413_);
  nor (_40422_, _40421_, _40135_);
  nor (_40423_, _40422_, _40410_);
  not (_40424_, _40423_);
  and (_40425_, _40424_, _40192_);
  and (_40426_, _40157_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_40427_, _40159_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_40428_, _40427_, _40426_);
  and (_40429_, _40162_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_40430_, _40164_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  or (_40431_, _40430_, _40429_);
  or (_40432_, _40431_, _40428_);
  and (_40433_, _40432_, _40265_);
  not (_40434_, _38253_);
  and (_40435_, _40156_, _40434_);
  or (_40436_, _40435_, _40433_);
  and (_40437_, _40436_, _40217_);
  or (_40438_, _40437_, _40425_);
  and (_40442_, _38741_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_40448_, _40442_, _38850_);
  and (_40454_, _40448_, _40236_);
  or (_40460_, _40454_, _40438_);
  or (_40466_, _40460_, _40409_);
  and (_40471_, _40466_, _40191_);
  and (_40472_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_40473_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_40474_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_40475_, _40474_, _40473_);
  and (_40476_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_40477_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_40478_, _40477_, _40476_);
  and (_40479_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_40480_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_40481_, _40480_, _40479_);
  and (_40482_, _40481_, _40478_);
  and (_40483_, _40482_, _40475_);
  nor (_40484_, _40483_, _40135_);
  nor (_40485_, _40484_, _40472_);
  not (_40488_, _40485_);
  and (_40492_, _40488_, _40192_);
  and (_40496_, _40162_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_40497_, _40159_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_40498_, _40497_, _40496_);
  and (_40499_, _40164_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_40504_, _40157_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_40509_, _40504_, _40499_);
  and (_40510_, _40509_, _40498_);
  nor (_40511_, _40510_, _40156_);
  and (_40513_, _40156_, _38277_);
  nor (_40519_, _40513_, _40511_);
  not (_40522_, _40519_);
  and (_40523_, _40522_, _40217_);
  nor (_40524_, _40523_, _40492_);
  not (_40529_, _38323_);
  and (_40534_, _40529_, _40116_);
  not (_40535_, _40534_);
  and (_40536_, _40142_, _40141_);
  and (_40538_, _40236_, _36786_);
  nor (_40544_, _40538_, _40536_);
  and (_40547_, _40544_, _40535_);
  and (_40548_, _40547_, _40524_);
  nor (_40549_, _40548_, _40190_);
  nor (_40555_, _40549_, _40471_);
  and (_40559_, _40274_, _25689_);
  nor (_40560_, _24764_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40561_, _40560_, _40559_);
  nand (_40567_, _40561_, _40555_);
  or (_40571_, _40561_, _40555_);
  and (_40572_, _40571_, _40567_);
  not (_40573_, _40572_);
  nor (_40578_, _25395_, _24437_);
  nor (_40583_, _40578_, _28519_);
  not (_40584_, _40583_);
  and (_40585_, _40357_, _40353_);
  nor (_40587_, _40585_, _40584_);
  and (_40593_, _40587_, _40573_);
  and (_40596_, _40593_, _40407_);
  and (_40597_, _40596_, _40359_);
  not (_40598_, _40273_);
  and (_40604_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_40608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_40609_, _40353_, _40608_);
  or (_40610_, _40609_, _40604_);
  and (_40616_, _40610_, _40555_);
  not (_40620_, _40555_);
  not (_40621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_40622_, _40353_, _40621_);
  and (_40627_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_40632_, _40627_, _40622_);
  and (_40633_, _40632_, _40620_);
  or (_40634_, _40633_, _40616_);
  or (_40638_, _40634_, _40598_);
  not (_40644_, _40399_);
  and (_40645_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not (_40646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_40649_, _40353_, _40646_);
  or (_40655_, _40649_, _40645_);
  and (_40657_, _40655_, _40555_);
  not (_40658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_40661_, _40353_, _40658_);
  and (_40667_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_40669_, _40667_, _40661_);
  and (_40670_, _40669_, _40620_);
  or (_40673_, _40670_, _40657_);
  or (_40679_, _40673_, _40273_);
  and (_40680_, _40679_, _40644_);
  and (_40681_, _40680_, _40638_);
  not (_40682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_40683_, _40353_, _40682_);
  or (_40684_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_40685_, _40684_, _40683_);
  and (_40686_, _40685_, _40555_);
  or (_40687_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_40688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_40689_, _40353_, _40688_);
  and (_40690_, _40689_, _40687_);
  and (_40691_, _40690_, _40620_);
  or (_40692_, _40691_, _40686_);
  or (_40693_, _40692_, _40598_);
  not (_40694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_40695_, _40353_, _40694_);
  or (_40696_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_40697_, _40696_, _40695_);
  and (_40698_, _40697_, _40555_);
  or (_40699_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_40700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_40701_, _40353_, _40700_);
  and (_40702_, _40701_, _40699_);
  and (_40703_, _40702_, _40620_);
  or (_40704_, _40703_, _40698_);
  or (_40705_, _40704_, _40273_);
  and (_40706_, _40705_, _40399_);
  and (_40707_, _40706_, _40693_);
  or (_40708_, _40707_, _40681_);
  or (_40709_, _40708_, _40597_);
  not (_40710_, _40597_);
  or (_40711_, _40710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_40712_, _40711_, _41654_);
  and (_42707_, _40712_, _40709_);
  nor (_40713_, _40356_, _40584_);
  nor (_40714_, _40584_, _40561_);
  and (_40715_, _40714_, _40713_);
  and (_40716_, _40402_, _40583_);
  nor (_40717_, _40584_, _40277_);
  and (_40718_, _40717_, _40716_);
  and (_40719_, _40718_, _40715_);
  and (_40720_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_40721_, _40720_, _26533_);
  nor (_40722_, _40721_, _29090_);
  nand (_40723_, _26533_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40724_, _17934_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40725_, _40724_, _40723_);
  nor (_40726_, _38307_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_40727_, _40726_, _40725_);
  or (_40728_, _40727_, _40722_);
  and (_40729_, _40728_, _40583_);
  and (_40730_, _40729_, _40719_);
  not (_40731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_40732_, _40719_, _40731_);
  or (_42719_, _40732_, _40730_);
  nor (_40733_, _40717_, _40716_);
  nor (_40734_, _40714_, _40713_);
  and (_40735_, _40734_, _40583_);
  and (_40736_, _40735_, _40733_);
  and (_40737_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _26512_);
  and (_40738_, _40737_, _26556_);
  nand (_40739_, _40738_, _29090_);
  not (_40740_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40741_, _38285_, _40740_);
  or (_40742_, _16778_, _40740_);
  and (_40743_, _40742_, _40741_);
  or (_40744_, _40743_, _40738_);
  and (_40745_, _40744_, _40739_);
  and (_40746_, _40745_, _40736_);
  not (_40747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_40748_, _40736_, _40747_);
  or (_42974_, _40748_, _40746_);
  nand (_40749_, _40737_, _26633_);
  nor (_40750_, _40749_, _29090_);
  nor (_40751_, _38276_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40752_, _40737_, _26589_);
  and (_40753_, _40737_, _26533_);
  or (_40754_, _40753_, _40720_);
  or (_40755_, _40754_, _40752_);
  and (_40756_, _40755_, _17760_);
  or (_40757_, _40756_, _40751_);
  or (_40758_, _40757_, _40750_);
  and (_40759_, _40758_, _40736_);
  not (_40760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_40761_, _40736_, _40760_);
  or (_42980_, _40761_, _40759_);
  not (_40762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_40763_, _40736_, _40762_);
  nand (_40764_, _40737_, _26600_);
  nor (_40765_, _40764_, _29090_);
  nor (_40766_, _38269_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40767_, _40737_, _26622_);
  or (_40768_, _40767_, _40754_);
  and (_40769_, _40768_, _16415_);
  or (_40770_, _40769_, _40766_);
  or (_40771_, _40770_, _40765_);
  and (_40772_, _40771_, _40736_);
  or (_42986_, _40772_, _40763_);
  not (_40773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_40774_, _40736_, _40773_);
  and (_40775_, _40753_, _29703_);
  nor (_40776_, _38261_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_40777_, _40752_, _40720_);
  or (_40778_, _40777_, _40767_);
  and (_40779_, _40778_, _17444_);
  or (_40780_, _40779_, _40776_);
  or (_40781_, _40780_, _40775_);
  and (_40782_, _40781_, _40736_);
  or (_42992_, _40782_, _40774_);
  not (_40783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_40784_, _40736_, _40783_);
  nand (_40785_, _40720_, _26556_);
  nor (_40786_, _40785_, _29090_);
  nor (_40787_, _38253_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40788_, _26556_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40789_, _16614_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40790_, _40789_, _40788_);
  or (_40791_, _40790_, _40787_);
  or (_40792_, _40791_, _40786_);
  and (_40793_, _40792_, _40736_);
  or (_42998_, _40793_, _40784_);
  nand (_40794_, _40720_, _26633_);
  nor (_40795_, _40794_, _29090_);
  nor (_40796_, _38246_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40797_, _26633_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40798_, _17596_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40799_, _40798_, _40797_);
  or (_40800_, _40799_, _40796_);
  or (_40801_, _40800_, _40795_);
  and (_40802_, _40801_, _40736_);
  not (_40803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_40804_, _40736_, _40803_);
  or (_43004_, _40804_, _40802_);
  not (_40805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_40806_, _40736_, _40805_);
  nand (_40807_, _40720_, _26600_);
  nor (_40808_, _40807_, _29090_);
  nor (_40809_, _38239_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40810_, _26600_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40811_, _16954_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40812_, _40811_, _40810_);
  or (_40813_, _40812_, _40809_);
  or (_40814_, _40813_, _40808_);
  and (_40815_, _40814_, _40736_);
  or (_43010_, _40815_, _40806_);
  not (_40816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_40817_, _40736_, _40816_);
  and (_40818_, _40736_, _40728_);
  or (_43013_, _40818_, _40817_);
  and (_40819_, _40745_, _40583_);
  and (_40820_, _40713_, _40561_);
  and (_40821_, _40820_, _40733_);
  and (_40822_, _40821_, _40819_);
  not (_40823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_40824_, _40821_, _40823_);
  or (_43021_, _40824_, _40822_);
  and (_40825_, _40758_, _40583_);
  and (_40826_, _40821_, _40825_);
  not (_40827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_40828_, _40821_, _40827_);
  or (_43025_, _40828_, _40826_);
  and (_40829_, _40771_, _40583_);
  and (_40830_, _40821_, _40829_);
  not (_40831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_40832_, _40821_, _40831_);
  or (_43029_, _40832_, _40830_);
  and (_40833_, _40781_, _40583_);
  and (_40834_, _40821_, _40833_);
  not (_40835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_40836_, _40821_, _40835_);
  or (_43033_, _40836_, _40834_);
  and (_40837_, _40792_, _40583_);
  and (_40838_, _40821_, _40837_);
  not (_40839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_40840_, _40821_, _40839_);
  or (_43034_, _40840_, _40838_);
  and (_40841_, _40801_, _40583_);
  and (_40842_, _40821_, _40841_);
  not (_40843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_40844_, _40821_, _40843_);
  or (_43038_, _40844_, _40842_);
  and (_40845_, _40814_, _40583_);
  and (_40846_, _40821_, _40845_);
  not (_40847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_40848_, _40821_, _40847_);
  or (_43042_, _40848_, _40846_);
  and (_40849_, _40821_, _40729_);
  nor (_40850_, _40821_, _40608_);
  or (_43045_, _40850_, _40849_);
  and (_40851_, _40714_, _40356_);
  and (_40852_, _40851_, _40733_);
  and (_40853_, _40852_, _40819_);
  not (_40854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_40855_, _40852_, _40854_);
  or (_43053_, _40855_, _40853_);
  and (_40856_, _40852_, _40825_);
  not (_40857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_40858_, _40852_, _40857_);
  or (_43057_, _40858_, _40856_);
  and (_40859_, _40852_, _40829_);
  not (_40860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_40861_, _40852_, _40860_);
  or (_43061_, _40861_, _40859_);
  and (_40862_, _40852_, _40833_);
  not (_40863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_40864_, _40852_, _40863_);
  or (_43065_, _40864_, _40862_);
  and (_40865_, _40852_, _40837_);
  not (_40866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_40867_, _40852_, _40866_);
  or (_43069_, _40867_, _40865_);
  and (_40868_, _40852_, _40841_);
  not (_40869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_40870_, _40852_, _40869_);
  or (_43073_, _40870_, _40868_);
  and (_40871_, _40852_, _40845_);
  not (_40872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_40873_, _40852_, _40872_);
  or (_43077_, _40873_, _40871_);
  and (_40874_, _40852_, _40729_);
  not (_40875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_40876_, _40852_, _40875_);
  or (_43080_, _40876_, _40874_);
  and (_40877_, _40733_, _40715_);
  and (_40878_, _40877_, _40819_);
  not (_40879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_40880_, _40877_, _40879_);
  or (_43086_, _40880_, _40878_);
  and (_40881_, _40877_, _40825_);
  not (_40882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_40883_, _40877_, _40882_);
  or (_43090_, _40883_, _40881_);
  and (_40884_, _40877_, _40829_);
  not (_40885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_40886_, _40877_, _40885_);
  or (_43094_, _40886_, _40884_);
  and (_40887_, _40877_, _40833_);
  not (_40888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_40889_, _40877_, _40888_);
  or (_43098_, _40889_, _40887_);
  and (_40890_, _40877_, _40837_);
  not (_40891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_40892_, _40877_, _40891_);
  or (_43102_, _40892_, _40890_);
  and (_40893_, _40877_, _40841_);
  not (_40894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_40895_, _40877_, _40894_);
  or (_43106_, _40895_, _40893_);
  and (_40896_, _40877_, _40845_);
  not (_40897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_40898_, _40877_, _40897_);
  or (_43110_, _40898_, _40896_);
  and (_40899_, _40877_, _40729_);
  nor (_40900_, _40877_, _40621_);
  or (_43113_, _40900_, _40899_);
  and (_40901_, _40717_, _40403_);
  and (_40902_, _40901_, _40734_);
  and (_40903_, _40902_, _40819_);
  not (_40904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_40905_, _40902_, _40904_);
  or (_43121_, _40905_, _40903_);
  and (_40906_, _40902_, _40825_);
  not (_40907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_40908_, _40902_, _40907_);
  or (_43125_, _40908_, _40906_);
  and (_40909_, _40902_, _40829_);
  not (_40910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_40911_, _40902_, _40910_);
  or (_43129_, _40911_, _40909_);
  and (_40912_, _40902_, _40833_);
  not (_40913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_40914_, _40902_, _40913_);
  or (_43133_, _40914_, _40912_);
  and (_40915_, _40902_, _40837_);
  not (_40916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_40917_, _40902_, _40916_);
  or (_43149_, _40917_, _40915_);
  and (_40918_, _40902_, _40841_);
  not (_40919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_40920_, _40902_, _40919_);
  or (_43169_, _40920_, _40918_);
  and (_40921_, _40902_, _40845_);
  not (_40922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_40923_, _40902_, _40922_);
  or (_43187_, _40923_, _40921_);
  and (_40924_, _40902_, _40729_);
  not (_40925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_40926_, _40902_, _40925_);
  or (_43198_, _40926_, _40924_);
  and (_40927_, _40901_, _40820_);
  and (_40928_, _40927_, _40819_);
  not (_40929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_40930_, _40927_, _40929_);
  or (_43223_, _40930_, _40928_);
  and (_40931_, _40927_, _40825_);
  not (_40932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_40933_, _40927_, _40932_);
  or (_43242_, _40933_, _40931_);
  and (_40934_, _40927_, _40829_);
  not (_40935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_40936_, _40927_, _40935_);
  or (_43262_, _40936_, _40934_);
  and (_40937_, _40927_, _40833_);
  not (_40938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_40939_, _40927_, _40938_);
  or (_43281_, _40939_, _40937_);
  and (_40940_, _40927_, _40837_);
  not (_40941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_40942_, _40927_, _40941_);
  or (_43301_, _40942_, _40940_);
  and (_40943_, _40927_, _40841_);
  not (_40944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_40945_, _40927_, _40944_);
  or (_43321_, _40945_, _40943_);
  and (_40946_, _40927_, _40845_);
  not (_40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_40948_, _40927_, _40947_);
  or (_43339_, _40948_, _40946_);
  and (_40949_, _40927_, _40729_);
  nor (_40950_, _40927_, _40646_);
  or (_43350_, _40950_, _40949_);
  and (_40951_, _40901_, _40851_);
  and (_40952_, _40951_, _40819_);
  not (_40953_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_40954_, _40951_, _40953_);
  or (_43375_, _40954_, _40952_);
  and (_40955_, _40951_, _40825_);
  not (_40956_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_40957_, _40951_, _40956_);
  or (_43379_, _40957_, _40955_);
  and (_40958_, _40951_, _40829_);
  not (_40959_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_40960_, _40951_, _40959_);
  or (_43383_, _40960_, _40958_);
  and (_40961_, _40951_, _40833_);
  not (_40962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_40963_, _40951_, _40962_);
  or (_43387_, _40963_, _40961_);
  and (_40964_, _40951_, _40837_);
  not (_40965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_40966_, _40951_, _40965_);
  or (_43391_, _40966_, _40964_);
  and (_40967_, _40951_, _40841_);
  not (_40968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_40969_, _40951_, _40968_);
  or (_43395_, _40969_, _40967_);
  and (_40970_, _40951_, _40845_);
  not (_40971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_40972_, _40951_, _40971_);
  or (_43399_, _40972_, _40970_);
  and (_40973_, _40951_, _40729_);
  not (_40974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_40975_, _40951_, _40974_);
  or (_43402_, _40975_, _40973_);
  and (_40976_, _40901_, _40715_);
  and (_40977_, _40976_, _40819_);
  not (_40978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_40979_, _40976_, _40978_);
  or (_43407_, _40979_, _40977_);
  and (_40980_, _40976_, _40825_);
  not (_40981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_40982_, _40976_, _40981_);
  or (_43411_, _40982_, _40980_);
  and (_40983_, _40976_, _40829_);
  not (_40984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_40985_, _40976_, _40984_);
  or (_43415_, _40985_, _40983_);
  and (_40986_, _40976_, _40833_);
  not (_40987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_40988_, _40976_, _40987_);
  or (_43419_, _40988_, _40986_);
  and (_40989_, _40976_, _40837_);
  not (_40990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_40991_, _40976_, _40990_);
  or (_43423_, _40991_, _40989_);
  and (_40992_, _40976_, _40841_);
  not (_40993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_40994_, _40976_, _40993_);
  or (_43427_, _40994_, _40992_);
  and (_40995_, _40976_, _40845_);
  not (_40996_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_40997_, _40976_, _40996_);
  or (_43431_, _40997_, _40995_);
  and (_40998_, _40976_, _40729_);
  nor (_40999_, _40976_, _40658_);
  or (_43434_, _40999_, _40998_);
  and (_41000_, _40716_, _40277_);
  and (_41001_, _41000_, _40734_);
  and (_41002_, _41001_, _40819_);
  not (_41003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_41004_, _41001_, _41003_);
  or (_43441_, _41004_, _41002_);
  and (_41005_, _41001_, _40825_);
  not (_41006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_41007_, _41001_, _41006_);
  or (_43445_, _41007_, _41005_);
  and (_41008_, _41001_, _40829_);
  not (_41009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_41010_, _41001_, _41009_);
  or (_43449_, _41010_, _41008_);
  and (_41011_, _41001_, _40833_);
  not (_41012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_41013_, _41001_, _41012_);
  or (_43453_, _41013_, _41011_);
  and (_41014_, _41001_, _40837_);
  not (_41015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_41016_, _41001_, _41015_);
  or (_43457_, _41016_, _41014_);
  and (_41017_, _41001_, _40841_);
  not (_41018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_41019_, _41001_, _41018_);
  or (_43461_, _41019_, _41017_);
  and (_41020_, _41001_, _40845_);
  not (_41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_41022_, _41001_, _41021_);
  or (_43465_, _41022_, _41020_);
  and (_41023_, _41001_, _40729_);
  nor (_41024_, _41001_, _40682_);
  or (_43468_, _41024_, _41023_);
  and (_41025_, _41000_, _40820_);
  and (_41026_, _41025_, _40819_);
  not (_41027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_41028_, _41025_, _41027_);
  or (_43473_, _41028_, _41026_);
  and (_41029_, _41025_, _40825_);
  not (_41030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_41031_, _41025_, _41030_);
  or (_43477_, _41031_, _41029_);
  and (_41032_, _41025_, _40829_);
  not (_41033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_41034_, _41025_, _41033_);
  or (_43481_, _41034_, _41032_);
  and (_41035_, _41025_, _40833_);
  not (_41036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_41037_, _41025_, _41036_);
  or (_43485_, _41037_, _41035_);
  and (_41038_, _41025_, _40837_);
  not (_41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_41040_, _41025_, _41039_);
  or (_43489_, _41040_, _41038_);
  and (_41041_, _41025_, _40841_);
  not (_41042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_41043_, _41025_, _41042_);
  or (_43493_, _41043_, _41041_);
  and (_41044_, _41025_, _40845_);
  not (_41045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_41046_, _41025_, _41045_);
  or (_43497_, _41046_, _41044_);
  and (_41047_, _41025_, _40729_);
  not (_41048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_41049_, _41025_, _41048_);
  or (_43500_, _41049_, _41047_);
  and (_41050_, _41000_, _40851_);
  and (_41051_, _41050_, _40819_);
  not (_41052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_41053_, _41050_, _41052_);
  or (_43505_, _41053_, _41051_);
  and (_41054_, _41050_, _40825_);
  not (_41055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_41056_, _41050_, _41055_);
  or (_43509_, _41056_, _41054_);
  and (_41057_, _41050_, _40829_);
  not (_41058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_41060_, _41050_, _41058_);
  or (_43513_, _41060_, _41057_);
  and (_41063_, _41050_, _40833_);
  not (_41065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_41067_, _41050_, _41065_);
  or (_43517_, _41067_, _41063_);
  and (_41070_, _41050_, _40837_);
  not (_41072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_41074_, _41050_, _41072_);
  or (_43521_, _41074_, _41070_);
  and (_41077_, _41050_, _40841_);
  not (_41079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_41081_, _41050_, _41079_);
  or (_43525_, _41081_, _41077_);
  and (_41084_, _41050_, _40845_);
  not (_41086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_41088_, _41050_, _41086_);
  or (_43529_, _41088_, _41084_);
  and (_41091_, _41050_, _40729_);
  nor (_41093_, _41050_, _40688_);
  or (_43532_, _41093_, _41091_);
  and (_41096_, _41000_, _40715_);
  and (_41098_, _41096_, _40819_);
  not (_41100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_41102_, _41096_, _41100_);
  or (_43537_, _41102_, _41098_);
  and (_41105_, _41096_, _40825_);
  not (_41107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_41108_, _41096_, _41107_);
  or (_43541_, _41108_, _41105_);
  and (_41109_, _41096_, _40829_);
  not (_41110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_41111_, _41096_, _41110_);
  or (_43545_, _41111_, _41109_);
  and (_41112_, _41096_, _40833_);
  not (_41113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_41114_, _41096_, _41113_);
  or (_43549_, _41114_, _41112_);
  and (_41115_, _41096_, _40837_);
  not (_41116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_41117_, _41096_, _41116_);
  or (_43553_, _41117_, _41115_);
  and (_41118_, _41096_, _40841_);
  not (_41119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_41120_, _41096_, _41119_);
  or (_43557_, _41120_, _41118_);
  and (_41121_, _41096_, _40845_);
  not (_41122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_41123_, _41096_, _41122_);
  or (_43561_, _41123_, _41121_);
  and (_41124_, _41096_, _40729_);
  not (_41125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_41126_, _41096_, _41125_);
  or (_43564_, _41126_, _41124_);
  and (_41127_, _40734_, _40718_);
  and (_41128_, _41127_, _40819_);
  not (_41129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_41130_, _41127_, _41129_);
  or (_43570_, _41130_, _41128_);
  and (_41131_, _41127_, _40825_);
  not (_41132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_41133_, _41127_, _41132_);
  or (_43574_, _41133_, _41131_);
  and (_41134_, _41127_, _40829_);
  not (_41135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_41136_, _41127_, _41135_);
  or (_43578_, _41136_, _41134_);
  and (_41137_, _41127_, _40833_);
  not (_41138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_41139_, _41127_, _41138_);
  or (_43582_, _41139_, _41137_);
  and (_41140_, _41127_, _40837_);
  not (_41141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_41142_, _41127_, _41141_);
  or (_43586_, _41142_, _41140_);
  and (_41143_, _41127_, _40841_);
  not (_41144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_41145_, _41127_, _41144_);
  or (_43590_, _41145_, _41143_);
  and (_41146_, _41127_, _40845_);
  not (_41147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_41148_, _41127_, _41147_);
  or (_43594_, _41148_, _41146_);
  and (_41149_, _41127_, _40729_);
  nor (_41150_, _41127_, _40694_);
  or (_43597_, _41150_, _41149_);
  and (_41151_, _40820_, _40718_);
  and (_41152_, _41151_, _40819_);
  not (_41153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_41154_, _41151_, _41153_);
  or (_43602_, _41154_, _41152_);
  and (_41155_, _41151_, _40825_);
  not (_41156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_41157_, _41151_, _41156_);
  or (_43606_, _41157_, _41155_);
  and (_41158_, _41151_, _40829_);
  not (_41159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_41160_, _41151_, _41159_);
  or (_43610_, _41160_, _41158_);
  and (_41161_, _41151_, _40833_);
  not (_41162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_41163_, _41151_, _41162_);
  or (_43614_, _41163_, _41161_);
  and (_41164_, _41151_, _40837_);
  not (_41165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_41166_, _41151_, _41165_);
  or (_43618_, _41166_, _41164_);
  and (_41167_, _41151_, _40841_);
  not (_41168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_41169_, _41151_, _41168_);
  or (_43622_, _41169_, _41167_);
  and (_41170_, _41151_, _40845_);
  not (_41171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_41172_, _41151_, _41171_);
  or (_43626_, _41172_, _41170_);
  and (_41173_, _41151_, _40729_);
  not (_41174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_41175_, _41151_, _41174_);
  or (_43629_, _41175_, _41173_);
  and (_41176_, _40851_, _40718_);
  and (_41177_, _41176_, _40819_);
  not (_41178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_41179_, _41176_, _41178_);
  or (_43634_, _41179_, _41177_);
  and (_41180_, _41176_, _40825_);
  not (_41181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_41182_, _41176_, _41181_);
  or (_43638_, _41182_, _41180_);
  and (_41183_, _41176_, _40829_);
  not (_41184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_41185_, _41176_, _41184_);
  or (_43642_, _41185_, _41183_);
  and (_41186_, _41176_, _40833_);
  not (_41187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_41188_, _41176_, _41187_);
  or (_43646_, _41188_, _41186_);
  and (_41189_, _41176_, _40837_);
  not (_41190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_41191_, _41176_, _41190_);
  or (_43650_, _41191_, _41189_);
  and (_41192_, _41176_, _40841_);
  not (_41193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_41194_, _41176_, _41193_);
  or (_43654_, _41194_, _41192_);
  and (_41195_, _41176_, _40845_);
  not (_41196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_41197_, _41176_, _41196_);
  or (_43658_, _41197_, _41195_);
  and (_41198_, _41176_, _40729_);
  nor (_41199_, _41176_, _40700_);
  or (_43661_, _41199_, _41198_);
  and (_41200_, _40819_, _40719_);
  not (_41201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_41202_, _40719_, _41201_);
  or (_43666_, _41202_, _41200_);
  and (_41203_, _40825_, _40719_);
  not (_41204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_41205_, _40719_, _41204_);
  or (_43670_, _41205_, _41203_);
  and (_41206_, _40829_, _40719_);
  not (_41207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_41208_, _40719_, _41207_);
  or (_43674_, _41208_, _41206_);
  and (_41209_, _40833_, _40719_);
  not (_41210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_41211_, _40719_, _41210_);
  or (_43678_, _41211_, _41209_);
  and (_41212_, _40837_, _40719_);
  not (_41213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_41214_, _40719_, _41213_);
  or (_43682_, _41214_, _41212_);
  and (_41215_, _40841_, _40719_);
  not (_41216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_41217_, _40719_, _41216_);
  or (_43686_, _41217_, _41215_);
  and (_41218_, _40845_, _40719_);
  not (_41219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_41220_, _40719_, _41219_);
  or (_43690_, _41220_, _41218_);
  and (_41221_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_41222_, _40353_, _40823_);
  or (_41223_, _41222_, _41221_);
  and (_41224_, _41223_, _40555_);
  nor (_41225_, _40353_, _40879_);
  and (_41226_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_41227_, _41226_, _41225_);
  and (_41228_, _41227_, _40620_);
  or (_41229_, _41228_, _41224_);
  or (_41230_, _41229_, _40598_);
  and (_41231_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_41232_, _40353_, _40929_);
  or (_41233_, _41232_, _41231_);
  and (_41234_, _41233_, _40555_);
  nor (_41235_, _40353_, _40978_);
  and (_41236_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_41237_, _41236_, _41235_);
  and (_41238_, _41237_, _40620_);
  or (_41239_, _41238_, _41234_);
  or (_41240_, _41239_, _40273_);
  and (_41241_, _41240_, _40644_);
  and (_41242_, _41241_, _41230_);
  nand (_41243_, _40353_, _41003_);
  or (_41244_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_41245_, _41244_, _41243_);
  and (_41246_, _41245_, _40555_);
  or (_41247_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand (_41248_, _40353_, _41052_);
  and (_41249_, _41248_, _41247_);
  and (_41250_, _41249_, _40620_);
  or (_41251_, _41250_, _41246_);
  or (_41252_, _41251_, _40598_);
  nand (_41253_, _40353_, _41129_);
  or (_41254_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_41255_, _41254_, _41253_);
  and (_41256_, _41255_, _40555_);
  or (_41257_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand (_41258_, _40353_, _41178_);
  and (_41259_, _41258_, _41257_);
  and (_41260_, _41259_, _40620_);
  or (_41261_, _41260_, _41256_);
  or (_41262_, _41261_, _40273_);
  and (_41263_, _41262_, _40399_);
  and (_41264_, _41263_, _41252_);
  or (_41265_, _41264_, _41242_);
  or (_41266_, _41265_, _40597_);
  or (_41267_, _40710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_41268_, _41267_, _41654_);
  and (_01364_, _41268_, _41266_);
  and (_41269_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_41270_, _40353_, _40827_);
  or (_41271_, _41270_, _41269_);
  and (_41272_, _41271_, _40555_);
  nor (_41273_, _40353_, _40882_);
  and (_41274_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_41275_, _41274_, _41273_);
  and (_41276_, _41275_, _40620_);
  or (_41277_, _41276_, _41272_);
  or (_41278_, _41277_, _40598_);
  and (_41279_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_41280_, _40353_, _40932_);
  or (_41281_, _41280_, _41279_);
  and (_41282_, _41281_, _40555_);
  nor (_41283_, _40353_, _40981_);
  and (_41284_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_41285_, _41284_, _41283_);
  and (_41286_, _41285_, _40620_);
  or (_41287_, _41286_, _41282_);
  or (_41288_, _41287_, _40273_);
  and (_41289_, _41288_, _40644_);
  and (_41290_, _41289_, _41278_);
  nand (_41291_, _40353_, _41006_);
  or (_41292_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_41293_, _41292_, _41291_);
  and (_41294_, _41293_, _40555_);
  or (_41295_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand (_41296_, _40353_, _41055_);
  and (_41297_, _41296_, _41295_);
  and (_41298_, _41297_, _40620_);
  or (_41299_, _41298_, _41294_);
  or (_41300_, _41299_, _40598_);
  nand (_41301_, _40353_, _41132_);
  or (_41302_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_41303_, _41302_, _41301_);
  and (_41304_, _41303_, _40555_);
  or (_41305_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand (_41306_, _40353_, _41181_);
  and (_41307_, _41306_, _41305_);
  and (_41308_, _41307_, _40620_);
  or (_41309_, _41308_, _41304_);
  or (_41310_, _41309_, _40273_);
  and (_41311_, _41310_, _40399_);
  and (_41312_, _41311_, _41300_);
  or (_41313_, _41312_, _41290_);
  or (_41314_, _41313_, _40597_);
  or (_41315_, _40710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_41316_, _41315_, _41654_);
  and (_01366_, _41316_, _41314_);
  and (_41317_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_41318_, _40353_, _40831_);
  or (_41319_, _41318_, _41317_);
  and (_41320_, _41319_, _40555_);
  nor (_41321_, _40353_, _40885_);
  and (_41322_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_41323_, _41322_, _41321_);
  and (_41324_, _41323_, _40620_);
  or (_41325_, _41324_, _41320_);
  or (_41326_, _41325_, _40598_);
  and (_41327_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_41328_, _40353_, _40935_);
  or (_41329_, _41328_, _41327_);
  and (_41330_, _41329_, _40555_);
  nor (_41331_, _40353_, _40984_);
  and (_41332_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_41333_, _41332_, _41331_);
  and (_41334_, _41333_, _40620_);
  or (_41335_, _41334_, _41330_);
  or (_41336_, _41335_, _40273_);
  and (_41337_, _41336_, _40644_);
  and (_41338_, _41337_, _41326_);
  nand (_41339_, _40353_, _41009_);
  or (_41340_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_41341_, _41340_, _41339_);
  and (_41342_, _41341_, _40555_);
  or (_41343_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_41344_, _40353_, _41058_);
  and (_41345_, _41344_, _41343_);
  and (_41346_, _41345_, _40620_);
  or (_41347_, _41346_, _41342_);
  or (_41348_, _41347_, _40598_);
  nand (_41349_, _40353_, _41135_);
  or (_41350_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_41351_, _41350_, _41349_);
  and (_41352_, _41351_, _40555_);
  or (_41353_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_41354_, _40353_, _41184_);
  and (_41355_, _41354_, _41353_);
  and (_41356_, _41355_, _40620_);
  or (_41357_, _41356_, _41352_);
  or (_41358_, _41357_, _40273_);
  and (_41359_, _41358_, _40399_);
  and (_41360_, _41359_, _41348_);
  or (_41361_, _41360_, _41338_);
  or (_41362_, _41361_, _40597_);
  or (_41363_, _40710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_41364_, _41363_, _41654_);
  and (_01368_, _41364_, _41362_);
  and (_41365_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_41366_, _40353_, _40835_);
  or (_41367_, _41366_, _41365_);
  and (_41368_, _41367_, _40555_);
  nor (_41369_, _40353_, _40888_);
  and (_41370_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_41371_, _41370_, _41369_);
  and (_41372_, _41371_, _40620_);
  or (_41373_, _41372_, _41368_);
  or (_41374_, _41373_, _40598_);
  and (_41375_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_41376_, _40353_, _40938_);
  or (_41377_, _41376_, _41375_);
  and (_41378_, _41377_, _40555_);
  nor (_41379_, _40353_, _40987_);
  and (_41380_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_41381_, _41380_, _41379_);
  and (_41382_, _41381_, _40620_);
  or (_41383_, _41382_, _41378_);
  or (_41384_, _41383_, _40273_);
  and (_41385_, _41384_, _40644_);
  and (_41386_, _41385_, _41374_);
  nand (_41387_, _40353_, _41012_);
  or (_41388_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_41389_, _41388_, _41387_);
  and (_41390_, _41389_, _40555_);
  or (_41391_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_41392_, _40353_, _41065_);
  and (_41393_, _41392_, _41391_);
  and (_41394_, _41393_, _40620_);
  or (_41395_, _41394_, _41390_);
  or (_41396_, _41395_, _40598_);
  nand (_41397_, _40353_, _41138_);
  or (_41398_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_41399_, _41398_, _41397_);
  and (_41400_, _41399_, _40555_);
  or (_41401_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_41402_, _40353_, _41187_);
  and (_41403_, _41402_, _41401_);
  and (_41404_, _41403_, _40620_);
  or (_41405_, _41404_, _41400_);
  or (_41406_, _41405_, _40273_);
  and (_41407_, _41406_, _40399_);
  and (_41408_, _41407_, _41396_);
  or (_41409_, _41408_, _41386_);
  or (_41410_, _41409_, _40597_);
  or (_41411_, _40710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_41412_, _41411_, _41654_);
  and (_01370_, _41412_, _41410_);
  and (_41413_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_41414_, _40353_, _40839_);
  or (_41415_, _41414_, _41413_);
  and (_41416_, _41415_, _40555_);
  nor (_41417_, _40353_, _40891_);
  and (_41418_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_41419_, _41418_, _41417_);
  and (_41420_, _41419_, _40620_);
  or (_41421_, _41420_, _41416_);
  or (_41422_, _41421_, _40598_);
  and (_41423_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_41424_, _40353_, _40941_);
  or (_41425_, _41424_, _41423_);
  and (_41426_, _41425_, _40555_);
  nor (_41427_, _40353_, _40990_);
  and (_41428_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_41429_, _41428_, _41427_);
  and (_41430_, _41429_, _40620_);
  or (_41431_, _41430_, _41426_);
  or (_41432_, _41431_, _40273_);
  and (_41433_, _41432_, _40644_);
  and (_41434_, _41433_, _41422_);
  nand (_41435_, _40353_, _41015_);
  or (_41436_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_41437_, _41436_, _41435_);
  and (_41438_, _41437_, _40555_);
  or (_41439_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_41440_, _40353_, _41072_);
  and (_41441_, _41440_, _41439_);
  and (_41442_, _41441_, _40620_);
  or (_41443_, _41442_, _41438_);
  or (_41444_, _41443_, _40598_);
  nand (_41445_, _40353_, _41141_);
  or (_41446_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_41447_, _41446_, _41445_);
  and (_41448_, _41447_, _40555_);
  or (_41449_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_41450_, _40353_, _41190_);
  and (_41451_, _41450_, _41449_);
  and (_41452_, _41451_, _40620_);
  or (_41453_, _41452_, _41448_);
  or (_41454_, _41453_, _40273_);
  and (_41455_, _41454_, _40399_);
  and (_41456_, _41455_, _41444_);
  or (_41457_, _41456_, _41434_);
  or (_41458_, _41457_, _40597_);
  or (_41459_, _40710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_41460_, _41459_, _41654_);
  and (_01372_, _41460_, _41458_);
  and (_41461_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_41462_, _40353_, _40843_);
  or (_41463_, _41462_, _41461_);
  and (_41464_, _41463_, _40555_);
  nor (_41465_, _40353_, _40894_);
  and (_41466_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_41467_, _41466_, _41465_);
  and (_41468_, _41467_, _40620_);
  or (_41469_, _41468_, _41464_);
  or (_41470_, _41469_, _40598_);
  and (_41471_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_41472_, _40353_, _40944_);
  or (_41473_, _41472_, _41471_);
  and (_41474_, _41473_, _40555_);
  nor (_41475_, _40353_, _40993_);
  and (_41476_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_41477_, _41476_, _41475_);
  and (_41478_, _41477_, _40620_);
  or (_41479_, _41478_, _41474_);
  or (_41480_, _41479_, _40273_);
  and (_41481_, _41480_, _40644_);
  and (_41482_, _41481_, _41470_);
  nand (_41483_, _40353_, _41018_);
  or (_41484_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_41485_, _41484_, _41483_);
  and (_41486_, _41485_, _40555_);
  or (_41487_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_41488_, _40353_, _41079_);
  and (_41489_, _41488_, _41487_);
  and (_41490_, _41489_, _40620_);
  or (_41491_, _41490_, _41486_);
  or (_41492_, _41491_, _40598_);
  nand (_41493_, _40353_, _41144_);
  or (_41494_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_41495_, _41494_, _41493_);
  and (_41496_, _41495_, _40555_);
  or (_41497_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_41498_, _40353_, _41193_);
  and (_41499_, _41498_, _41497_);
  and (_41500_, _41499_, _40620_);
  or (_41501_, _41500_, _41496_);
  or (_41502_, _41501_, _40273_);
  and (_41503_, _41502_, _40399_);
  and (_41504_, _41503_, _41492_);
  or (_41505_, _41504_, _41482_);
  or (_41506_, _41505_, _40597_);
  or (_41507_, _40710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_41508_, _41507_, _41654_);
  and (_01374_, _41508_, _41506_);
  and (_41509_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_41510_, _40353_, _40847_);
  or (_41511_, _41510_, _41509_);
  and (_41512_, _41511_, _40555_);
  nor (_41513_, _40353_, _40897_);
  and (_41514_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_41515_, _41514_, _41513_);
  and (_41516_, _41515_, _40620_);
  or (_41517_, _41516_, _41512_);
  or (_41518_, _41517_, _40598_);
  and (_41519_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_41520_, _40353_, _40947_);
  or (_41521_, _41520_, _41519_);
  and (_41522_, _41521_, _40555_);
  nor (_41523_, _40353_, _40996_);
  and (_41524_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_41525_, _41524_, _41523_);
  and (_41526_, _41525_, _40620_);
  or (_41527_, _41526_, _41522_);
  or (_41528_, _41527_, _40273_);
  and (_41529_, _41528_, _40644_);
  and (_41530_, _41529_, _41518_);
  nand (_41531_, _40353_, _41021_);
  or (_41532_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_41533_, _41532_, _41531_);
  and (_41534_, _41533_, _40555_);
  or (_41535_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_41536_, _40353_, _41086_);
  and (_41537_, _41536_, _41535_);
  and (_41538_, _41537_, _40620_);
  or (_41539_, _41538_, _41534_);
  or (_41540_, _41539_, _40598_);
  nand (_41541_, _40353_, _41147_);
  or (_41542_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_41543_, _41542_, _41541_);
  and (_41544_, _41543_, _40555_);
  or (_41545_, _40353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_41546_, _40353_, _41196_);
  and (_41547_, _41546_, _41545_);
  and (_41548_, _41547_, _40620_);
  or (_41549_, _41548_, _41544_);
  or (_41550_, _41549_, _40273_);
  and (_41551_, _41550_, _40399_);
  and (_41552_, _41551_, _41540_);
  or (_41553_, _41552_, _41530_);
  or (_41554_, _41553_, _40597_);
  or (_41555_, _40710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_41556_, _41555_, _41654_);
  and (_01376_, _41556_, _41554_);
  or (_41557_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_41558_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_41559_, _41558_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_41560_, _41559_, _41557_);
  nand (_41561_, _41560_, _41654_);
  or (_41562_, \oc8051_gm_cxrom_1.cell0.data [7], _41654_);
  and (_01384_, _41562_, _41561_);
  or (_41563_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41564_, \oc8051_gm_cxrom_1.cell0.data [0], _41558_);
  nand (_41565_, _41564_, _41563_);
  nand (_41566_, _41565_, _41654_);
  or (_41567_, \oc8051_gm_cxrom_1.cell0.data [0], _41654_);
  and (_01391_, _41567_, _41566_);
  or (_41568_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41569_, \oc8051_gm_cxrom_1.cell0.data [1], _41558_);
  nand (_41570_, _41569_, _41568_);
  nand (_41571_, _41570_, _41654_);
  or (_41572_, \oc8051_gm_cxrom_1.cell0.data [1], _41654_);
  and (_01395_, _41572_, _41571_);
  or (_41573_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41574_, \oc8051_gm_cxrom_1.cell0.data [2], _41558_);
  nand (_41575_, _41574_, _41573_);
  nand (_41576_, _41575_, _41654_);
  or (_41577_, \oc8051_gm_cxrom_1.cell0.data [2], _41654_);
  and (_01399_, _41577_, _41576_);
  or (_41578_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41579_, \oc8051_gm_cxrom_1.cell0.data [3], _41558_);
  nand (_41580_, _41579_, _41578_);
  nand (_41581_, _41580_, _41654_);
  or (_41582_, \oc8051_gm_cxrom_1.cell0.data [3], _41654_);
  and (_01403_, _41582_, _41581_);
  or (_41583_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41584_, \oc8051_gm_cxrom_1.cell0.data [4], _41558_);
  nand (_41585_, _41584_, _41583_);
  nand (_41586_, _41585_, _41654_);
  or (_41587_, \oc8051_gm_cxrom_1.cell0.data [4], _41654_);
  and (_01407_, _41587_, _41586_);
  or (_41588_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41589_, \oc8051_gm_cxrom_1.cell0.data [5], _41558_);
  nand (_41590_, _41589_, _41588_);
  nand (_41591_, _41590_, _41654_);
  or (_41592_, \oc8051_gm_cxrom_1.cell0.data [5], _41654_);
  and (_01411_, _41592_, _41591_);
  or (_41593_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41594_, \oc8051_gm_cxrom_1.cell0.data [6], _41558_);
  nand (_41595_, _41594_, _41593_);
  nand (_41596_, _41595_, _41654_);
  or (_41598_, \oc8051_gm_cxrom_1.cell0.data [6], _41654_);
  and (_01415_, _41598_, _41596_);
  or (_41600_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_41602_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_41603_, _41602_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_41605_, _41603_, _41600_);
  nand (_41607_, _41605_, _41654_);
  or (_41609_, \oc8051_gm_cxrom_1.cell1.data [7], _41654_);
  and (_01437_, _41609_, _41607_);
  or (_41611_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41612_, \oc8051_gm_cxrom_1.cell1.data [0], _41602_);
  nand (_41613_, _41612_, _41611_);
  nand (_41614_, _41613_, _41654_);
  or (_41615_, \oc8051_gm_cxrom_1.cell1.data [0], _41654_);
  and (_01444_, _41615_, _41614_);
  or (_41616_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41617_, \oc8051_gm_cxrom_1.cell1.data [1], _41602_);
  nand (_41618_, _41617_, _41616_);
  nand (_41619_, _41618_, _41654_);
  or (_41620_, \oc8051_gm_cxrom_1.cell1.data [1], _41654_);
  and (_01448_, _41620_, _41619_);
  or (_41621_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41622_, \oc8051_gm_cxrom_1.cell1.data [2], _41602_);
  nand (_41623_, _41622_, _41621_);
  nand (_41624_, _41623_, _41654_);
  or (_41625_, \oc8051_gm_cxrom_1.cell1.data [2], _41654_);
  and (_01452_, _41625_, _41624_);
  or (_41626_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41627_, \oc8051_gm_cxrom_1.cell1.data [3], _41602_);
  nand (_41628_, _41627_, _41626_);
  nand (_41629_, _41628_, _41654_);
  or (_41630_, \oc8051_gm_cxrom_1.cell1.data [3], _41654_);
  and (_01456_, _41630_, _41629_);
  or (_41631_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41632_, \oc8051_gm_cxrom_1.cell1.data [4], _41602_);
  nand (_41633_, _41632_, _41631_);
  nand (_41634_, _41633_, _41654_);
  or (_41635_, \oc8051_gm_cxrom_1.cell1.data [4], _41654_);
  and (_01460_, _41635_, _41634_);
  or (_41636_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41637_, \oc8051_gm_cxrom_1.cell1.data [5], _41602_);
  nand (_41638_, _41637_, _41636_);
  nand (_41639_, _41638_, _41654_);
  or (_41640_, \oc8051_gm_cxrom_1.cell1.data [5], _41654_);
  and (_01464_, _41640_, _41639_);
  or (_41642_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41644_, \oc8051_gm_cxrom_1.cell1.data [6], _41602_);
  nand (_41646_, _41644_, _41642_);
  nand (_41648_, _41646_, _41654_);
  or (_41650_, \oc8051_gm_cxrom_1.cell1.data [6], _41654_);
  and (_01468_, _41650_, _41648_);
  or (_41653_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_41655_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_41656_, _41655_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_41657_, _41656_, _41653_);
  nand (_41658_, _41657_, _41654_);
  or (_41659_, \oc8051_gm_cxrom_1.cell2.data [7], _41654_);
  and (_01490_, _41659_, _41658_);
  or (_41660_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41661_, \oc8051_gm_cxrom_1.cell2.data [0], _41655_);
  nand (_41662_, _41661_, _41660_);
  nand (_41663_, _41662_, _41654_);
  or (_41664_, \oc8051_gm_cxrom_1.cell2.data [0], _41654_);
  and (_01497_, _41664_, _41663_);
  or (_41665_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41666_, \oc8051_gm_cxrom_1.cell2.data [1], _41655_);
  nand (_41667_, _41666_, _41665_);
  nand (_41668_, _41667_, _41654_);
  or (_41669_, \oc8051_gm_cxrom_1.cell2.data [1], _41654_);
  and (_01501_, _41669_, _41668_);
  or (_41670_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41671_, \oc8051_gm_cxrom_1.cell2.data [2], _41655_);
  nand (_41672_, _41671_, _41670_);
  nand (_41673_, _41672_, _41654_);
  or (_41674_, \oc8051_gm_cxrom_1.cell2.data [2], _41654_);
  and (_01505_, _41674_, _41673_);
  or (_41675_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41676_, \oc8051_gm_cxrom_1.cell2.data [3], _41655_);
  nand (_41677_, _41676_, _41675_);
  nand (_41678_, _41677_, _41654_);
  or (_41679_, \oc8051_gm_cxrom_1.cell2.data [3], _41654_);
  and (_01509_, _41679_, _41678_);
  or (_41680_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41681_, \oc8051_gm_cxrom_1.cell2.data [4], _41655_);
  nand (_41682_, _41681_, _41680_);
  nand (_41683_, _41682_, _41654_);
  or (_41684_, \oc8051_gm_cxrom_1.cell2.data [4], _41654_);
  and (_01513_, _41684_, _41683_);
  or (_41685_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41686_, \oc8051_gm_cxrom_1.cell2.data [5], _41655_);
  nand (_41687_, _41686_, _41685_);
  nand (_41688_, _41687_, _41654_);
  or (_41689_, \oc8051_gm_cxrom_1.cell2.data [5], _41654_);
  and (_01517_, _41689_, _41688_);
  or (_41690_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41691_, \oc8051_gm_cxrom_1.cell2.data [6], _41655_);
  nand (_41692_, _41691_, _41690_);
  nand (_41693_, _41692_, _41654_);
  or (_41694_, \oc8051_gm_cxrom_1.cell2.data [6], _41654_);
  and (_01521_, _41694_, _41693_);
  or (_41695_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_41696_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_41697_, _41696_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_41698_, _41697_, _41695_);
  nand (_41699_, _41698_, _41654_);
  or (_41700_, \oc8051_gm_cxrom_1.cell3.data [7], _41654_);
  and (_01542_, _41700_, _41699_);
  or (_41701_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41702_, \oc8051_gm_cxrom_1.cell3.data [0], _41696_);
  nand (_41703_, _41702_, _41701_);
  nand (_41704_, _41703_, _41654_);
  or (_41705_, \oc8051_gm_cxrom_1.cell3.data [0], _41654_);
  and (_01549_, _41705_, _41704_);
  or (_41706_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41707_, \oc8051_gm_cxrom_1.cell3.data [1], _41696_);
  nand (_41708_, _41707_, _41706_);
  nand (_41709_, _41708_, _41654_);
  or (_41710_, \oc8051_gm_cxrom_1.cell3.data [1], _41654_);
  and (_01552_, _41710_, _41709_);
  or (_41711_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41712_, \oc8051_gm_cxrom_1.cell3.data [2], _41696_);
  nand (_41713_, _41712_, _41711_);
  nand (_41714_, _41713_, _41654_);
  or (_41715_, \oc8051_gm_cxrom_1.cell3.data [2], _41654_);
  and (_01556_, _41715_, _41714_);
  or (_41716_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41717_, \oc8051_gm_cxrom_1.cell3.data [3], _41696_);
  nand (_41718_, _41717_, _41716_);
  nand (_41719_, _41718_, _41654_);
  or (_41720_, \oc8051_gm_cxrom_1.cell3.data [3], _41654_);
  and (_01560_, _41720_, _41719_);
  or (_41721_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41722_, \oc8051_gm_cxrom_1.cell3.data [4], _41696_);
  nand (_41723_, _41722_, _41721_);
  nand (_41724_, _41723_, _41654_);
  or (_41725_, \oc8051_gm_cxrom_1.cell3.data [4], _41654_);
  and (_01564_, _41725_, _41724_);
  or (_41726_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41727_, \oc8051_gm_cxrom_1.cell3.data [5], _41696_);
  nand (_41728_, _41727_, _41726_);
  nand (_41729_, _41728_, _41654_);
  or (_41730_, \oc8051_gm_cxrom_1.cell3.data [5], _41654_);
  and (_01568_, _41730_, _41729_);
  or (_41731_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41732_, \oc8051_gm_cxrom_1.cell3.data [6], _41696_);
  nand (_41733_, _41732_, _41731_);
  nand (_41734_, _41733_, _41654_);
  or (_41735_, \oc8051_gm_cxrom_1.cell3.data [6], _41654_);
  and (_01572_, _41735_, _41734_);
  or (_41736_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_41737_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_41738_, _41737_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_41739_, _41738_, _41736_);
  nand (_41740_, _41739_, _41654_);
  or (_41741_, \oc8051_gm_cxrom_1.cell4.data [7], _41654_);
  and (_01594_, _41741_, _41740_);
  or (_41742_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41743_, \oc8051_gm_cxrom_1.cell4.data [0], _41737_);
  nand (_41744_, _41743_, _41742_);
  nand (_41745_, _41744_, _41654_);
  or (_41746_, \oc8051_gm_cxrom_1.cell4.data [0], _41654_);
  and (_01601_, _41746_, _41745_);
  or (_41747_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41748_, \oc8051_gm_cxrom_1.cell4.data [1], _41737_);
  nand (_41749_, _41748_, _41747_);
  nand (_41750_, _41749_, _41654_);
  or (_41751_, \oc8051_gm_cxrom_1.cell4.data [1], _41654_);
  and (_01605_, _41751_, _41750_);
  or (_41752_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41753_, \oc8051_gm_cxrom_1.cell4.data [2], _41737_);
  nand (_41754_, _41753_, _41752_);
  nand (_41755_, _41754_, _41654_);
  or (_41756_, \oc8051_gm_cxrom_1.cell4.data [2], _41654_);
  and (_01609_, _41756_, _41755_);
  or (_41757_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41758_, \oc8051_gm_cxrom_1.cell4.data [3], _41737_);
  nand (_41759_, _41758_, _41757_);
  nand (_41760_, _41759_, _41654_);
  or (_41761_, \oc8051_gm_cxrom_1.cell4.data [3], _41654_);
  and (_01613_, _41761_, _41760_);
  or (_41762_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41763_, \oc8051_gm_cxrom_1.cell4.data [4], _41737_);
  nand (_41764_, _41763_, _41762_);
  nand (_41765_, _41764_, _41654_);
  or (_41766_, \oc8051_gm_cxrom_1.cell4.data [4], _41654_);
  and (_01617_, _41766_, _41765_);
  or (_41767_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41768_, \oc8051_gm_cxrom_1.cell4.data [5], _41737_);
  nand (_41769_, _41768_, _41767_);
  nand (_41770_, _41769_, _41654_);
  or (_41771_, \oc8051_gm_cxrom_1.cell4.data [5], _41654_);
  and (_01621_, _41771_, _41770_);
  or (_41772_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41773_, \oc8051_gm_cxrom_1.cell4.data [6], _41737_);
  nand (_41774_, _41773_, _41772_);
  nand (_41775_, _41774_, _41654_);
  or (_41776_, \oc8051_gm_cxrom_1.cell4.data [6], _41654_);
  and (_01624_, _41776_, _41775_);
  or (_41777_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_41778_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_41779_, _41778_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_41780_, _41779_, _41777_);
  nand (_41781_, _41780_, _41654_);
  or (_41782_, \oc8051_gm_cxrom_1.cell5.data [7], _41654_);
  and (_01646_, _41782_, _41781_);
  or (_41783_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41784_, \oc8051_gm_cxrom_1.cell5.data [0], _41778_);
  nand (_41785_, _41784_, _41783_);
  nand (_41786_, _41785_, _41654_);
  or (_41787_, \oc8051_gm_cxrom_1.cell5.data [0], _41654_);
  and (_01653_, _41787_, _41786_);
  or (_41788_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41789_, \oc8051_gm_cxrom_1.cell5.data [1], _41778_);
  nand (_41790_, _41789_, _41788_);
  nand (_41791_, _41790_, _41654_);
  or (_41792_, \oc8051_gm_cxrom_1.cell5.data [1], _41654_);
  and (_01657_, _41792_, _41791_);
  or (_41793_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41794_, \oc8051_gm_cxrom_1.cell5.data [2], _41778_);
  nand (_41795_, _41794_, _41793_);
  nand (_41796_, _41795_, _41654_);
  or (_41797_, \oc8051_gm_cxrom_1.cell5.data [2], _41654_);
  and (_01661_, _41797_, _41796_);
  or (_41798_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41799_, \oc8051_gm_cxrom_1.cell5.data [3], _41778_);
  nand (_41800_, _41799_, _41798_);
  nand (_41801_, _41800_, _41654_);
  or (_41802_, \oc8051_gm_cxrom_1.cell5.data [3], _41654_);
  and (_01665_, _41802_, _41801_);
  or (_41803_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41804_, \oc8051_gm_cxrom_1.cell5.data [4], _41778_);
  nand (_41805_, _41804_, _41803_);
  nand (_41806_, _41805_, _41654_);
  or (_41807_, \oc8051_gm_cxrom_1.cell5.data [4], _41654_);
  and (_01668_, _41807_, _41806_);
  or (_41808_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41809_, \oc8051_gm_cxrom_1.cell5.data [5], _41778_);
  nand (_41810_, _41809_, _41808_);
  nand (_41811_, _41810_, _41654_);
  or (_41812_, \oc8051_gm_cxrom_1.cell5.data [5], _41654_);
  and (_01672_, _41812_, _41811_);
  or (_41813_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41814_, \oc8051_gm_cxrom_1.cell5.data [6], _41778_);
  nand (_41815_, _41814_, _41813_);
  nand (_41816_, _41815_, _41654_);
  or (_41817_, \oc8051_gm_cxrom_1.cell5.data [6], _41654_);
  and (_01676_, _41817_, _41816_);
  or (_41818_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_41819_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_41820_, _41819_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_41821_, _41820_, _41818_);
  nand (_41822_, _41821_, _41654_);
  or (_41823_, \oc8051_gm_cxrom_1.cell6.data [7], _41654_);
  and (_01698_, _41823_, _41822_);
  or (_41824_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41825_, \oc8051_gm_cxrom_1.cell6.data [0], _41819_);
  nand (_41826_, _41825_, _41824_);
  nand (_41827_, _41826_, _41654_);
  or (_41828_, \oc8051_gm_cxrom_1.cell6.data [0], _41654_);
  and (_01704_, _41828_, _41827_);
  or (_41829_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41830_, \oc8051_gm_cxrom_1.cell6.data [1], _41819_);
  nand (_41831_, _41830_, _41829_);
  nand (_41832_, _41831_, _41654_);
  or (_41833_, \oc8051_gm_cxrom_1.cell6.data [1], _41654_);
  and (_01708_, _41833_, _41832_);
  or (_41834_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41835_, \oc8051_gm_cxrom_1.cell6.data [2], _41819_);
  nand (_41836_, _41835_, _41834_);
  nand (_41837_, _41836_, _41654_);
  or (_41838_, \oc8051_gm_cxrom_1.cell6.data [2], _41654_);
  and (_01712_, _41838_, _41837_);
  or (_41839_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41840_, \oc8051_gm_cxrom_1.cell6.data [3], _41819_);
  nand (_41841_, _41840_, _41839_);
  nand (_41842_, _41841_, _41654_);
  or (_41843_, \oc8051_gm_cxrom_1.cell6.data [3], _41654_);
  and (_01716_, _41843_, _41842_);
  or (_41844_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41845_, \oc8051_gm_cxrom_1.cell6.data [4], _41819_);
  nand (_41846_, _41845_, _41844_);
  nand (_41847_, _41846_, _41654_);
  or (_41848_, \oc8051_gm_cxrom_1.cell6.data [4], _41654_);
  and (_01720_, _41848_, _41847_);
  or (_41849_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41850_, \oc8051_gm_cxrom_1.cell6.data [5], _41819_);
  nand (_41851_, _41850_, _41849_);
  nand (_41852_, _41851_, _41654_);
  or (_41853_, \oc8051_gm_cxrom_1.cell6.data [5], _41654_);
  and (_01724_, _41853_, _41852_);
  or (_41854_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41855_, \oc8051_gm_cxrom_1.cell6.data [6], _41819_);
  nand (_41856_, _41855_, _41854_);
  nand (_41857_, _41856_, _41654_);
  or (_41858_, \oc8051_gm_cxrom_1.cell6.data [6], _41654_);
  and (_01728_, _41858_, _41857_);
  or (_41859_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_41860_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_41861_, _41860_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_41862_, _41861_, _41859_);
  nand (_41863_, _41862_, _41654_);
  or (_41864_, \oc8051_gm_cxrom_1.cell7.data [7], _41654_);
  and (_01749_, _41864_, _41863_);
  or (_41865_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41866_, \oc8051_gm_cxrom_1.cell7.data [0], _41860_);
  nand (_41867_, _41866_, _41865_);
  nand (_41868_, _41867_, _41654_);
  or (_41869_, \oc8051_gm_cxrom_1.cell7.data [0], _41654_);
  and (_01756_, _41869_, _41868_);
  or (_41870_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41871_, \oc8051_gm_cxrom_1.cell7.data [1], _41860_);
  nand (_41872_, _41871_, _41870_);
  nand (_41873_, _41872_, _41654_);
  or (_41874_, \oc8051_gm_cxrom_1.cell7.data [1], _41654_);
  and (_01760_, _41874_, _41873_);
  or (_41875_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41876_, \oc8051_gm_cxrom_1.cell7.data [2], _41860_);
  nand (_41877_, _41876_, _41875_);
  nand (_41878_, _41877_, _41654_);
  or (_41879_, \oc8051_gm_cxrom_1.cell7.data [2], _41654_);
  and (_01764_, _41879_, _41878_);
  or (_41880_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41881_, \oc8051_gm_cxrom_1.cell7.data [3], _41860_);
  nand (_41882_, _41881_, _41880_);
  nand (_41883_, _41882_, _41654_);
  or (_41884_, \oc8051_gm_cxrom_1.cell7.data [3], _41654_);
  and (_01768_, _41884_, _41883_);
  or (_41885_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41886_, \oc8051_gm_cxrom_1.cell7.data [4], _41860_);
  nand (_41887_, _41886_, _41885_);
  nand (_41888_, _41887_, _41654_);
  or (_41889_, \oc8051_gm_cxrom_1.cell7.data [4], _41654_);
  and (_01772_, _41889_, _41888_);
  or (_41890_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41891_, \oc8051_gm_cxrom_1.cell7.data [5], _41860_);
  nand (_41892_, _41891_, _41890_);
  nand (_41893_, _41892_, _41654_);
  or (_41894_, \oc8051_gm_cxrom_1.cell7.data [5], _41654_);
  and (_01776_, _41894_, _41893_);
  or (_41895_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41896_, \oc8051_gm_cxrom_1.cell7.data [6], _41860_);
  nand (_41897_, _41896_, _41895_);
  nand (_41898_, _41897_, _41654_);
  or (_41899_, \oc8051_gm_cxrom_1.cell7.data [6], _41654_);
  and (_01780_, _41899_, _41898_);
  or (_41900_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_41901_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_41902_, _41901_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_41903_, _41902_, _41900_);
  nand (_41904_, _41903_, _41654_);
  or (_41905_, \oc8051_gm_cxrom_1.cell8.data [7], _41654_);
  and (_01801_, _41905_, _41904_);
  or (_41906_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41907_, \oc8051_gm_cxrom_1.cell8.data [0], _41901_);
  nand (_41908_, _41907_, _41906_);
  nand (_41909_, _41908_, _41654_);
  or (_41910_, \oc8051_gm_cxrom_1.cell8.data [0], _41654_);
  and (_01808_, _41910_, _41909_);
  or (_41911_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41912_, \oc8051_gm_cxrom_1.cell8.data [1], _41901_);
  nand (_41913_, _41912_, _41911_);
  nand (_41914_, _41913_, _41654_);
  or (_41915_, \oc8051_gm_cxrom_1.cell8.data [1], _41654_);
  and (_01812_, _41915_, _41914_);
  or (_41916_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41917_, \oc8051_gm_cxrom_1.cell8.data [2], _41901_);
  nand (_41918_, _41917_, _41916_);
  nand (_41919_, _41918_, _41654_);
  or (_41920_, \oc8051_gm_cxrom_1.cell8.data [2], _41654_);
  and (_01816_, _41920_, _41919_);
  or (_41921_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41922_, \oc8051_gm_cxrom_1.cell8.data [3], _41901_);
  nand (_41923_, _41922_, _41921_);
  nand (_41924_, _41923_, _41654_);
  or (_41925_, \oc8051_gm_cxrom_1.cell8.data [3], _41654_);
  and (_01819_, _41925_, _41924_);
  or (_41926_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41927_, \oc8051_gm_cxrom_1.cell8.data [4], _41901_);
  nand (_41928_, _41927_, _41926_);
  nand (_41929_, _41928_, _41654_);
  or (_41930_, \oc8051_gm_cxrom_1.cell8.data [4], _41654_);
  and (_01823_, _41930_, _41929_);
  or (_41931_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41932_, \oc8051_gm_cxrom_1.cell8.data [5], _41901_);
  nand (_41933_, _41932_, _41931_);
  nand (_41934_, _41933_, _41654_);
  or (_41935_, \oc8051_gm_cxrom_1.cell8.data [5], _41654_);
  and (_01827_, _41935_, _41934_);
  or (_41936_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_41937_, \oc8051_gm_cxrom_1.cell8.data [6], _41901_);
  nand (_41938_, _41937_, _41936_);
  nand (_41939_, _41938_, _41654_);
  or (_41940_, \oc8051_gm_cxrom_1.cell8.data [6], _41654_);
  and (_01831_, _41940_, _41939_);
  or (_41941_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_41942_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_41943_, _41942_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_41944_, _41943_, _41941_);
  nand (_41945_, _41944_, _41654_);
  or (_41946_, \oc8051_gm_cxrom_1.cell9.data [7], _41654_);
  and (_01852_, _41946_, _41945_);
  or (_41947_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41948_, \oc8051_gm_cxrom_1.cell9.data [0], _41942_);
  nand (_41949_, _41948_, _41947_);
  nand (_41950_, _41949_, _41654_);
  or (_41951_, \oc8051_gm_cxrom_1.cell9.data [0], _41654_);
  and (_01859_, _41951_, _41950_);
  or (_41952_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41953_, \oc8051_gm_cxrom_1.cell9.data [1], _41942_);
  nand (_41954_, _41953_, _41952_);
  nand (_41955_, _41954_, _41654_);
  or (_41956_, \oc8051_gm_cxrom_1.cell9.data [1], _41654_);
  and (_01863_, _41956_, _41955_);
  or (_41957_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41958_, \oc8051_gm_cxrom_1.cell9.data [2], _41942_);
  nand (_41959_, _41958_, _41957_);
  nand (_41960_, _41959_, _41654_);
  or (_41961_, \oc8051_gm_cxrom_1.cell9.data [2], _41654_);
  and (_01867_, _41961_, _41960_);
  or (_41962_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41963_, \oc8051_gm_cxrom_1.cell9.data [3], _41942_);
  nand (_41964_, _41963_, _41962_);
  nand (_41965_, _41964_, _41654_);
  or (_41966_, \oc8051_gm_cxrom_1.cell9.data [3], _41654_);
  and (_01871_, _41966_, _41965_);
  or (_41967_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41968_, \oc8051_gm_cxrom_1.cell9.data [4], _41942_);
  nand (_41969_, _41968_, _41967_);
  nand (_41970_, _41969_, _41654_);
  or (_41971_, \oc8051_gm_cxrom_1.cell9.data [4], _41654_);
  and (_01875_, _41971_, _41970_);
  or (_41972_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41973_, \oc8051_gm_cxrom_1.cell9.data [5], _41942_);
  nand (_41974_, _41973_, _41972_);
  nand (_41975_, _41974_, _41654_);
  or (_41976_, \oc8051_gm_cxrom_1.cell9.data [5], _41654_);
  and (_01879_, _41976_, _41975_);
  or (_41977_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_41978_, \oc8051_gm_cxrom_1.cell9.data [6], _41942_);
  nand (_41979_, _41978_, _41977_);
  nand (_41980_, _41979_, _41654_);
  or (_41981_, \oc8051_gm_cxrom_1.cell9.data [6], _41654_);
  and (_01883_, _41981_, _41980_);
  or (_41982_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_41983_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_41984_, _41983_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_41985_, _41984_, _41982_);
  nand (_41986_, _41985_, _41654_);
  or (_41987_, \oc8051_gm_cxrom_1.cell10.data [7], _41654_);
  and (_01892_, _41987_, _41986_);
  or (_41988_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41989_, \oc8051_gm_cxrom_1.cell10.data [0], _41983_);
  nand (_41990_, _41989_, _41988_);
  nand (_41991_, _41990_, _41654_);
  or (_41992_, \oc8051_gm_cxrom_1.cell10.data [0], _41654_);
  and (_01898_, _41992_, _41991_);
  or (_41993_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41994_, \oc8051_gm_cxrom_1.cell10.data [1], _41983_);
  nand (_41995_, _41994_, _41993_);
  nand (_41996_, _41995_, _41654_);
  or (_41997_, \oc8051_gm_cxrom_1.cell10.data [1], _41654_);
  and (_01902_, _41997_, _41996_);
  or (_41998_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_41999_, \oc8051_gm_cxrom_1.cell10.data [2], _41983_);
  nand (_42000_, _41999_, _41998_);
  nand (_42001_, _42000_, _41654_);
  or (_42002_, \oc8051_gm_cxrom_1.cell10.data [2], _41654_);
  and (_01906_, _42002_, _42001_);
  or (_42003_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42004_, \oc8051_gm_cxrom_1.cell10.data [3], _41983_);
  nand (_42005_, _42004_, _42003_);
  nand (_42006_, _42005_, _41654_);
  or (_42007_, \oc8051_gm_cxrom_1.cell10.data [3], _41654_);
  and (_01910_, _42007_, _42006_);
  or (_42008_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42009_, \oc8051_gm_cxrom_1.cell10.data [4], _41983_);
  nand (_42010_, _42009_, _42008_);
  nand (_42011_, _42010_, _41654_);
  or (_42012_, \oc8051_gm_cxrom_1.cell10.data [4], _41654_);
  and (_01914_, _42012_, _42011_);
  or (_42013_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42014_, \oc8051_gm_cxrom_1.cell10.data [5], _41983_);
  nand (_42015_, _42014_, _42013_);
  nand (_42016_, _42015_, _41654_);
  or (_42017_, \oc8051_gm_cxrom_1.cell10.data [5], _41654_);
  and (_01918_, _42017_, _42016_);
  or (_42018_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42019_, \oc8051_gm_cxrom_1.cell10.data [6], _41983_);
  nand (_42020_, _42019_, _42018_);
  nand (_42021_, _42020_, _41654_);
  or (_42022_, \oc8051_gm_cxrom_1.cell10.data [6], _41654_);
  and (_01922_, _42022_, _42021_);
  or (_42023_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_42024_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_42025_, _42024_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_42026_, _42025_, _42023_);
  nand (_42027_, _42026_, _41654_);
  or (_42028_, \oc8051_gm_cxrom_1.cell11.data [7], _41654_);
  and (_01944_, _42028_, _42027_);
  or (_42029_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42030_, \oc8051_gm_cxrom_1.cell11.data [0], _42024_);
  nand (_42031_, _42030_, _42029_);
  nand (_42032_, _42031_, _41654_);
  or (_42033_, \oc8051_gm_cxrom_1.cell11.data [0], _41654_);
  and (_01951_, _42033_, _42032_);
  or (_42034_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42035_, \oc8051_gm_cxrom_1.cell11.data [1], _42024_);
  nand (_42036_, _42035_, _42034_);
  nand (_42037_, _42036_, _41654_);
  or (_42038_, \oc8051_gm_cxrom_1.cell11.data [1], _41654_);
  and (_01955_, _42038_, _42037_);
  or (_42039_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42040_, \oc8051_gm_cxrom_1.cell11.data [2], _42024_);
  nand (_42041_, _42040_, _42039_);
  nand (_42042_, _42041_, _41654_);
  or (_42043_, \oc8051_gm_cxrom_1.cell11.data [2], _41654_);
  and (_01959_, _42043_, _42042_);
  or (_42044_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42045_, \oc8051_gm_cxrom_1.cell11.data [3], _42024_);
  nand (_42046_, _42045_, _42044_);
  nand (_42047_, _42046_, _41654_);
  or (_42048_, \oc8051_gm_cxrom_1.cell11.data [3], _41654_);
  and (_01963_, _42048_, _42047_);
  or (_42049_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42050_, \oc8051_gm_cxrom_1.cell11.data [4], _42024_);
  nand (_42051_, _42050_, _42049_);
  nand (_42052_, _42051_, _41654_);
  or (_42053_, \oc8051_gm_cxrom_1.cell11.data [4], _41654_);
  and (_01967_, _42053_, _42052_);
  or (_42054_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42055_, \oc8051_gm_cxrom_1.cell11.data [5], _42024_);
  nand (_42056_, _42055_, _42054_);
  nand (_42057_, _42056_, _41654_);
  or (_42058_, \oc8051_gm_cxrom_1.cell11.data [5], _41654_);
  and (_01971_, _42058_, _42057_);
  or (_42059_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42060_, \oc8051_gm_cxrom_1.cell11.data [6], _42024_);
  nand (_42061_, _42060_, _42059_);
  nand (_42062_, _42061_, _41654_);
  or (_42063_, \oc8051_gm_cxrom_1.cell11.data [6], _41654_);
  and (_01975_, _42063_, _42062_);
  or (_42064_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_42065_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_42066_, _42065_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_42067_, _42066_, _42064_);
  nand (_42068_, _42067_, _41654_);
  or (_42069_, \oc8051_gm_cxrom_1.cell12.data [7], _41654_);
  and (_01997_, _42069_, _42068_);
  or (_42070_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42071_, \oc8051_gm_cxrom_1.cell12.data [0], _42065_);
  nand (_42072_, _42071_, _42070_);
  nand (_42073_, _42072_, _41654_);
  or (_42074_, \oc8051_gm_cxrom_1.cell12.data [0], _41654_);
  and (_02004_, _42074_, _42073_);
  or (_42075_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42076_, \oc8051_gm_cxrom_1.cell12.data [1], _42065_);
  nand (_42077_, _42076_, _42075_);
  nand (_42078_, _42077_, _41654_);
  or (_42079_, \oc8051_gm_cxrom_1.cell12.data [1], _41654_);
  and (_02007_, _42079_, _42078_);
  or (_42080_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42081_, \oc8051_gm_cxrom_1.cell12.data [2], _42065_);
  nand (_42082_, _42081_, _42080_);
  nand (_42083_, _42082_, _41654_);
  or (_42084_, \oc8051_gm_cxrom_1.cell12.data [2], _41654_);
  and (_02011_, _42084_, _42083_);
  or (_42085_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42086_, \oc8051_gm_cxrom_1.cell12.data [3], _42065_);
  nand (_42087_, _42086_, _42085_);
  nand (_42088_, _42087_, _41654_);
  or (_42089_, \oc8051_gm_cxrom_1.cell12.data [3], _41654_);
  and (_02015_, _42089_, _42088_);
  or (_42090_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42091_, \oc8051_gm_cxrom_1.cell12.data [4], _42065_);
  nand (_42092_, _42091_, _42090_);
  nand (_42093_, _42092_, _41654_);
  or (_42094_, \oc8051_gm_cxrom_1.cell12.data [4], _41654_);
  and (_02019_, _42094_, _42093_);
  or (_42095_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42096_, \oc8051_gm_cxrom_1.cell12.data [5], _42065_);
  nand (_42097_, _42096_, _42095_);
  nand (_42098_, _42097_, _41654_);
  or (_42099_, \oc8051_gm_cxrom_1.cell12.data [5], _41654_);
  and (_02023_, _42099_, _42098_);
  or (_42100_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42101_, \oc8051_gm_cxrom_1.cell12.data [6], _42065_);
  nand (_42102_, _42101_, _42100_);
  nand (_42103_, _42102_, _41654_);
  or (_42104_, \oc8051_gm_cxrom_1.cell12.data [6], _41654_);
  and (_02027_, _42104_, _42103_);
  or (_42105_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_42106_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_42107_, _42106_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_42108_, _42107_, _42105_);
  nand (_42109_, _42108_, _41654_);
  or (_42110_, \oc8051_gm_cxrom_1.cell13.data [7], _41654_);
  and (_02048_, _42110_, _42109_);
  or (_42111_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42112_, \oc8051_gm_cxrom_1.cell13.data [0], _42106_);
  nand (_42113_, _42112_, _42111_);
  nand (_42114_, _42113_, _41654_);
  or (_42115_, \oc8051_gm_cxrom_1.cell13.data [0], _41654_);
  and (_02055_, _42115_, _42114_);
  or (_42116_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42117_, \oc8051_gm_cxrom_1.cell13.data [1], _42106_);
  nand (_42118_, _42117_, _42116_);
  nand (_42119_, _42118_, _41654_);
  or (_42120_, \oc8051_gm_cxrom_1.cell13.data [1], _41654_);
  and (_02059_, _42120_, _42119_);
  or (_42121_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42122_, \oc8051_gm_cxrom_1.cell13.data [2], _42106_);
  nand (_42123_, _42122_, _42121_);
  nand (_42124_, _42123_, _41654_);
  or (_42125_, \oc8051_gm_cxrom_1.cell13.data [2], _41654_);
  and (_02063_, _42125_, _42124_);
  or (_42126_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42127_, \oc8051_gm_cxrom_1.cell13.data [3], _42106_);
  nand (_42128_, _42127_, _42126_);
  nand (_42129_, _42128_, _41654_);
  or (_42130_, \oc8051_gm_cxrom_1.cell13.data [3], _41654_);
  and (_02067_, _42130_, _42129_);
  or (_42131_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42132_, \oc8051_gm_cxrom_1.cell13.data [4], _42106_);
  nand (_42133_, _42132_, _42131_);
  nand (_42134_, _42133_, _41654_);
  or (_42135_, \oc8051_gm_cxrom_1.cell13.data [4], _41654_);
  and (_02071_, _42135_, _42134_);
  or (_42136_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42137_, \oc8051_gm_cxrom_1.cell13.data [5], _42106_);
  nand (_42138_, _42137_, _42136_);
  nand (_42139_, _42138_, _41654_);
  or (_42140_, \oc8051_gm_cxrom_1.cell13.data [5], _41654_);
  and (_02075_, _42140_, _42139_);
  or (_42141_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42142_, \oc8051_gm_cxrom_1.cell13.data [6], _42106_);
  nand (_42143_, _42142_, _42141_);
  nand (_42144_, _42143_, _41654_);
  or (_42145_, \oc8051_gm_cxrom_1.cell13.data [6], _41654_);
  and (_02079_, _42145_, _42144_);
  or (_42146_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_42147_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_42148_, _42147_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_42149_, _42148_, _42146_);
  nand (_42150_, _42149_, _41654_);
  or (_42151_, \oc8051_gm_cxrom_1.cell14.data [7], _41654_);
  and (_02100_, _42151_, _42150_);
  or (_42152_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42153_, \oc8051_gm_cxrom_1.cell14.data [0], _42147_);
  nand (_42154_, _42153_, _42152_);
  nand (_42155_, _42154_, _41654_);
  or (_42156_, \oc8051_gm_cxrom_1.cell14.data [0], _41654_);
  and (_02107_, _42156_, _42155_);
  or (_42157_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42158_, \oc8051_gm_cxrom_1.cell14.data [1], _42147_);
  nand (_42159_, _42158_, _42157_);
  nand (_42160_, _42159_, _41654_);
  or (_42161_, \oc8051_gm_cxrom_1.cell14.data [1], _41654_);
  and (_02111_, _42161_, _42160_);
  or (_42162_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42163_, \oc8051_gm_cxrom_1.cell14.data [2], _42147_);
  nand (_42164_, _42163_, _42162_);
  nand (_42165_, _42164_, _41654_);
  or (_42166_, \oc8051_gm_cxrom_1.cell14.data [2], _41654_);
  and (_02115_, _42166_, _42165_);
  or (_42167_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42168_, \oc8051_gm_cxrom_1.cell14.data [3], _42147_);
  nand (_42169_, _42168_, _42167_);
  nand (_42170_, _42169_, _41654_);
  or (_42171_, \oc8051_gm_cxrom_1.cell14.data [3], _41654_);
  and (_02118_, _42171_, _42170_);
  or (_42172_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42173_, \oc8051_gm_cxrom_1.cell14.data [4], _42147_);
  nand (_42174_, _42173_, _42172_);
  nand (_42175_, _42174_, _41654_);
  or (_42176_, \oc8051_gm_cxrom_1.cell14.data [4], _41654_);
  and (_02122_, _42176_, _42175_);
  or (_42177_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42178_, \oc8051_gm_cxrom_1.cell14.data [5], _42147_);
  nand (_42179_, _42178_, _42177_);
  nand (_42180_, _42179_, _41654_);
  or (_42181_, \oc8051_gm_cxrom_1.cell14.data [5], _41654_);
  and (_02126_, _42181_, _42180_);
  or (_42182_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42183_, \oc8051_gm_cxrom_1.cell14.data [6], _42147_);
  nand (_42184_, _42183_, _42182_);
  nand (_42185_, _42184_, _41654_);
  or (_42186_, \oc8051_gm_cxrom_1.cell14.data [6], _41654_);
  and (_02130_, _42186_, _42185_);
  or (_42187_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_42188_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_42189_, _42188_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_42190_, _42189_, _42187_);
  nand (_42191_, _42190_, _41654_);
  or (_42192_, \oc8051_gm_cxrom_1.cell15.data [7], _41654_);
  and (_02152_, _42192_, _42191_);
  or (_42193_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42194_, \oc8051_gm_cxrom_1.cell15.data [0], _42188_);
  nand (_42195_, _42194_, _42193_);
  nand (_42196_, _42195_, _41654_);
  or (_42197_, \oc8051_gm_cxrom_1.cell15.data [0], _41654_);
  and (_02159_, _42197_, _42196_);
  or (_42198_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42199_, \oc8051_gm_cxrom_1.cell15.data [1], _42188_);
  nand (_42200_, _42199_, _42198_);
  nand (_42201_, _42200_, _41654_);
  or (_42202_, \oc8051_gm_cxrom_1.cell15.data [1], _41654_);
  and (_02163_, _42202_, _42201_);
  or (_42203_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42204_, \oc8051_gm_cxrom_1.cell15.data [2], _42188_);
  nand (_42205_, _42204_, _42203_);
  nand (_42206_, _42205_, _41654_);
  or (_42207_, \oc8051_gm_cxrom_1.cell15.data [2], _41654_);
  and (_02167_, _42207_, _42206_);
  or (_42208_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42209_, \oc8051_gm_cxrom_1.cell15.data [3], _42188_);
  nand (_42210_, _42209_, _42208_);
  nand (_42211_, _42210_, _41654_);
  or (_42212_, \oc8051_gm_cxrom_1.cell15.data [3], _41654_);
  and (_02171_, _42212_, _42211_);
  or (_42213_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42214_, \oc8051_gm_cxrom_1.cell15.data [4], _42188_);
  nand (_42215_, _42214_, _42213_);
  nand (_42216_, _42215_, _41654_);
  or (_42217_, \oc8051_gm_cxrom_1.cell15.data [4], _41654_);
  and (_02174_, _42217_, _42216_);
  or (_42218_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42219_, \oc8051_gm_cxrom_1.cell15.data [5], _42188_);
  nand (_42220_, _42219_, _42218_);
  nand (_42221_, _42220_, _41654_);
  or (_42222_, \oc8051_gm_cxrom_1.cell15.data [5], _41654_);
  and (_02178_, _42222_, _42221_);
  or (_42223_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42224_, \oc8051_gm_cxrom_1.cell15.data [6], _42188_);
  nand (_42225_, _42224_, _42223_);
  nand (_42226_, _42225_, _41654_);
  or (_42227_, \oc8051_gm_cxrom_1.cell15.data [6], _41654_);
  and (_02182_, _42227_, _42226_);
  nor (_05950_, _38210_, rst);
  and (_42228_, _34293_, _41654_);
  nand (_42229_, _42228_, _37058_);
  nor (_42230_, _36796_, _36742_);
  or (_05953_, _42230_, _42229_);
  and (_42231_, _35678_, _35446_);
  and (_42232_, _42231_, _35931_);
  and (_42233_, _42232_, _36677_);
  and (_42234_, _35157_, _34664_);
  and (_42235_, _36184_, _34915_);
  and (_42236_, _42235_, _42234_);
  and (_42237_, _42236_, _42233_);
  not (_42238_, _36677_);
  nor (_42239_, _36184_, _34915_);
  not (_42240_, _35157_);
  and (_42241_, _42240_, _34664_);
  and (_42242_, _42241_, _42239_);
  nor (_42243_, _42242_, _42238_);
  not (_42244_, _35446_);
  and (_42245_, _35931_, _35678_);
  and (_42246_, _42245_, _42244_);
  not (_42247_, _42246_);
  nor (_42248_, _42247_, _42243_);
  not (_42249_, _42248_);
  and (_42250_, _36677_, _42244_);
  and (_42251_, _42250_, _42245_);
  not (_42252_, _36184_);
  nor (_42253_, _42252_, _34915_);
  and (_42254_, _42253_, _42234_);
  and (_42255_, _42254_, _42251_);
  and (_42256_, _42252_, _34915_);
  and (_42257_, _42256_, _42241_);
  and (_42258_, _42257_, _42251_);
  nor (_42259_, _42258_, _42255_);
  and (_42260_, _42259_, _42249_);
  and (_42261_, _42241_, _36184_);
  and (_42262_, _42261_, _42251_);
  nor (_42263_, _35157_, _34664_);
  and (_42264_, _42263_, _42235_);
  not (_42265_, _35678_);
  and (_42266_, _35931_, _42265_);
  and (_42267_, _42266_, _42244_);
  and (_42268_, _42267_, _42238_);
  and (_42269_, _42268_, _42264_);
  not (_42270_, _34915_);
  and (_42271_, _42263_, _42270_);
  and (_42272_, _42271_, _42251_);
  or (_42273_, _42272_, _42269_);
  nor (_42274_, _42273_, _42262_);
  nand (_42275_, _42274_, _42260_);
  or (_42276_, _42275_, _42237_);
  not (_42277_, _34664_);
  and (_42278_, _35157_, _42277_);
  and (_42279_, _42266_, _42250_);
  and (_42280_, _42279_, _42252_);
  and (_42281_, _42280_, _42278_);
  not (_42282_, _42251_);
  and (_42283_, _42239_, _42234_);
  nor (_42284_, _42283_, _42236_);
  nor (_42285_, _42284_, _42282_);
  not (_42286_, _42285_);
  and (_42287_, _42278_, _42256_);
  and (_42288_, _42287_, _42251_);
  and (_42289_, _42278_, _42253_);
  not (_42290_, _35931_);
  and (_42291_, _42265_, _35446_);
  nor (_42292_, _42291_, _42290_);
  not (_42293_, _42292_);
  and (_42294_, _42293_, _42289_);
  nor (_42295_, _42294_, _42288_);
  nand (_42296_, _42295_, _42286_);
  or (_42297_, _42296_, _42281_);
  and (_42298_, _42278_, _34915_);
  and (_42299_, _42232_, _42238_);
  and (_42300_, _42299_, _42298_);
  and (_42301_, _42264_, _42290_);
  or (_42302_, _42301_, _42300_);
  and (_42303_, _42253_, _42241_);
  and (_42304_, _42299_, _42303_);
  and (_42305_, _42289_, _42267_);
  or (_42306_, _42305_, _42304_);
  or (_42307_, _42306_, _42302_);
  and (_42308_, _42271_, _42232_);
  nand (_42309_, _42233_, _42234_);
  nor (_42310_, _42235_, _42309_);
  or (_42311_, _42310_, _42308_);
  or (_42312_, _42311_, _42307_);
  or (_42313_, _42312_, _42297_);
  or (_42314_, _42313_, _42276_);
  and (_42315_, _42314_, _34304_);
  not (_42316_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_42317_, _34282_, _16098_);
  and (_42318_, _42317_, _37189_);
  nor (_42319_, _42318_, _42316_);
  or (_42320_, _42319_, rst);
  or (_05956_, _42320_, _42315_);
  nand (_42321_, _34664_, _34238_);
  or (_42322_, _34238_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_42323_, _42322_, _41654_);
  and (_05959_, _42323_, _42321_);
  and (_42324_, \oc8051_top_1.oc8051_sfr1.wait_data , _41654_);
  and (_42325_, _42324_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_42326_, _36873_, _36446_);
  and (_42327_, _38200_, _37331_);
  or (_42328_, _42327_, _42326_);
  and (_42329_, _36742_, _36446_);
  or (_42330_, _42329_, _38171_);
  or (_42331_, _42330_, _37755_);
  and (_42332_, _37546_, _36873_);
  and (_42333_, _36796_, _36764_);
  or (_42334_, _42333_, _42332_);
  nor (_42335_, _42334_, _42331_);
  nand (_42336_, _42335_, _38030_);
  or (_42337_, _42336_, _42328_);
  and (_42338_, _42337_, _42228_);
  or (_05962_, _42338_, _42325_);
  and (_42339_, _36916_, _36742_);
  or (_42340_, _42339_, _36895_);
  and (_42341_, _37458_, _36753_);
  or (_42342_, _42341_, _37091_);
  and (_42343_, _37298_, _35491_);
  and (_42344_, _42343_, _37546_);
  or (_42345_, _42344_, _42342_);
  or (_42346_, _42345_, _42340_);
  and (_42347_, _42346_, _34293_);
  and (_42348_, \oc8051_top_1.oc8051_decoder1.state [0], _16098_);
  and (_42349_, _42348_, _42316_);
  not (_42350_, _38203_);
  and (_42351_, _42350_, _42349_);
  and (_42352_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42353_, _42352_, _42351_);
  or (_42354_, _42353_, _42347_);
  and (_05965_, _42354_, _41654_);
  and (_42355_, _42324_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_42356_, _38200_, _37480_);
  nor (_42357_, _37480_, _36764_);
  nor (_42358_, _42357_, _37419_);
  or (_42359_, _42358_, _42356_);
  and (_42360_, _42343_, _37777_);
  or (_42361_, _42360_, _42359_);
  nor (_42362_, _42357_, _35975_);
  not (_42363_, _35975_);
  and (_42364_, _37777_, _42363_);
  or (_42365_, _42364_, _42362_);
  or (_42366_, _42365_, _36425_);
  nor (_42367_, _36228_, _35975_);
  and (_42368_, _42367_, _36392_);
  and (_42369_, _38200_, _37353_);
  or (_42370_, _42369_, _42368_);
  or (_42371_, _42370_, _42340_);
  or (_42372_, _42371_, _42366_);
  or (_42373_, _42372_, _42361_);
  and (_42374_, _42373_, _42228_);
  or (_05968_, _42374_, _42355_);
  and (_42375_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42376_, _37931_, _34293_);
  or (_42377_, _42376_, _42375_);
  or (_42378_, _42377_, _42351_);
  and (_05971_, _42378_, _41654_);
  and (_42379_, _36873_, _36436_);
  not (_42380_, _37331_);
  nor (_42381_, _42230_, _42380_);
  nor (_42382_, _42381_, _42379_);
  not (_42383_, _42382_);
  and (_42384_, _42383_, _42349_);
  and (_42385_, _36807_, _37777_);
  and (_42386_, _37309_, _36479_);
  and (_42387_, _42386_, _36239_);
  or (_42388_, _42387_, _42385_);
  or (_42389_, _42388_, _42326_);
  and (_42390_, _42389_, _38207_);
  or (_42391_, _42390_, _42384_);
  and (_42392_, _42388_, _37205_);
  or (_42393_, _42392_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42394_, _42393_, _42391_);
  or (_42395_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _16098_);
  and (_42396_, _42395_, _41654_);
  and (_05974_, _42396_, _42394_);
  and (_42397_, _42324_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_42398_, _42364_, _36895_);
  and (_42399_, _36764_, _42363_);
  or (_42400_, _42399_, _37799_);
  or (_42401_, _42400_, _42398_);
  and (_42402_, _37546_, _36283_);
  or (_42403_, _42333_, _37744_);
  or (_42404_, _42403_, _42402_);
  or (_42405_, _42341_, _37557_);
  and (_42406_, _36348_, _36261_);
  or (_42407_, _42360_, _42406_);
  or (_42408_, _42407_, _37579_);
  or (_42409_, _42408_, _42405_);
  or (_42410_, _42409_, _42404_);
  or (_42411_, _42410_, _42401_);
  and (_42412_, _42411_, _42228_);
  or (_05977_, _42412_, _42397_);
  and (_42413_, _42324_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_42414_, _42344_, _37832_);
  and (_42415_, _36873_, _36294_);
  and (_42416_, _42343_, _37004_);
  or (_42417_, _42416_, _42415_);
  or (_42418_, _42417_, _42414_);
  or (_42419_, _42418_, _42365_);
  and (_42420_, _38200_, _37656_);
  and (_42421_, _37656_, _36796_);
  or (_42422_, _37843_, _42421_);
  or (_42423_, _42422_, _42420_);
  and (_42424_, _37036_, _35212_);
  or (_42425_, _42424_, _37014_);
  and (_42426_, _36764_, _36283_);
  or (_42427_, _42426_, _42425_);
  or (_42428_, _42427_, _42423_);
  or (_42429_, _42428_, _42419_);
  and (_42430_, _37458_, _35212_);
  and (_42431_, _37458_, _36949_);
  or (_42432_, _42431_, _42430_);
  nor (_42433_, _38052_, _36359_);
  nand (_42434_, _42433_, _37678_);
  or (_42435_, _42434_, _42432_);
  or (_42436_, _42435_, _42361_);
  or (_42437_, _42436_, _42429_);
  and (_42438_, _42437_, _42228_);
  or (_05980_, _42438_, _42413_);
  and (_42439_, _42367_, _36436_);
  or (_42440_, _42439_, _36316_);
  and (_42441_, _42343_, _36305_);
  and (_42442_, _36305_, _42363_);
  or (_42443_, _42442_, _37102_);
  or (_42444_, _42443_, _42441_);
  or (_42445_, _42444_, _42440_);
  and (_42446_, _42343_, _36916_);
  or (_42447_, _42446_, _42445_);
  and (_42448_, _42447_, _34293_);
  and (_42449_, _38202_, _16098_);
  and (_42450_, _38201_, _16098_);
  or (_42451_, _42450_, _42449_);
  and (_42452_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_42453_, _42452_, _42451_);
  or (_42454_, _42453_, _42448_);
  and (_05983_, _42454_, _41654_);
  or (_42455_, _37590_, _37557_);
  not (_42456_, _38063_);
  or (_42457_, _42358_, _42456_);
  or (_42458_, _42457_, _42455_);
  and (_42459_, _36938_, _36239_);
  and (_42460_, _42459_, _37320_);
  or (_42461_, _42460_, _37788_);
  or (_42462_, _42461_, _42421_);
  or (_42463_, _42462_, _42385_);
  nand (_42464_, _37942_, _37766_);
  or (_42465_, _42464_, _42463_);
  or (_42466_, _42465_, _42458_);
  and (_42467_, _36446_, _42363_);
  and (_42468_, _42367_, _36938_);
  or (_42469_, _42468_, _37469_);
  or (_42470_, _42469_, _42467_);
  or (_42471_, _42470_, _42342_);
  and (_42472_, _42459_, _36283_);
  or (_42473_, _42472_, _36359_);
  or (_42474_, _42473_, _37265_);
  or (_42475_, _42387_, _36457_);
  or (_42476_, _42475_, _37898_);
  or (_42477_, _42476_, _42474_);
  or (_42478_, _42477_, _42471_);
  or (_42479_, _42478_, _42365_);
  or (_42480_, _42479_, _42466_);
  and (_42481_, _42480_, _34293_);
  and (_42482_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42483_, _42392_, _42351_);
  and (_42484_, _38189_, _37205_);
  or (_42485_, _42484_, _42483_);
  or (_42486_, _42485_, _42482_);
  or (_42487_, _42486_, _42481_);
  and (_05986_, _42487_, _41654_);
  nor (_06045_, _37251_, rst);
  nor (_06047_, _38195_, rst);
  nand (_06050_, _42383_, _42228_);
  and (_42488_, _37058_, _36742_);
  or (_42489_, _42488_, _42379_);
  nand (_06053_, _42489_, _42228_);
  and (_42490_, _42234_, _42270_);
  and (_42491_, _42490_, _42233_);
  or (_42492_, _42300_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_42493_, _42492_, _42491_);
  or (_42494_, _42493_, _42281_);
  and (_42495_, _42494_, _42318_);
  nor (_42496_, _42317_, _37189_);
  or (_42497_, _42496_, rst);
  or (_06056_, _42497_, _42495_);
  nand (_42498_, _36677_, _34238_);
  or (_42499_, _34238_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_42500_, _42499_, _41654_);
  and (_06059_, _42500_, _42498_);
  not (_42501_, _34238_);
  or (_42502_, _35446_, _42501_);
  or (_42503_, _34238_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_42504_, _42503_, _41654_);
  and (_06062_, _42504_, _42502_);
  nand (_42505_, _35678_, _34238_);
  or (_42506_, _34238_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_42507_, _42506_, _41654_);
  and (_06065_, _42507_, _42505_);
  nand (_42508_, _35931_, _34238_);
  or (_42509_, _34238_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_42510_, _42509_, _41654_);
  and (_06068_, _42510_, _42508_);
  or (_42511_, _36184_, _42501_);
  or (_42512_, _34238_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_42513_, _42512_, _41654_);
  and (_06071_, _42513_, _42511_);
  nand (_42514_, _34915_, _34238_);
  or (_42515_, _34238_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_42516_, _42515_, _41654_);
  and (_06074_, _42516_, _42514_);
  nand (_42517_, _35157_, _34238_);
  or (_42518_, _34238_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_42519_, _42518_, _41654_);
  and (_06077_, _42519_, _42517_);
  and (_42520_, _42430_, _34707_);
  or (_42521_, _42441_, _37102_);
  or (_42522_, _42521_, _42520_);
  or (_42523_, _37080_, _36895_);
  or (_42524_, _42523_, _42522_);
  and (_42525_, _42343_, _37656_);
  or (_42526_, _42525_, _42339_);
  or (_42527_, _36764_, _36348_);
  and (_42528_, _42527_, _38200_);
  or (_42529_, _42528_, _42526_);
  or (_42530_, _42529_, _42524_);
  or (_42531_, _42431_, _42416_);
  and (_42532_, _38200_, _36960_);
  or (_42533_, _42532_, _42440_);
  or (_42534_, _42533_, _42531_);
  or (_42535_, _37342_, _37014_);
  or (_42536_, _42415_, _42327_);
  or (_42537_, _42536_, _42535_);
  or (_42538_, _42537_, _42534_);
  nor (_42539_, _37408_, _35975_);
  or (_42540_, _42539_, _42446_);
  and (_42541_, _42343_, _37397_);
  or (_42542_, _42541_, _36272_);
  and (_42543_, _37058_, _36239_);
  and (_42544_, _42543_, _38200_);
  and (_42545_, _37458_, _37058_);
  or (_42546_, _42545_, _42544_);
  or (_42547_, _42546_, _42542_);
  or (_42548_, _42547_, _42540_);
  or (_42549_, _42548_, _42538_);
  or (_42550_, _42549_, _42530_);
  and (_42551_, _42550_, _34293_);
  and (_42552_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42553_, _42552_, _42384_);
  or (_42554_, _42553_, _42551_);
  and (_30380_, _42554_, _41654_);
  and (_42555_, _42324_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_42556_, _37656_, _37004_);
  and (_42557_, _42556_, _36807_);
  or (_42558_, _42526_, _42432_);
  or (_42559_, _42558_, _42557_);
  nor (_42560_, _42368_, _36403_);
  not (_42561_, _42560_);
  nor (_42562_, _42561_, _42369_);
  nand (_42563_, _42562_, _37568_);
  or (_42564_, _42563_, _42328_);
  not (_42565_, _37004_);
  nand (_42566_, _42565_, _37408_);
  and (_42567_, _42566_, _38200_);
  or (_42568_, _42567_, _42427_);
  or (_42569_, _42568_, _42564_);
  or (_42570_, _42569_, _42559_);
  and (_42572_, _42570_, _42228_);
  or (_30383_, _42572_, _42555_);
  or (_42575_, _42476_, _42467_);
  or (_42577_, _42575_, _42466_);
  and (_42579_, _42577_, _34293_);
  and (_42581_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42583_, _42581_, _42485_);
  or (_42585_, _42583_, _42579_);
  and (_30385_, _42585_, _41654_);
  and (_42588_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42590_, _38041_, _36228_);
  or (_42592_, _42590_, _37091_);
  or (_42594_, _42592_, _42474_);
  or (_42596_, _42594_, _42388_);
  and (_42598_, _42596_, _34293_);
  or (_42600_, _42598_, _42588_);
  or (_42602_, _42600_, _42483_);
  and (_30387_, _42602_, _41654_);
  or (_42605_, _42439_, _36326_);
  or (_42607_, _42605_, _42388_);
  or (_42609_, _42379_, _38202_);
  and (_42611_, _42441_, _36239_);
  or (_42613_, _42611_, _42541_);
  or (_42615_, _42613_, _42609_);
  or (_42617_, _42556_, _36960_);
  and (_42619_, _42617_, _38200_);
  or (_42621_, _42619_, _42615_);
  or (_42623_, _42621_, _42607_);
  and (_42625_, _38200_, _37546_);
  or (_42627_, _42415_, _42625_);
  or (_42629_, _42627_, _42540_);
  and (_42630_, _42343_, _37733_);
  or (_42631_, _42630_, _42327_);
  or (_42632_, _42544_, _38201_);
  or (_42633_, _42632_, _42528_);
  or (_42634_, _42633_, _42631_);
  and (_42635_, _42441_, _36228_);
  or (_42636_, _42635_, _36971_);
  or (_42637_, _42472_, _37102_);
  or (_42638_, _42637_, _42468_);
  and (_42639_, _36807_, _37397_);
  and (_42640_, _42543_, _37320_);
  or (_42641_, _42640_, _42639_);
  or (_42642_, _42641_, _42638_);
  or (_42643_, _42642_, _42636_);
  or (_42644_, _42643_, _42634_);
  or (_42645_, _42644_, _42629_);
  or (_42646_, _42645_, _42623_);
  and (_42647_, _42646_, _34293_);
  and (_42648_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42649_, _42384_, _38208_);
  or (_42650_, _42649_, _42648_);
  or (_42651_, _42650_, _42647_);
  and (_30389_, _42651_, _41654_);
  or (_42652_, _38202_, _37102_);
  or (_42653_, _42460_, _42339_);
  or (_42654_, _42653_, _42652_);
  or (_42655_, _35733_, _42363_);
  and (_42656_, _42655_, _42543_);
  or (_42657_, _42656_, _37898_);
  or (_42658_, _42657_, _42654_);
  nand (_42659_, _37436_, _36982_);
  or (_42660_, _42659_, _42658_);
  or (_42661_, _38052_, _42421_);
  and (_42662_, _42661_, _36862_);
  or (_42663_, _42662_, _42605_);
  or (_42664_, _42663_, _42660_);
  or (_42665_, _42634_, _42629_);
  or (_42666_, _42665_, _42664_);
  and (_42667_, _42666_, _34293_);
  and (_42668_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42669_, _42668_, _42649_);
  or (_42670_, _42669_, _42667_);
  and (_30391_, _42670_, _41654_);
  and (_42671_, _42324_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_42672_, _40180_);
  or (_42673_, _42446_, _42672_);
  and (_42674_, _36873_, _36348_);
  and (_42675_, _42674_, _36239_);
  and (_42676_, _42333_, _36862_);
  or (_42677_, _42676_, _42675_);
  or (_42678_, _42677_, _42401_);
  or (_42679_, _42678_, _42673_);
  and (_42680_, _37997_, _42363_);
  or (_42681_, _37102_, _42406_);
  nor (_42682_, _42681_, _42680_);
  nand (_42683_, _42682_, _40179_);
  and (_42684_, _38200_, _36764_);
  or (_42685_, _42684_, _42360_);
  or (_42686_, _42685_, _42455_);
  or (_42687_, _42686_, _42683_);
  and (_42688_, _37997_, _36873_);
  and (_42689_, _36873_, _37733_);
  and (_42690_, _36316_, _36239_);
  or (_42691_, _42690_, _42689_);
  or (_42692_, _42691_, _42688_);
  or (_42693_, _42439_, _42341_);
  or (_42694_, _42693_, _42611_);
  or (_42695_, _42402_, _37920_);
  or (_42696_, _42695_, _42694_);
  or (_42697_, _42696_, _42692_);
  or (_42698_, _42697_, _42687_);
  or (_42699_, _42698_, _42679_);
  and (_42700_, _42699_, _42228_);
  or (_30393_, _42700_, _42671_);
  or (_42701_, _42344_, _37667_);
  or (_42702_, _42426_, _42424_);
  or (_42703_, _42702_, _42701_);
  or (_42704_, _42703_, _42423_);
  or (_42705_, _42704_, _42615_);
  or (_42706_, _42684_, _42688_);
  or (_42708_, _42675_, _42636_);
  or (_42709_, _42708_, _42706_);
  or (_42710_, _42430_, _36895_);
  or (_42711_, _42710_, _36326_);
  not (_42712_, _37909_);
  or (_42713_, _42539_, _42712_);
  or (_42714_, _42713_, _42711_);
  or (_42715_, _42714_, _42709_);
  or (_42716_, _42715_, _42705_);
  and (_42717_, _42716_, _42228_);
  and (_42718_, _42324_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_42720_, _34249_, _41654_);
  and (_42721_, _42720_, _38202_);
  or (_42722_, _42721_, _42718_);
  or (_30395_, _42722_, _42717_);
  or (_42723_, _42368_, _37645_);
  or (_42724_, _42723_, _42446_);
  or (_42725_, _42724_, _42631_);
  and (_42726_, _42367_, _35223_);
  or (_42727_, _42726_, _36272_);
  and (_42728_, _36796_, _37733_);
  or (_42729_, _42728_, _42544_);
  or (_42730_, _42729_, _42727_);
  or (_42731_, _42730_, _42725_);
  nor (_42732_, _42541_, _37898_);
  not (_42733_, _42732_);
  nor (_42734_, _42733_, _37887_);
  or (_42735_, _42344_, _37124_);
  and (_42736_, _36873_, _36305_);
  or (_42737_, _42693_, _42736_);
  nor (_42738_, _42737_, _42735_);
  nand (_42739_, _42738_, _42734_);
  or (_42740_, _42739_, _42731_);
  or (_42741_, _42366_, _42361_);
  or (_42742_, _42741_, _42740_);
  and (_42743_, _42742_, _34293_);
  and (_42744_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42745_, _42744_, _42449_);
  or (_42746_, _42745_, _42743_);
  and (_30397_, _42746_, _41654_);
  or (_42747_, _42733_, _42727_);
  or (_42748_, _42747_, _42729_);
  or (_42749_, _37091_, _36359_);
  nor (_42750_, _42749_, _42674_);
  nand (_42751_, _42750_, _40180_);
  or (_42752_, _42685_, _42405_);
  or (_42753_, _42752_, _42751_);
  or (_42754_, _42365_, _42359_);
  or (_42755_, _42754_, _42753_);
  or (_42756_, _42755_, _42748_);
  and (_42757_, _42756_, _34293_);
  and (_42758_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42759_, _42758_, _42450_);
  or (_42760_, _42759_, _42757_);
  and (_30399_, _42760_, _41654_);
  and (_42761_, _42324_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_42762_, _42630_, _37579_);
  nand (_42763_, _42762_, _40179_);
  or (_42764_, _42763_, _42706_);
  or (_42765_, _42561_, _42332_);
  or (_42766_, _42765_, _42689_);
  or (_42767_, _42766_, _42445_);
  or (_42768_, _42677_, _42673_);
  or (_42769_, _42768_, _42767_);
  or (_42770_, _42769_, _42764_);
  and (_42771_, _42770_, _42228_);
  or (_30401_, _42771_, _42761_);
  nor (_38625_, _34664_, rst);
  nor (_38627_, _40137_, rst);
  and (_42772_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_42773_, _34347_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_42774_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_42775_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_42776_, _42775_, _42774_);
  and (_42777_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_42778_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_42779_, _42778_, _42777_);
  and (_42780_, _42779_, _42776_);
  and (_42781_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_42782_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_42783_, _42782_, _42781_);
  and (_42784_, _42783_, _42780_);
  nor (_42785_, _42784_, _34347_);
  nor (_42786_, _42785_, _42773_);
  nor (_42787_, _42786_, _40121_);
  nor (_42788_, _42787_, _42772_);
  nor (_38628_, _42788_, rst);
  nor (_38639_, _36677_, rst);
  and (_38640_, _35446_, _41654_);
  nor (_38641_, _35678_, rst);
  nor (_38642_, _35931_, rst);
  and (_38643_, _36184_, _41654_);
  nor (_38644_, _34915_, rst);
  nor (_38645_, _35157_, rst);
  nor (_38646_, _40332_, rst);
  nor (_38648_, _40485_, rst);
  nor (_38649_, _40251_, rst);
  nor (_38650_, _40295_, rst);
  nor (_38651_, _40423_, rst);
  nor (_38652_, _40206_, rst);
  nor (_38654_, _40388_, rst);
  and (_42789_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_42790_, _34347_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_42791_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42792_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42793_, _42792_, _42791_);
  and (_42794_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_42795_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_42796_, _42795_, _42794_);
  and (_42797_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_42798_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_42799_, _42798_, _42797_);
  and (_42800_, _42799_, _42796_);
  and (_42801_, _42800_, _42793_);
  nor (_42802_, _42801_, _34347_);
  nor (_42803_, _42802_, _42790_);
  nor (_42804_, _42803_, _40121_);
  nor (_42805_, _42804_, _42789_);
  nor (_38655_, _42805_, rst);
  and (_42806_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_42807_, _34347_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_42808_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_42809_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_42810_, _42809_, _42808_);
  and (_42811_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_42812_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_42813_, _42812_, _42811_);
  and (_42814_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42815_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_42816_, _42815_, _42814_);
  and (_42817_, _42816_, _42813_);
  and (_42818_, _42817_, _42810_);
  nor (_42819_, _42818_, _34347_);
  nor (_42820_, _42819_, _42807_);
  nor (_42821_, _42820_, _40121_);
  nor (_42822_, _42821_, _42806_);
  nor (_38656_, _42822_, rst);
  and (_42823_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_42824_, _34347_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_42825_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_42826_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_42827_, _42826_, _42825_);
  and (_42828_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_42829_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_42830_, _42829_, _42828_);
  and (_42831_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_42832_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_42833_, _42832_, _42831_);
  and (_42834_, _42833_, _42830_);
  and (_42835_, _42834_, _42827_);
  nor (_42836_, _42835_, _34347_);
  nor (_42837_, _42836_, _42824_);
  nor (_42838_, _42837_, _40121_);
  nor (_42839_, _42838_, _42823_);
  nor (_38657_, _42839_, rst);
  and (_42840_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_42841_, _34347_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_42842_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_42843_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_42844_, _42843_, _42842_);
  and (_42845_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_42846_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_42847_, _42846_, _42845_);
  and (_42848_, _42847_, _42844_);
  and (_42849_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_42850_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_42851_, _42850_, _42849_);
  and (_42852_, _42851_, _42848_);
  nor (_42853_, _42852_, _34347_);
  nor (_42854_, _42853_, _42841_);
  nor (_42855_, _42854_, _40121_);
  nor (_42856_, _42855_, _42840_);
  nor (_38658_, _42856_, rst);
  and (_42857_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_42858_, _34347_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_42859_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_42860_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_42861_, _42860_, _42859_);
  and (_42862_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42863_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_42864_, _42863_, _42862_);
  and (_42865_, _42864_, _42861_);
  and (_42866_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_42867_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_42868_, _42867_, _42866_);
  and (_42869_, _42868_, _42865_);
  nor (_42870_, _42869_, _34347_);
  nor (_42871_, _42870_, _42858_);
  nor (_42872_, _42871_, _40121_);
  nor (_42873_, _42872_, _42857_);
  nor (_38660_, _42873_, rst);
  and (_42874_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_42875_, _34347_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_42876_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_42877_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_42878_, _42877_, _42876_);
  and (_42879_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42880_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_42881_, _42880_, _42879_);
  and (_42882_, _42881_, _42878_);
  and (_42883_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_42884_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_42885_, _42884_, _42883_);
  and (_42886_, _42885_, _42882_);
  nor (_42887_, _42886_, _34347_);
  nor (_42888_, _42887_, _42875_);
  nor (_42889_, _42888_, _40121_);
  nor (_42890_, _42889_, _42874_);
  nor (_38661_, _42890_, rst);
  and (_42891_, _40121_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_42892_, _34347_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_42893_, _34478_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_42894_, _34434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_42895_, _42894_, _42893_);
  and (_42896_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42897_, _34522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_42898_, _42897_, _42896_);
  and (_42899_, _42898_, _42895_);
  and (_42900_, _34391_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_42901_, _34555_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42902_, _42901_, _42900_);
  and (_42903_, _42902_, _42899_);
  nor (_42904_, _42903_, _34347_);
  nor (_42905_, _42904_, _42892_);
  nor (_42906_, _42905_, _40121_);
  nor (_42907_, _42906_, _42891_);
  nor (_38662_, _42907_, rst);
  and (_42908_, _34304_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_42909_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_42910_, _42908_, _38435_);
  and (_42911_, _42910_, _41654_);
  and (_38685_, _42911_, _42909_);
  not (_42912_, _42908_);
  or (_42913_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _42908_, _41654_);
  and (_42914_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _41654_);
  or (_42915_, _42914_, _00000_);
  and (_38687_, _42915_, _42913_);
  nor (_38720_, _40176_, rst);
  and (_38722_, _40448_, _41654_);
  nor (_38723_, _40171_, rst);
  nor (_42916_, _40315_, _25548_);
  and (_42917_, _40315_, _25548_);
  nor (_42918_, _42917_, _42916_);
  not (_42919_, _42918_);
  and (_42920_, _40396_, _38758_);
  nor (_42921_, _40396_, _38758_);
  and (_42922_, _40232_, _38882_);
  or (_42923_, _42922_, _42921_);
  or (_42924_, _42923_, _42920_);
  and (_42925_, _40176_, _25406_);
  nor (_42926_, _40176_, _25406_);
  and (_42927_, _40466_, _25678_);
  nor (_42928_, _40466_, _25678_);
  nor (_42929_, _42928_, _42927_);
  nor (_42930_, _40232_, _38882_);
  not (_42931_, _42930_);
  nand (_42932_, _42931_, _42929_);
  or (_42933_, _42932_, _42926_);
  or (_42934_, _42933_, _42925_);
  nor (_42935_, _42934_, _42924_);
  and (_42936_, _42935_, _42919_);
  nor (_42937_, _38030_, _42348_);
  and (_42938_, _38708_, _28541_);
  and (_42939_, _42938_, _42937_);
  and (_42940_, _42939_, _42936_);
  or (_42941_, _26435_, _26083_);
  nor (_42942_, _42941_, _29483_);
  and (_42943_, _42942_, _30676_);
  nand (_42944_, _42943_, _31298_);
  nor (_42945_, _42944_, _32007_);
  nor (_42946_, _42937_, _38182_);
  and (_42947_, _42946_, _42945_);
  and (_42948_, _42947_, _33542_);
  and (_42949_, _42948_, _27060_);
  and (_42950_, _42937_, _26808_);
  not (_42951_, _38182_);
  nor (_42952_, _42937_, _34959_);
  nor (_42953_, _42952_, _42951_);
  and (_42954_, _42953_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_42955_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_42956_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_42957_, _42956_, _42955_);
  nor (_42958_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_42959_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_42960_, _42959_, _42958_);
  and (_42961_, _42960_, _42957_);
  and (_42962_, _42961_, _37220_);
  or (_42963_, _42962_, _42954_);
  or (_42964_, _42963_, _42950_);
  nor (_42965_, _42964_, _42949_);
  not (_42966_, _42399_);
  nor (_42967_, _42630_, _37799_);
  and (_42968_, _42967_, _42966_);
  or (_42969_, _37997_, _36960_);
  nor (_42970_, _42969_, _37397_);
  nor (_42971_, _42970_, _37986_);
  nor (_42972_, _42971_, _42561_);
  and (_42973_, _42972_, _42968_);
  not (_42975_, _42973_);
  and (_42976_, _42975_, _42965_);
  not (_42977_, _42976_);
  and (_42978_, _38171_, _36228_);
  not (_42979_, _42978_);
  and (_42981_, _42979_, _38190_);
  nor (_42982_, _42981_, _42965_);
  nor (_42983_, _42329_, _36971_);
  not (_42984_, _42983_);
  nor (_42985_, _42984_, _42982_);
  and (_42987_, _42985_, _42977_);
  nor (_42988_, _42987_, _38186_);
  and (_42989_, _36807_, _36348_);
  nor (_42990_, _42989_, _42386_);
  nor (_42991_, _42990_, _34249_);
  nor (_42993_, _42991_, _37228_);
  not (_42994_, _42993_);
  nor (_42995_, _42994_, _42988_);
  nor (_42996_, _38762_, _38715_);
  and (_42997_, _42996_, _38741_);
  not (_42999_, _42997_);
  and (_43000_, _42999_, _42953_);
  not (_43001_, _38941_);
  and (_43002_, _43001_, _37220_);
  nor (_43003_, _43002_, _43000_);
  not (_43005_, _43003_);
  nor (_43006_, _43005_, _42995_);
  not (_43007_, _43006_);
  nor (_43008_, _43007_, _42940_);
  nor (_43009_, _42918_, _38999_);
  and (_43011_, _40548_, _31103_);
  nor (_43012_, _40548_, _31103_);
  or (_43014_, _43012_, _43011_);
  or (_43015_, _40351_, _24884_);
  nand (_43016_, _40351_, _24884_);
  and (_43017_, _43016_, _43015_);
  or (_43018_, _40271_, _24645_);
  nand (_43019_, _40271_, _24645_);
  and (_43020_, _43019_, _43018_);
  or (_43022_, _43020_, _43017_);
  nor (_43023_, _43022_, _43014_);
  and (_43024_, _43023_, _43009_);
  and (_43026_, _43024_, _42935_);
  nor (_43027_, _25395_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_43028_, _43027_, _43026_);
  not (_43030_, _43028_);
  and (_43031_, _43030_, _43008_);
  nor (_43032_, _37235_, rst);
  and (_38727_, _43032_, _43031_);
  and (_38728_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _41654_);
  and (_38729_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _41654_);
  and (_43035_, _37235_, _28475_);
  and (_43036_, _37205_, _36971_);
  not (_43037_, _43036_);
  nor (_43039_, _43037_, _38446_);
  and (_43040_, _42560_, _38030_);
  and (_43041_, _43040_, _42967_);
  nor (_43043_, _43041_, _38186_);
  and (_43044_, _42989_, _38207_);
  nor (_43046_, _43044_, _38138_);
  not (_43047_, _43046_);
  nor (_43048_, _43047_, _43043_);
  and (_43049_, _43048_, _42991_);
  and (_43050_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43051_, _43050_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_43052_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43054_, _43052_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_43055_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43056_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_43058_, _43056_, _43055_);
  and (_43059_, _43058_, _43054_);
  and (_43060_, _43059_, _43051_);
  and (_43062_, _43060_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43063_, _43062_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43064_, _43063_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_43066_, _43064_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43067_, _43066_, _38435_);
  or (_43068_, _43066_, _38435_);
  and (_43070_, _43068_, _43067_);
  and (_43071_, _43070_, _43049_);
  nor (_43072_, _43036_, _42991_);
  nand (_43074_, _43048_, _43072_);
  nor (_43075_, _42984_, _38171_);
  and (_43076_, _43075_, _42968_);
  and (_43078_, _43076_, _43040_);
  nor (_43079_, _43078_, _38186_);
  and (_43081_, _37964_, _38207_);
  or (_43082_, _43081_, _43079_);
  nor (_43083_, _43082_, _43074_);
  and (_43084_, _43083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43085_, _43044_, _40138_);
  or (_43087_, _43085_, _43084_);
  or (_43088_, _43087_, _43071_);
  nor (_43089_, _43088_, _43039_);
  nand (_43091_, _43089_, _43031_);
  or (_43092_, _43091_, _43035_);
  and (_43093_, _36742_, _38207_);
  and (_43095_, _43093_, _36305_);
  not (_43096_, _43095_);
  and (_43097_, _43048_, _43096_);
  and (_43099_, _43097_, _40137_);
  not (_43100_, _42788_);
  nor (_43101_, _43097_, _43100_);
  nor (_43103_, _43101_, _43099_);
  and (_43104_, _43103_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_43105_, _43103_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_43107_, _43097_, _40388_);
  not (_43108_, _42907_);
  nor (_43109_, _43097_, _43108_);
  nor (_43111_, _43109_, _43107_);
  and (_43112_, _43111_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_43114_, _43111_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_43115_, _43114_, _43112_);
  and (_43116_, _43097_, _40206_);
  not (_43117_, _42890_);
  nor (_43118_, _43097_, _43117_);
  nor (_43119_, _43118_, _43116_);
  and (_43120_, _43119_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_43122_, _43119_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_43123_, _43097_, _40423_);
  not (_43124_, _42873_);
  nor (_43126_, _43097_, _43124_);
  nor (_43127_, _43126_, _43123_);
  nand (_43128_, _43127_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43130_, _43097_, _40295_);
  not (_43131_, _42856_);
  nor (_43132_, _43097_, _43131_);
  nor (_43134_, _43132_, _43130_);
  and (_43135_, _43134_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_43148_, _43134_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_43153_, _43097_, _40251_);
  not (_43154_, _42839_);
  nor (_43168_, _43097_, _43154_);
  nor (_43173_, _43168_, _43153_);
  and (_43174_, _43173_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43186_, _43097_, _40485_);
  not (_43193_, _42822_);
  nor (_43194_, _43097_, _43193_);
  nor (_43205_, _43194_, _43186_);
  and (_43206_, _43205_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_43214_, _43097_, _40332_);
  not (_43222_, _42805_);
  nor (_43231_, _43097_, _43222_);
  nor (_43232_, _43231_, _43214_);
  and (_43241_, _43232_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_43249_, _43205_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_43250_, _43249_, _43206_);
  and (_43261_, _43250_, _43241_);
  nor (_43267_, _43261_, _43206_);
  not (_43268_, _43267_);
  nor (_43280_, _43173_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_43286_, _43280_, _43174_);
  and (_43287_, _43286_, _43268_);
  nor (_43300_, _43287_, _43174_);
  nor (_43305_, _43300_, _43148_);
  or (_43306_, _43305_, _43135_);
  or (_43320_, _43127_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43325_, _43320_, _43128_);
  nand (_43326_, _43325_, _43306_);
  and (_43338_, _43326_, _43128_);
  nor (_43345_, _43338_, _43122_);
  or (_43346_, _43345_, _43120_);
  and (_43357_, _43346_, _43115_);
  nor (_43358_, _43357_, _43112_);
  nor (_43366_, _43358_, _43105_);
  or (_43374_, _43366_, _43104_);
  and (_43376_, _43374_, _43051_);
  and (_43377_, _43376_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43378_, _43377_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43380_, _43378_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_43381_, _43380_, _43103_);
  not (_43382_, _43103_);
  nor (_43384_, _43374_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43385_, _43384_, _38413_);
  and (_43386_, _43385_, _38418_);
  and (_43388_, _43386_, _38403_);
  nor (_43389_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43390_, _43389_, _43388_);
  nor (_43392_, _43390_, _43382_);
  nor (_43393_, _43392_, _43381_);
  or (_43394_, _43103_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43396_, _43103_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_43397_, _43396_, _43394_);
  and (_43398_, _43397_, _43393_);
  or (_43400_, _43398_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_43401_, _43398_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_43403_, _43401_, _43400_);
  not (_43404_, _43072_);
  and (_43405_, _43097_, _43404_);
  nor (_43406_, _43095_, _43079_);
  nor (_43408_, _43406_, _43405_);
  and (_43409_, _43408_, _43403_);
  or (_43410_, _43409_, _43092_);
  not (_43412_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_43414_, _43413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_43416_, _43414_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_43417_, _43416_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_43418_, _43417_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_43420_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_43421_, _43420_, _43418_);
  and (_43422_, _43421_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_43424_, _43422_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_43425_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_43426_, _34467_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43428_, _43426_, _40121_);
  nor (_43429_, _43428_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_43430_, _43429_);
  and (_43432_, _43430_, _43425_);
  and (_43433_, _43432_, _43424_);
  nand (_43435_, _43433_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_43436_, _43435_, _43412_);
  or (_43437_, _43435_, _43412_);
  and (_43438_, _43437_, _43436_);
  or (_43439_, _43438_, _43031_);
  and (_43440_, _43439_, _41654_);
  and (_38731_, _43440_, _43410_);
  and (_43442_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _41654_);
  and (_43443_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_43444_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_43446_, _34293_, _43444_);
  not (_43447_, _43446_);
  not (_43448_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_43450_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_43451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_43452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_43454_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_43455_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_43456_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_43458_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_43459_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_43460_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_43462_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43463_, _43462_, _43460_);
  and (_43464_, _43463_, _43459_);
  and (_43466_, _43464_, _43458_);
  and (_43467_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_43469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_43470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43471_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_43472_, _43471_, _43469_);
  and (_43474_, _43472_, _43470_);
  nor (_43475_, _43474_, _43469_);
  nor (_43476_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43478_, _43476_, _43467_);
  not (_43479_, _43478_);
  nor (_43480_, _43479_, _43475_);
  nor (_43482_, _43480_, _43467_);
  and (_43483_, _43482_, _43466_);
  and (_43484_, _43483_, _43456_);
  and (_43486_, _43484_, _43455_);
  and (_43487_, _43486_, _43454_);
  and (_43488_, _43487_, _43452_);
  and (_43490_, _43488_, _43451_);
  and (_43491_, _43490_, _43450_);
  and (_43492_, _43491_, _43448_);
  nor (_43494_, _43492_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43495_, _43492_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_43496_, _43495_, _43494_);
  nor (_43498_, _43491_, _43448_);
  nor (_43499_, _43498_, _43492_);
  not (_43501_, _43499_);
  nor (_43502_, _43490_, _43450_);
  or (_43503_, _43502_, _43491_);
  nor (_43504_, _43488_, _43451_);
  nor (_43506_, _43504_, _43490_);
  not (_43507_, _43506_);
  nor (_43508_, _43487_, _43452_);
  or (_43510_, _43508_, _43488_);
  nor (_43511_, _43486_, _43454_);
  nor (_43512_, _43511_, _43487_);
  not (_43514_, _43512_);
  nor (_43515_, _43484_, _43455_);
  nor (_43516_, _43515_, _43486_);
  not (_43518_, _43516_);
  and (_43519_, _43482_, _43463_);
  and (_43520_, _43519_, _43459_);
  nor (_43522_, _43520_, _43458_);
  or (_43523_, _43522_, _43483_);
  nor (_43524_, _43519_, _43459_);
  nor (_43526_, _43524_, _43520_);
  not (_43527_, _43526_);
  and (_43528_, _43482_, _43462_);
  nor (_43530_, _43528_, _43460_);
  nor (_43531_, _43530_, _43519_);
  not (_43533_, _43531_);
  not (_43534_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43535_, _43482_, _43534_);
  nor (_43536_, _43482_, _43534_);
  nor (_43538_, _43536_, _43535_);
  not (_43539_, _43538_);
  and (_43540_, _42242_, _42232_);
  nor (_43542_, _42279_, _42233_);
  not (_43543_, _42257_);
  not (_43544_, _42233_);
  nor (_43546_, _42264_, _42303_);
  or (_43547_, _43546_, _43544_);
  and (_43548_, _43547_, _43543_);
  nor (_43550_, _43548_, _43542_);
  nor (_43551_, _43550_, _43540_);
  not (_43552_, _42267_);
  and (_43554_, _42278_, _42235_);
  nor (_43555_, _43554_, _42242_);
  nor (_43556_, _43555_, _43552_);
  or (_43558_, _42301_, _42288_);
  nor (_43559_, _43558_, _42262_);
  nand (_43560_, _43559_, _42260_);
  nor (_43562_, _43560_, _43556_);
  and (_43563_, _43562_, _43551_);
  not (_43565_, _42268_);
  nor (_43566_, _42287_, _42303_);
  nor (_43567_, _43566_, _43565_);
  not (_43568_, _43567_);
  and (_43569_, _42268_, _42490_);
  and (_43571_, _42263_, _42256_);
  nor (_43572_, _43571_, _42289_);
  nor (_43573_, _43572_, _43544_);
  nor (_43575_, _43573_, _43569_);
  and (_43576_, _42289_, _42268_);
  and (_43577_, _42241_, _42235_);
  and (_43579_, _42299_, _43577_);
  nor (_43580_, _43579_, _43576_);
  and (_43581_, _42234_, _34915_);
  nand (_43583_, _42268_, _43581_);
  and (_43584_, _43583_, _43580_);
  and (_43585_, _43584_, _43575_);
  and (_43587_, _42278_, _42239_);
  or (_43588_, _43554_, _43587_);
  nand (_43589_, _43588_, _42233_);
  and (_43591_, _43581_, _42233_);
  and (_43592_, _42263_, _42253_);
  or (_43593_, _43592_, _42257_);
  and (_43595_, _43593_, _42268_);
  nor (_43596_, _43595_, _43591_);
  and (_43598_, _43596_, _43589_);
  and (_43599_, _43598_, _43585_);
  and (_43600_, _43599_, _43568_);
  and (_43601_, _43600_, _43563_);
  and (_43603_, _42279_, _42303_);
  and (_43604_, _42289_, _42251_);
  nor (_43605_, _43604_, _43603_);
  and (_43607_, _42263_, _42239_);
  and (_43608_, _43607_, _42268_);
  and (_43609_, _43554_, _42251_);
  nor (_43611_, _43609_, _43608_);
  and (_43612_, _43611_, _43605_);
  and (_43613_, _42299_, _42257_);
  and (_43615_, _43571_, _42268_);
  or (_43616_, _43615_, _43613_);
  nor (_43617_, _43616_, _42294_);
  and (_43619_, _43617_, _43612_);
  not (_43620_, _43587_);
  and (_43621_, _43566_, _43620_);
  nor (_43623_, _43621_, _35931_);
  and (_43624_, _42252_, _35931_);
  and (_43625_, _42291_, _42278_);
  and (_43627_, _43625_, _43624_);
  nor (_43628_, _43627_, _43623_);
  and (_43630_, _42289_, _42279_);
  not (_43631_, _43630_);
  nor (_43632_, _42285_, _42269_);
  and (_43633_, _43632_, _43631_);
  not (_43635_, _43577_);
  nor (_43636_, _42267_, _42233_);
  nor (_43637_, _43636_, _43635_);
  and (_43639_, _42263_, _34915_);
  nor (_43640_, _43587_, _43639_);
  nor (_43641_, _43640_, _42282_);
  nor (_43643_, _43641_, _43637_);
  and (_43644_, _43643_, _43633_);
  and (_43645_, _42280_, _42490_);
  and (_43647_, _42279_, _42254_);
  and (_43648_, _42287_, _42233_);
  and (_43649_, _36184_, _35931_);
  and (_43651_, _42241_, _42270_);
  and (_43652_, _42291_, _43651_);
  and (_43653_, _43652_, _43649_);
  or (_43655_, _43653_, _43648_);
  or (_43656_, _43655_, _43647_);
  nor (_43657_, _43656_, _43645_);
  and (_43659_, _43657_, _43644_);
  and (_43660_, _43659_, _43628_);
  and (_43662_, _43660_, _43619_);
  and (_43663_, _43662_, _43601_);
  nor (_43664_, _43472_, _43470_);
  nor (_43665_, _43664_, _43474_);
  not (_43667_, _43665_);
  nor (_43668_, _43667_, _43663_);
  and (_43669_, _43580_, _43633_);
  nor (_43671_, _42294_, _43591_);
  and (_43672_, _43671_, _43568_);
  nor (_43673_, _43613_, _42255_);
  and (_43675_, _42299_, _42242_);
  nor (_43676_, _43609_, _43675_);
  and (_43677_, _43676_, _43673_);
  and (_43679_, _43677_, _43672_);
  and (_43680_, _43679_, _43669_);
  not (_43681_, _43680_);
  nor (_43683_, _43681_, _43663_);
  not (_43684_, _43683_);
  nor (_43685_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43687_, _43685_, _43470_);
  and (_43688_, _43687_, _43684_);
  and (_43689_, _43667_, _43663_);
  nor (_43691_, _43689_, _43668_);
  and (_43692_, _43691_, _43688_);
  nor (_43693_, _43692_, _43668_);
  not (_43694_, _43693_);
  and (_43695_, _43479_, _43475_);
  nor (_43696_, _43695_, _43480_);
  and (_43697_, _43696_, _43694_);
  and (_43698_, _43697_, _43539_);
  not (_43699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_43700_, _43535_, _43699_);
  or (_43701_, _43700_, _43528_);
  and (_43702_, _43701_, _43698_);
  and (_43703_, _43702_, _43533_);
  and (_43704_, _43703_, _43527_);
  and (_43705_, _43704_, _43523_);
  nor (_43706_, _43483_, _43456_);
  or (_43707_, _43706_, _43484_);
  and (_43708_, _43707_, _43705_);
  and (_43709_, _43708_, _43518_);
  and (_43710_, _43709_, _43514_);
  and (_43711_, _43710_, _43510_);
  and (_43712_, _43711_, _43507_);
  and (_43713_, _43712_, _43503_);
  and (_43714_, _43713_, _43501_);
  or (_43715_, _43714_, _43496_);
  nand (_43716_, _43714_, _43496_);
  and (_43717_, _43716_, _43715_);
  or (_43718_, _43717_, _43447_);
  or (_43719_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_43720_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_43721_, _43720_, _43719_);
  and (_43722_, _43721_, _43718_);
  or (_38732_, _43722_, _43443_);
  nor (_43723_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_38733_, _43723_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_38734_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _41654_);
  nor (_43724_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_43725_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_43726_, _43725_, _43724_);
  nor (_43727_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_43728_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_43729_, _43728_, _43727_);
  and (_43730_, _43729_, _43726_);
  nor (_43731_, _43730_, rst);
  and (_43732_, \oc8051_top_1.oc8051_rom1.ea_int , _34260_);
  nand (_43733_, _43732_, _34293_);
  and (_43734_, _43733_, _38734_);
  or (_38735_, _43734_, _43731_);
  and (_43735_, _43730_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_43736_, _43735_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_38736_, _43736_, _41654_);
  nor (_43737_, _43429_, _40121_);
  nor (_43738_, _43663_, _34413_);
  nor (_43739_, _43683_, _34500_);
  and (_43740_, _43663_, _34413_);
  nor (_43741_, _43740_, _43738_);
  and (_43742_, _43741_, _43739_);
  nor (_43743_, _43742_, _43738_);
  nor (_43744_, _43743_, _40121_);
  and (_43745_, _43744_, _34369_);
  nor (_43746_, _43744_, _34369_);
  nor (_43747_, _43746_, _43745_);
  nor (_43748_, _43747_, _43737_);
  and (_43749_, _34424_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_43750_, _43749_, _43737_);
  nor (_43751_, _43750_, _43680_);
  or (_43752_, _43751_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_43753_, _43752_, _43748_);
  and (_38737_, _43753_, _41654_);
  not (_43754_, _35366_);
  and (_43755_, _34620_, _43754_);
  not (_43756_, _36118_);
  and (_43757_, _43756_, _35113_);
  and (_43758_, _43757_, _43755_);
  and (_43759_, _34304_, _41654_);
  nand (_43760_, _43759_, _35634_);
  nor (_43761_, _43760_, _35887_);
  not (_43762_, _34871_);
  nor (_43763_, _36633_, _43762_);
  and (_43764_, _43763_, _43761_);
  and (_38740_, _43764_, _43758_);
  nor (_43765_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_43766_, _43765_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_43767_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_38743_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _41654_);
  and (_43768_, _38743_, _43767_);
  or (_38742_, _43768_, _43766_);
  not (_43769_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_43770_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43771_, _43770_, _43769_);
  and (_43772_, _43770_, _43769_);
  nor (_43773_, _43772_, _43771_);
  not (_43774_, _43773_);
  and (_43775_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_43776_, _43775_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43777_, _43775_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43778_, _43777_, _43776_);
  or (_43779_, _43778_, _43770_);
  and (_43780_, _43779_, _43774_);
  nor (_43781_, _43771_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_43782_, _43771_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_43783_, _43782_, _43781_);
  or (_43784_, _43776_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_38745_, _43784_, _41654_);
  and (_43785_, _38745_, _43783_);
  and (_38744_, _43785_, _43780_);
  not (_43786_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_43787_, _43429_, _43786_);
  and (_43788_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_43789_, _43787_);
  and (_43790_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_43791_, _43790_, _43788_);
  and (_38746_, _43791_, _41654_);
  and (_43792_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_43793_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_43794_, _43793_, _43792_);
  and (_38747_, _43794_, _41654_);
  and (_43795_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_43796_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_43797_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _43796_);
  and (_43798_, _43797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_43799_, _43798_, _43795_);
  and (_38749_, _43799_, _41654_);
  and (_43800_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_43801_, _43800_, _43797_);
  and (_38750_, _43801_, _41654_);
  or (_43802_, _43796_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_38751_, _43802_, _41654_);
  not (_43803_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_43804_, _43803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_43805_, _43804_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_43806_, _43796_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_43807_, _43806_, _41654_);
  and (_38752_, _43807_, _43805_);
  or (_43808_, _43796_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_38753_, _43808_, _41654_);
  nor (_43809_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_43810_, _43809_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_43811_, _43810_, _41654_);
  and (_43812_, _38743_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_38754_, _43812_, _43811_);
  and (_43813_, _43786_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_43814_, _43813_, _43810_);
  and (_38755_, _43814_, _41654_);
  nand (_43815_, _43810_, _38446_);
  or (_43816_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_43817_, _43816_, _41654_);
  and (_38756_, _43817_, _43815_);
  and (_38757_, _38213_, _40119_);
  or (_43818_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_43819_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_43820_, _42908_, _43819_);
  and (_43821_, _43820_, _41654_);
  and (_38795_, _43821_, _43818_);
  or (_43822_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_43823_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_43824_, _42908_, _43823_);
  and (_43825_, _43824_, _41654_);
  and (_38796_, _43825_, _43822_);
  or (_43826_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_43827_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_43828_, _42908_, _43827_);
  and (_43829_, _43828_, _41654_);
  and (_38797_, _43829_, _43826_);
  or (_43830_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_43831_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_43832_, _42908_, _43831_);
  and (_43833_, _43832_, _41654_);
  and (_38799_, _43833_, _43830_);
  or (_43834_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43835_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4], _41654_);
  or (_43836_, _43835_, _00000_);
  and (_38800_, _43836_, _43834_);
  or (_43837_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_43838_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_43839_, _42908_, _43838_);
  and (_43840_, _43839_, _41654_);
  and (_38801_, _43840_, _43837_);
  or (_43841_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_43842_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6], _41654_);
  or (_43843_, _43842_, _00000_);
  and (_38802_, _43843_, _43841_);
  or (_43844_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_43845_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_43846_, _42908_, _43845_);
  and (_43847_, _43846_, _41654_);
  and (_38803_, _43847_, _43844_);
  or (_43848_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_43849_, _42908_, _38407_);
  and (_43850_, _43849_, _41654_);
  and (_38804_, _43850_, _43848_);
  or (_43851_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_43852_, _42908_, _38413_);
  and (_43853_, _43852_, _41654_);
  and (_38805_, _43853_, _43851_);
  or (_43854_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_43855_, _42908_, _38418_);
  and (_43856_, _43855_, _41654_);
  and (_38806_, _43856_, _43854_);
  or (_43857_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_43858_, _42908_, _38403_);
  and (_43859_, _43858_, _41654_);
  and (_38807_, _43859_, _43857_);
  or (_43860_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_43861_, _42908_, _38424_);
  and (_43862_, _43861_, _41654_);
  and (_38808_, _43862_, _43860_);
  or (_43863_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_43864_, _42908_, _38399_);
  and (_43865_, _43864_, _41654_);
  and (_38810_, _43865_, _43863_);
  or (_43866_, _42908_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_43867_, _42908_, _38430_);
  and (_43868_, _43867_, _41654_);
  and (_38811_, _43868_, _43866_);
  or (_43869_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_43870_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _41654_);
  or (_43871_, _43870_, _00000_);
  and (_38815_, _43871_, _43869_);
  or (_43872_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_43873_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _41654_);
  or (_43874_, _43873_, _00000_);
  and (_38816_, _43874_, _43872_);
  or (_43875_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_43876_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _41654_);
  or (_43877_, _43876_, _00000_);
  and (_38817_, _43877_, _43875_);
  or (_43878_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_43879_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _41654_);
  or (_43880_, _43879_, _00000_);
  and (_38818_, _43880_, _43878_);
  or (_43881_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_43882_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _41654_);
  or (_43883_, _43882_, _00000_);
  and (_38819_, _43883_, _43881_);
  or (_43884_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_43885_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _41654_);
  or (_43886_, _43885_, _00000_);
  and (_38820_, _43886_, _43884_);
  or (_43887_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_43888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _41654_);
  or (_43889_, _43888_, _00000_);
  and (_38821_, _43889_, _43887_);
  or (_43890_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_43891_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _41654_);
  or (_43892_, _43891_, _00000_);
  and (_38822_, _43892_, _43890_);
  or (_43893_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_43894_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _41654_);
  or (_43895_, _43894_, _00000_);
  and (_38824_, _43895_, _43893_);
  or (_43896_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_43897_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _41654_);
  or (_43898_, _43897_, _00000_);
  and (_38825_, _43898_, _43896_);
  or (_43899_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_43900_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _41654_);
  or (_43901_, _43900_, _00000_);
  and (_38826_, _43901_, _43899_);
  or (_43902_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_43903_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _41654_);
  or (_43904_, _43903_, _00000_);
  and (_38827_, _43904_, _43902_);
  or (_43905_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_43906_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _41654_);
  or (_43907_, _43906_, _00000_);
  and (_38828_, _43907_, _43905_);
  or (_43908_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_43909_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _41654_);
  or (_43910_, _43909_, _00000_);
  and (_38829_, _43910_, _43908_);
  or (_00006_, _42912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_00007_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _41654_);
  or (_00008_, _00007_, _00000_);
  and (_38830_, _00008_, _00006_);
  nor (_39005_, _36720_, rst);
  nor (_39006_, _35491_, rst);
  nor (_39007_, _35722_, rst);
  nor (_39008_, _40152_, rst);
  and (_00009_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00010_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_00011_, _00010_, _00009_);
  and (_39009_, _00011_, _41654_);
  and (_00012_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00013_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00014_, _00013_, _43787_);
  or (_00015_, _00014_, _00012_);
  and (_39010_, _00015_, _41654_);
  and (_00016_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00017_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_00018_, _00017_, _00016_);
  and (_39012_, _00018_, _41654_);
  and (_00019_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00020_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_00021_, _00020_, _43787_);
  or (_00022_, _00021_, _00019_);
  and (_39013_, _00022_, _41654_);
  and (_00023_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00024_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_00025_, _00024_, _00023_);
  and (_39014_, _00025_, _41654_);
  and (_00026_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00027_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_00028_, _00027_, _00026_);
  and (_39015_, _00028_, _41654_);
  and (_00029_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00030_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_00031_, _00030_, _00029_);
  and (_39016_, _00031_, _41654_);
  and (_00032_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00033_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_00034_, _00033_, _00032_);
  and (_39017_, _00034_, _41654_);
  and (_00035_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_00036_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_00037_, _00036_, _00035_);
  and (_39018_, _00037_, _41654_);
  and (_00038_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_00039_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_00040_, _00039_, _00038_);
  and (_39019_, _00040_, _41654_);
  and (_00041_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_00042_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_00043_, _00042_, _00041_);
  and (_39020_, _00043_, _41654_);
  and (_00044_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_00045_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_00046_, _00045_, _00044_);
  and (_39021_, _00046_, _41654_);
  and (_00047_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_00048_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_00049_, _00048_, _00047_);
  and (_39023_, _00049_, _41654_);
  and (_00050_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_00051_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_00052_, _00051_, _00050_);
  and (_39024_, _00052_, _41654_);
  and (_00053_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_00054_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_00055_, _00054_, _00053_);
  and (_39025_, _00055_, _41654_);
  and (_00056_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_00057_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_00058_, _00057_, _00056_);
  and (_39026_, _00058_, _41654_);
  and (_00059_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_00060_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_00061_, _00060_, _00059_);
  and (_39027_, _00061_, _41654_);
  and (_00062_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_00063_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_00064_, _00063_, _00062_);
  and (_39028_, _00064_, _41654_);
  and (_00065_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_00066_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_00067_, _00066_, _00065_);
  and (_39029_, _00067_, _41654_);
  and (_00068_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_00069_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_00070_, _00069_, _00068_);
  and (_39030_, _00070_, _41654_);
  and (_00071_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_00072_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_00073_, _00072_, _00071_);
  and (_39031_, _00073_, _41654_);
  and (_00074_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_00075_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_00076_, _00075_, _00074_);
  and (_39032_, _00076_, _41654_);
  and (_00077_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_00078_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_00079_, _00078_, _00077_);
  and (_39034_, _00079_, _41654_);
  and (_00080_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_00081_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_00082_, _00081_, _00080_);
  and (_39035_, _00082_, _41654_);
  and (_00083_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_00084_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_00085_, _00084_, _00083_);
  and (_39036_, _00085_, _41654_);
  and (_00086_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_00087_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_00088_, _00087_, _00086_);
  and (_39037_, _00088_, _41654_);
  and (_00089_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_00090_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_00091_, _00090_, _00089_);
  and (_39038_, _00091_, _41654_);
  and (_00092_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_00093_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_00094_, _00093_, _00092_);
  and (_39039_, _00094_, _41654_);
  and (_00095_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_00096_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_00097_, _00096_, _00095_);
  and (_39040_, _00097_, _41654_);
  and (_00098_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_00099_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_00100_, _00099_, _00098_);
  and (_39041_, _00100_, _41654_);
  and (_00101_, _43787_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_00102_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_00103_, _00102_, _00101_);
  and (_39042_, _00103_, _41654_);
  nor (_39044_, _40347_, rst);
  nor (_39045_, _40519_, rst);
  nor (_39046_, _40267_, rst);
  nor (_39047_, _40311_, rst);
  and (_39048_, _40436_, _41654_);
  nor (_39050_, _40228_, rst);
  nor (_39051_, _40372_, rst);
  and (_39067_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _41654_);
  and (_39068_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _41654_);
  and (_39069_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _41654_);
  and (_39071_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _41654_);
  and (_39072_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _41654_);
  and (_39073_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _41654_);
  and (_39074_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _41654_);
  nor (_00104_, _43083_, _43036_);
  nor (_00105_, _00104_, _29615_);
  and (_00106_, _38138_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00107_, _43049_, _40333_);
  and (_00108_, _43044_, _43222_);
  or (_00109_, _00108_, _00107_);
  or (_00110_, _00109_, _00106_);
  nor (_00111_, _43232_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00112_, _00111_, _43241_);
  and (_00113_, _00112_, _43408_);
  nor (_00114_, _00113_, _00110_);
  nand (_00115_, _00114_, _43031_);
  or (_00116_, _00115_, _00105_);
  or (_00117_, _43031_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00118_, _00117_, _41654_);
  and (_39075_, _00118_, _00116_);
  nor (_00119_, _00104_, _30294_);
  and (_00120_, _43049_, _40488_);
  and (_00121_, _43044_, _43193_);
  and (_00122_, _37235_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00123_, _00122_, _00121_);
  or (_00124_, _00123_, _00120_);
  or (_00125_, _43250_, _43241_);
  not (_00126_, _43408_);
  nor (_00127_, _00126_, _43261_);
  and (_00128_, _00127_, _00125_);
  nor (_00129_, _00128_, _00124_);
  nand (_00130_, _00129_, _43031_);
  or (_00131_, _00130_, _00119_);
  or (_00132_, _43031_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00133_, _00132_, _41654_);
  and (_39076_, _00133_, _00131_);
  nor (_00134_, _00104_, _30993_);
  nand (_00135_, _38138_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_00136_, _43049_, _40252_);
  and (_00137_, _43044_, _43154_);
  nor (_00138_, _00137_, _00136_);
  and (_00139_, _00138_, _00135_);
  or (_00140_, _43286_, _43268_);
  nor (_00141_, _00126_, _43287_);
  nand (_00142_, _00141_, _00140_);
  and (_00143_, _00142_, _00139_);
  nand (_00144_, _00143_, _43031_);
  or (_00145_, _00144_, _00134_);
  not (_00146_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00147_, _43429_, _00146_);
  and (_00148_, _43429_, _00146_);
  nor (_00149_, _00148_, _00147_);
  or (_00150_, _00149_, _43031_);
  and (_00151_, _00150_, _41654_);
  and (_39077_, _00151_, _00145_);
  nor (_00152_, _00104_, _31724_);
  or (_00153_, _43148_, _43135_);
  and (_00154_, _00153_, _43300_);
  not (_00155_, _43405_);
  and (_00156_, _43082_, _00155_);
  or (_00157_, _00153_, _43300_);
  nand (_00158_, _00157_, _00156_);
  or (_00159_, _00158_, _00154_);
  and (_00160_, _43049_, _40296_);
  and (_00161_, _43044_, _43131_);
  and (_00162_, _37235_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_00163_, _00162_, _00161_);
  nor (_00164_, _00163_, _00160_);
  and (_00165_, _00164_, _00159_);
  nand (_00166_, _00165_, _43031_);
  or (_00167_, _00166_, _00152_);
  and (_00168_, _00147_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00169_, _00147_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00170_, _00169_, _00168_);
  or (_00171_, _00170_, _43031_);
  and (_00172_, _00171_, _41654_);
  and (_39078_, _00172_, _00167_);
  nor (_00173_, _00104_, _32486_);
  and (_00174_, _43049_, _40424_);
  and (_00175_, _43044_, _43124_);
  and (_00176_, _37235_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00177_, _00176_, _00175_);
  or (_00178_, _00177_, _00174_);
  or (_00179_, _43325_, _43306_);
  and (_00180_, _00156_, _43326_);
  and (_00181_, _00180_, _00179_);
  nor (_00182_, _00181_, _00178_);
  nand (_00183_, _00182_, _43031_);
  or (_00184_, _00183_, _00173_);
  and (_00185_, _43414_, _43430_);
  nor (_00186_, _00168_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00187_, _00186_, _00185_);
  or (_00188_, _00187_, _43031_);
  and (_00189_, _00188_, _41654_);
  and (_39079_, _00189_, _00184_);
  nor (_00190_, _00104_, _33314_);
  and (_00191_, _43049_, _40207_);
  and (_00192_, _43044_, _43117_);
  and (_00193_, _37235_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00194_, _00193_, _00192_);
  or (_00195_, _00194_, _00191_);
  or (_00196_, _43122_, _43120_);
  or (_00197_, _00196_, _43338_);
  nand (_00198_, _00196_, _43338_);
  and (_00199_, _00198_, _00156_);
  and (_00200_, _00199_, _00197_);
  nor (_00201_, _00200_, _00195_);
  nand (_00202_, _00201_, _43031_);
  or (_00203_, _00202_, _00190_);
  and (_00204_, _43416_, _43430_);
  nor (_00205_, _00185_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00206_, _00205_, _00204_);
  or (_00207_, _00206_, _43031_);
  and (_00208_, _00207_, _41654_);
  and (_39080_, _00208_, _00203_);
  nor (_00209_, _00104_, _34032_);
  and (_00210_, _43049_, _40389_);
  and (_00211_, _43044_, _43108_);
  and (_00212_, _37235_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00213_, _00212_, _00211_);
  or (_00214_, _00213_, _00210_);
  or (_00215_, _43346_, _43115_);
  nor (_00216_, _00126_, _43357_);
  and (_00217_, _00216_, _00215_);
  nor (_00218_, _00217_, _00214_);
  nand (_00219_, _00218_, _43031_);
  or (_00220_, _00219_, _00209_);
  and (_00221_, _00204_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00222_, _00204_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00223_, _00222_, _00221_);
  or (_00224_, _00223_, _43031_);
  and (_00225_, _00224_, _41654_);
  and (_39082_, _00225_, _00220_);
  or (_00226_, _43104_, _43105_);
  nor (_00227_, _00226_, _43358_);
  and (_00228_, _00226_, _43358_);
  or (_00229_, _00228_, _00227_);
  or (_00230_, _00229_, _00126_);
  or (_00231_, _00104_, _28465_);
  nand (_00232_, _38138_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nand (_00233_, _43049_, _40138_);
  nand (_00234_, _43044_, _43100_);
  and (_00235_, _00234_, _00233_);
  and (_00236_, _00235_, _00232_);
  and (_00237_, _00236_, _00231_);
  and (_00238_, _00237_, _00230_);
  nand (_00239_, _00238_, _43031_);
  and (_00240_, _00221_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00241_, _00221_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00242_, _00241_, _00240_);
  or (_00243_, _00242_, _43031_);
  and (_00244_, _00243_, _41654_);
  and (_39083_, _00244_, _00239_);
  not (_00245_, _43031_);
  nor (_00246_, _38149_, _29615_);
  and (_00247_, _43374_, _38407_);
  nor (_00248_, _43374_, _38407_);
  nor (_00249_, _00248_, _00247_);
  or (_00250_, _00249_, _43382_);
  nand (_00251_, _00249_, _43382_);
  and (_00252_, _00251_, _43408_);
  and (_00253_, _00252_, _00250_);
  nor (_00254_, _43037_, _38480_);
  and (_00255_, _43049_, _42270_);
  and (_00256_, _43083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_00257_, _43044_, _40333_);
  or (_00258_, _00257_, _00256_);
  or (_00259_, _00258_, _00255_);
  or (_00260_, _00259_, _00254_);
  or (_00261_, _00260_, _00253_);
  or (_00262_, _00261_, _00246_);
  or (_00263_, _00262_, _00245_);
  and (_00264_, _00240_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00265_, _00240_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00266_, _00265_, _00264_);
  or (_00267_, _00266_, _43031_);
  and (_00268_, _00267_, _41654_);
  and (_39084_, _00268_, _00263_);
  and (_00269_, _43374_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00270_, _00269_, _43382_);
  and (_00271_, _43384_, _43103_);
  nor (_00272_, _00271_, _00270_);
  nand (_00273_, _00272_, _38413_);
  or (_00274_, _00272_, _38413_);
  and (_00275_, _00274_, _00156_);
  and (_00276_, _00275_, _00273_);
  nor (_00277_, _43037_, _38509_);
  and (_00278_, _43049_, _42240_);
  and (_00279_, _43083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_00280_, _43044_, _40488_);
  or (_00281_, _00280_, _00279_);
  or (_00282_, _00281_, _00278_);
  nor (_00283_, _00282_, _00277_);
  nand (_00284_, _00283_, _43031_);
  or (_00285_, _00284_, _00276_);
  nor (_00286_, _38149_, _30294_);
  or (_00287_, _00286_, _00285_);
  and (_00288_, _43421_, _43430_);
  nor (_00289_, _00264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00290_, _00289_, _00288_);
  or (_00291_, _00290_, _43031_);
  and (_00292_, _00291_, _41654_);
  and (_39085_, _00292_, _00287_);
  or (_00293_, _38149_, _30993_);
  or (_00294_, _43037_, _38537_);
  nand (_00295_, _43049_, _42277_);
  nand (_00296_, _43083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nand (_00297_, _43044_, _40252_);
  and (_00298_, _00297_, _00296_);
  and (_00299_, _00298_, _00295_);
  and (_00300_, _00299_, _00294_);
  and (_00301_, _43385_, _43103_);
  and (_00302_, _00270_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_00303_, _00302_, _00301_);
  and (_00304_, _00303_, _38418_);
  nor (_00305_, _00303_, _38418_);
  or (_00306_, _00305_, _00304_);
  or (_00307_, _00306_, _00126_);
  and (_00308_, _00307_, _00300_);
  and (_00309_, _00308_, _00293_);
  nand (_00310_, _00309_, _43031_);
  and (_00311_, _00288_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00312_, _00288_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00313_, _00312_, _00311_);
  or (_00314_, _00313_, _43031_);
  and (_00315_, _00314_, _41654_);
  and (_39086_, _00315_, _00310_);
  or (_00316_, _38149_, _31724_);
  or (_00317_, _43037_, _38565_);
  nor (_00318_, _43060_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00319_, _00318_, _43062_);
  nand (_00320_, _00319_, _43049_);
  nand (_00321_, _43083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand (_00322_, _43044_, _40296_);
  and (_00323_, _00322_, _00321_);
  and (_00324_, _00323_, _00320_);
  and (_00325_, _00324_, _00317_);
  and (_00326_, _43376_, _43382_);
  and (_00327_, _43386_, _43103_);
  nor (_00328_, _00327_, _00326_);
  and (_00329_, _00328_, _38403_);
  nor (_00330_, _00328_, _38403_);
  or (_00331_, _00330_, _00126_);
  or (_00332_, _00331_, _00329_);
  and (_00333_, _00332_, _00325_);
  and (_00334_, _00333_, _00316_);
  nand (_00335_, _00334_, _43031_);
  and (_00336_, _00311_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00337_, _00311_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00338_, _00337_, _00336_);
  or (_00339_, _00338_, _43031_);
  and (_00340_, _00339_, _41654_);
  and (_39087_, _00340_, _00335_);
  and (_00341_, _37235_, _32497_);
  and (_00342_, _43377_, _43382_);
  and (_00343_, _43388_, _43103_);
  nor (_00344_, _00343_, _00342_);
  nor (_00345_, _00344_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00346_, _00344_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_00347_, _00346_, _00345_);
  and (_00348_, _00347_, _00156_);
  nor (_00349_, _43037_, _38594_);
  nor (_00350_, _43062_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00351_, _00350_, _43063_);
  and (_00352_, _00351_, _43049_);
  and (_00353_, _43083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_00354_, _43044_, _40424_);
  or (_00355_, _00354_, _00353_);
  or (_00356_, _00355_, _00352_);
  nor (_00357_, _00356_, _00349_);
  nand (_00358_, _00357_, _43031_);
  or (_00359_, _00358_, _00348_);
  or (_00360_, _00359_, _00341_);
  and (_00361_, _00336_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00362_, _00336_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00363_, _00362_, _00361_);
  or (_00364_, _00363_, _43031_);
  and (_00365_, _00364_, _41654_);
  and (_39088_, _00365_, _00360_);
  and (_00366_, _43378_, _43382_);
  and (_00367_, _00343_, _38424_);
  nor (_00368_, _00367_, _00366_);
  nand (_00369_, _00368_, _38399_);
  or (_00370_, _00368_, _38399_);
  and (_00371_, _00370_, _00156_);
  and (_00372_, _00371_, _00369_);
  and (_00373_, _37235_, _33325_);
  nor (_00374_, _43037_, _38626_);
  nor (_00375_, _43063_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00376_, _00375_, _43064_);
  and (_00377_, _00376_, _43049_);
  and (_00378_, _43083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_00379_, _43044_, _40207_);
  or (_00380_, _00379_, _00378_);
  or (_00381_, _00380_, _00377_);
  nor (_00382_, _00381_, _00374_);
  nand (_00383_, _00382_, _43031_);
  or (_00384_, _00383_, _00373_);
  or (_00385_, _00384_, _00372_);
  or (_00386_, _00361_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_00387_, _00361_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_00388_, _00387_, _00386_);
  or (_00389_, _00388_, _43031_);
  and (_00390_, _00389_, _41654_);
  and (_39089_, _00390_, _00385_);
  or (_00391_, _43393_, _38430_);
  nand (_00392_, _43393_, _38430_);
  nand (_00393_, _00392_, _00391_);
  and (_00394_, _00393_, _00156_);
  and (_00395_, _37235_, _34043_);
  or (_00396_, _43037_, _38675_);
  or (_00397_, _43064_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00398_, _00397_, _43066_);
  nand (_00399_, _00398_, _43049_);
  nand (_00400_, _43083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_00401_, _43044_, _40389_);
  and (_00402_, _00401_, _00400_);
  and (_00403_, _00402_, _00399_);
  and (_00404_, _00403_, _00396_);
  nand (_00405_, _00404_, _43031_);
  or (_00406_, _00405_, _00395_);
  or (_00407_, _00406_, _00394_);
  or (_00408_, _43433_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00409_, _00408_, _43435_);
  or (_00410_, _00409_, _43031_);
  and (_00411_, _00410_, _41654_);
  and (_39090_, _00411_, _00407_);
  and (_00412_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_00413_, _43687_, _43684_);
  nor (_00414_, _00413_, _43688_);
  or (_00415_, _00414_, _43447_);
  or (_00416_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00417_, _00416_, _43720_);
  and (_00418_, _00417_, _00415_);
  or (_39091_, _00418_, _00412_);
  nor (_00419_, _43691_, _43688_);
  nor (_00420_, _00419_, _43692_);
  or (_00421_, _00420_, _43447_);
  or (_00422_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00423_, _00422_, _43720_);
  and (_00424_, _00423_, _00421_);
  and (_00425_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39093_, _00425_, _00424_);
  and (_00426_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00427_, _43696_, _43694_);
  nor (_00428_, _00427_, _43697_);
  or (_00429_, _00428_, _43447_);
  or (_00430_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00431_, _00430_, _43720_);
  and (_00432_, _00431_, _00429_);
  or (_39094_, _00432_, _00426_);
  and (_00433_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00434_, _43697_, _43539_);
  nor (_00435_, _00434_, _43698_);
  or (_00436_, _00435_, _43447_);
  or (_00437_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00438_, _00437_, _43720_);
  and (_00439_, _00438_, _00436_);
  or (_39095_, _00439_, _00433_);
  and (_00440_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00441_, _43701_, _43698_);
  nor (_00442_, _00441_, _43702_);
  or (_00443_, _00442_, _43447_);
  or (_00444_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00445_, _00444_, _43720_);
  and (_00446_, _00445_, _00443_);
  or (_39096_, _00446_, _00440_);
  or (_00447_, _43702_, _43533_);
  nor (_00448_, _43703_, _43447_);
  and (_00449_, _00448_, _00447_);
  nor (_00450_, _43446_, _43838_);
  or (_00451_, _00450_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00452_, _00451_, _00449_);
  or (_00453_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _34260_);
  and (_00454_, _00453_, _41654_);
  and (_39097_, _00454_, _00452_);
  nor (_00455_, _43703_, _43527_);
  nor (_00456_, _00455_, _43704_);
  or (_00457_, _00456_, _43447_);
  or (_00458_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00459_, _00458_, _43720_);
  and (_00460_, _00459_, _00457_);
  and (_00461_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39098_, _00461_, _00460_);
  and (_00462_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00463_, _43704_, _43523_);
  nor (_00464_, _00463_, _43705_);
  or (_00465_, _00464_, _43447_);
  or (_00466_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_00467_, _00466_, _43720_);
  and (_00468_, _00467_, _00465_);
  or (_39099_, _00468_, _00462_);
  nor (_00469_, _43707_, _43705_);
  nor (_00470_, _00469_, _43708_);
  or (_00471_, _00470_, _43447_);
  or (_00472_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00473_, _00472_, _43720_);
  and (_00474_, _00473_, _00471_);
  and (_00475_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_39100_, _00475_, _00474_);
  nor (_00476_, _43708_, _43518_);
  nor (_00477_, _00476_, _43709_);
  or (_00478_, _00477_, _43447_);
  or (_00479_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00480_, _00479_, _43720_);
  and (_00481_, _00480_, _00478_);
  and (_00482_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39101_, _00482_, _00481_);
  and (_00483_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00484_, _43709_, _43514_);
  nor (_00485_, _00484_, _43710_);
  or (_00486_, _00485_, _43447_);
  or (_00487_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00488_, _00487_, _43720_);
  and (_00489_, _00488_, _00486_);
  or (_39102_, _00489_, _00483_);
  nor (_00490_, _43710_, _43510_);
  nor (_00491_, _00490_, _43711_);
  or (_00492_, _00491_, _43447_);
  or (_00493_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00494_, _00493_, _43720_);
  and (_00495_, _00494_, _00492_);
  and (_00496_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39104_, _00496_, _00495_);
  nor (_00497_, _43711_, _43507_);
  nor (_00498_, _00497_, _43712_);
  or (_00499_, _00498_, _43447_);
  or (_00500_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00501_, _00500_, _43720_);
  and (_00502_, _00501_, _00499_);
  and (_00503_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_39105_, _00503_, _00502_);
  nor (_00504_, _43712_, _43503_);
  nor (_00505_, _00504_, _43713_);
  or (_00506_, _00505_, _43447_);
  or (_00507_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00508_, _00507_, _43720_);
  and (_00509_, _00508_, _00506_);
  and (_00510_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_39106_, _00510_, _00509_);
  and (_00511_, _43442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_00512_, _43713_, _43501_);
  nor (_00513_, _00512_, _43714_);
  or (_00514_, _00513_, _43447_);
  or (_00515_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00516_, _00515_, _43720_);
  and (_00517_, _00516_, _00514_);
  or (_39107_, _00517_, _00511_);
  and (_00518_, _43730_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_00519_, _00518_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39108_, _00519_, _41654_);
  and (_00520_, _43730_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_00521_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39109_, _00521_, _41654_);
  and (_00522_, _43730_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_00523_, _00522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39110_, _00523_, _41654_);
  and (_00524_, _43730_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_00525_, _00524_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39111_, _00525_, _41654_);
  and (_00526_, _43730_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_00527_, _00526_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39112_, _00527_, _41654_);
  and (_00528_, _43730_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_00529_, _00528_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39113_, _00529_, _41654_);
  and (_00530_, _43730_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_00531_, _00530_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39115_, _00531_, _41654_);
  nor (_00532_, _43683_, _40121_);
  nand (_00533_, _00532_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00534_, _00532_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00535_, _00534_, _43720_);
  and (_39116_, _00535_, _00533_);
  nor (_00536_, _43741_, _43739_);
  nor (_00537_, _00536_, _43742_);
  or (_00538_, _00537_, _40121_);
  or (_00539_, _34293_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00540_, _00539_, _43720_);
  and (_39117_, _00540_, _00538_);
  and (_00541_, _43765_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_00542_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_00543_, _00542_, _38743_);
  or (_39133_, _00543_, _00541_);
  and (_00544_, _43765_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00545_, _00013_, _38743_);
  or (_39134_, _00545_, _00544_);
  and (_00546_, _43765_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00547_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00548_, _00547_, _38743_);
  or (_39135_, _00548_, _00546_);
  and (_00549_, _43765_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00550_, _00020_, _38743_);
  or (_39137_, _00550_, _00549_);
  and (_00551_, _43765_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00552_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_00553_, _00552_, _38743_);
  or (_39138_, _00553_, _00551_);
  and (_00554_, _43765_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00555_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_00556_, _00555_, _38743_);
  or (_39139_, _00556_, _00554_);
  and (_00557_, _43765_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00558_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_00559_, _00558_, _38743_);
  or (_39140_, _00559_, _00557_);
  and (_39141_, _43773_, _41654_);
  nor (_39142_, _43783_, rst);
  and (_39143_, _43779_, _41654_);
  and (_00560_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00561_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00562_, _00561_, _00560_);
  and (_39144_, _00562_, _41654_);
  and (_00563_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00564_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00565_, _00564_, _00563_);
  and (_39145_, _00565_, _41654_);
  and (_00566_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00567_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00568_, _00567_, _00566_);
  and (_39146_, _00568_, _41654_);
  and (_00569_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00570_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00571_, _00570_, _00569_);
  and (_39148_, _00571_, _41654_);
  and (_00572_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00573_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00574_, _00573_, _00572_);
  and (_39149_, _00574_, _41654_);
  and (_00575_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00576_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00577_, _00576_, _00575_);
  and (_39150_, _00577_, _41654_);
  and (_00578_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00579_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00580_, _00579_, _00578_);
  and (_39151_, _00580_, _41654_);
  and (_00581_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00582_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00583_, _00582_, _00581_);
  and (_39152_, _00583_, _41654_);
  and (_00584_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00585_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00586_, _00585_, _00584_);
  and (_39153_, _00586_, _41654_);
  and (_00587_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00588_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00589_, _00588_, _00587_);
  and (_39154_, _00589_, _41654_);
  and (_00590_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00591_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00592_, _00591_, _00590_);
  and (_39155_, _00592_, _41654_);
  and (_00593_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00594_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00595_, _00594_, _00593_);
  and (_39156_, _00595_, _41654_);
  and (_00596_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00597_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00598_, _00597_, _00596_);
  and (_39157_, _00598_, _41654_);
  and (_00599_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00600_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00601_, _00600_, _00599_);
  and (_39158_, _00601_, _41654_);
  and (_00602_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00603_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00604_, _00603_, _00602_);
  and (_39159_, _00604_, _41654_);
  and (_00605_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00606_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00607_, _00606_, _00605_);
  and (_39160_, _00607_, _41654_);
  and (_00608_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00609_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00610_, _00609_, _00608_);
  and (_39161_, _00610_, _41654_);
  and (_00611_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00612_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00613_, _00612_, _00611_);
  and (_39162_, _00613_, _41654_);
  and (_00614_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00615_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00616_, _00615_, _00614_);
  and (_39163_, _00616_, _41654_);
  and (_00617_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00618_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00619_, _00618_, _00617_);
  and (_39164_, _00619_, _41654_);
  and (_00620_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00621_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00622_, _00621_, _00620_);
  and (_39165_, _00622_, _41654_);
  and (_00623_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00624_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00625_, _00624_, _00623_);
  and (_39166_, _00625_, _41654_);
  and (_00626_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00627_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00628_, _00627_, _00626_);
  and (_39167_, _00628_, _41654_);
  and (_00629_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00630_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00631_, _00630_, _00629_);
  and (_39169_, _00631_, _41654_);
  and (_00632_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00633_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00634_, _00633_, _00632_);
  and (_39170_, _00634_, _41654_);
  and (_00635_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00636_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00637_, _00636_, _00635_);
  and (_39171_, _00637_, _41654_);
  and (_00638_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00639_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00640_, _00639_, _00638_);
  and (_39172_, _00640_, _41654_);
  and (_00641_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00642_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00643_, _00642_, _00641_);
  and (_39173_, _00643_, _41654_);
  and (_00644_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00645_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00646_, _00645_, _00644_);
  and (_39174_, _00646_, _41654_);
  and (_00647_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00648_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00649_, _00648_, _00647_);
  and (_39175_, _00649_, _41654_);
  and (_00650_, _43787_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00651_, _43789_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00652_, _00651_, _00650_);
  and (_39176_, _00652_, _41654_);
  and (_00653_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00654_, _43797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00655_, _00654_, _00653_);
  and (_39177_, _00655_, _41654_);
  and (_00656_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00657_, _43797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00658_, _00657_, _00656_);
  and (_39178_, _00658_, _41654_);
  and (_00659_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00660_, _43797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00661_, _00660_, _00659_);
  and (_39180_, _00661_, _41654_);
  and (_00662_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00663_, _43797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00664_, _00663_, _00662_);
  and (_39181_, _00664_, _41654_);
  and (_00665_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00666_, _43797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00667_, _00666_, _00665_);
  and (_39182_, _00667_, _41654_);
  and (_00668_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00669_, _43797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00670_, _00669_, _00668_);
  and (_39183_, _00670_, _41654_);
  and (_00671_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00672_, _43797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00673_, _00672_, _00671_);
  and (_39184_, _00673_, _41654_);
  and (_00674_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00675_, _40347_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00676_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00677_, _00676_, _43796_);
  and (_00678_, _00677_, _00675_);
  or (_00679_, _00678_, _00674_);
  and (_39185_, _00679_, _41654_);
  and (_00680_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00681_, _40519_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00682_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00683_, _00682_, _43796_);
  and (_00684_, _00683_, _00681_);
  or (_00685_, _00684_, _00680_);
  and (_39186_, _00685_, _41654_);
  and (_00686_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00687_, _40267_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00688_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00689_, _00688_, _43796_);
  and (_00690_, _00689_, _00687_);
  or (_00691_, _00690_, _00686_);
  and (_39187_, _00691_, _41654_);
  and (_00692_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00693_, _40311_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00694_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00695_, _00694_, _43796_);
  and (_00696_, _00695_, _00693_);
  or (_00697_, _00696_, _00692_);
  and (_39188_, _00697_, _41654_);
  and (_00698_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00699_, _40436_, _43803_);
  or (_00700_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00701_, _00700_, _43796_);
  and (_00702_, _00701_, _00699_);
  or (_00703_, _00702_, _00698_);
  and (_39189_, _00703_, _41654_);
  and (_00704_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00705_, _40228_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00706_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00707_, _00706_, _43796_);
  and (_00708_, _00707_, _00705_);
  or (_00709_, _00708_, _00704_);
  and (_39191_, _00709_, _41654_);
  and (_00710_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00711_, _40372_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00712_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00713_, _00712_, _43796_);
  and (_00714_, _00713_, _00711_);
  or (_00715_, _00714_, _00710_);
  and (_39192_, _00715_, _41654_);
  and (_00716_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00717_, _40171_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00718_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00719_, _00718_, _43796_);
  and (_00720_, _00719_, _00717_);
  or (_00721_, _00720_, _00716_);
  and (_39193_, _00721_, _41654_);
  and (_00722_, _43803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00723_, _00722_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00724_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _43796_);
  and (_00725_, _00724_, _41654_);
  and (_39194_, _00725_, _00723_);
  and (_00726_, _43803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00727_, _00726_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00728_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _43796_);
  and (_00729_, _00728_, _41654_);
  and (_39195_, _00729_, _00727_);
  and (_00730_, _43803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00731_, _00730_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00732_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _43796_);
  and (_00733_, _00732_, _41654_);
  and (_39196_, _00733_, _00731_);
  and (_00734_, _43803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00735_, _00734_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00736_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _43796_);
  and (_00737_, _00736_, _41654_);
  and (_39197_, _00737_, _00735_);
  and (_00738_, _43803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00739_, _00738_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00740_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _43796_);
  and (_00741_, _00740_, _41654_);
  and (_39198_, _00741_, _00739_);
  and (_00742_, _43803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_00743_, _00742_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00744_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _43796_);
  and (_00745_, _00744_, _41654_);
  and (_39199_, _00745_, _00743_);
  and (_00746_, _43803_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_00747_, _00746_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00748_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _43796_);
  and (_00749_, _00748_, _41654_);
  and (_39200_, _00749_, _00747_);
  nand (_00750_, _43810_, _29615_);
  or (_00751_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00752_, _00751_, _41654_);
  and (_39202_, _00752_, _00750_);
  nand (_00753_, _43810_, _30294_);
  or (_00754_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00755_, _00754_, _41654_);
  and (_39203_, _00755_, _00753_);
  nand (_00756_, _43810_, _30993_);
  or (_00757_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00758_, _00757_, _41654_);
  and (_39204_, _00758_, _00756_);
  nand (_00759_, _43810_, _31724_);
  or (_00760_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00761_, _00760_, _41654_);
  and (_39205_, _00761_, _00759_);
  nand (_00762_, _43810_, _32486_);
  or (_00763_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00764_, _00763_, _41654_);
  and (_39206_, _00764_, _00762_);
  nand (_00765_, _43810_, _33314_);
  or (_00766_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00767_, _00766_, _41654_);
  and (_39207_, _00767_, _00765_);
  nand (_00768_, _43810_, _34032_);
  or (_00769_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00770_, _00769_, _41654_);
  and (_39208_, _00770_, _00768_);
  nand (_00771_, _43810_, _28465_);
  or (_00772_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00773_, _00772_, _41654_);
  and (_39209_, _00773_, _00771_);
  nand (_00774_, _43810_, _38480_);
  or (_00775_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00776_, _00775_, _41654_);
  and (_39210_, _00776_, _00774_);
  nand (_00777_, _43810_, _38509_);
  or (_00778_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00779_, _00778_, _41654_);
  and (_39211_, _00779_, _00777_);
  nand (_00780_, _43810_, _38537_);
  or (_00781_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00782_, _00781_, _41654_);
  and (_39213_, _00782_, _00780_);
  nand (_00783_, _43810_, _38565_);
  or (_00784_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00785_, _00784_, _41654_);
  and (_39214_, _00785_, _00783_);
  nand (_00786_, _43810_, _38594_);
  or (_00787_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00788_, _00787_, _41654_);
  and (_39215_, _00788_, _00786_);
  nand (_00789_, _43810_, _38626_);
  or (_00790_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00791_, _00790_, _41654_);
  and (_39216_, _00791_, _00789_);
  nand (_00792_, _43810_, _38675_);
  or (_00793_, _43810_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00794_, _00793_, _41654_);
  and (_39217_, _00794_, _00792_);
  nor (_39429_, _40189_, rst);
  and (_00795_, _38993_, _25395_);
  and (_00796_, _00795_, _40146_);
  nand (_00797_, _00796_, _38307_);
  or (_00798_, _00796_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_00799_, _00798_, _41654_);
  and (_39430_, _00799_, _00797_);
  and (_00800_, _38218_, _25395_);
  not (_00801_, _00800_);
  nor (_00802_, _00801_, _38307_);
  not (_00803_, _40146_);
  and (_00804_, _00801_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_00805_, _00804_, _00803_);
  or (_00806_, _00805_, _00802_);
  or (_00807_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_00808_, _00807_, _41654_);
  and (_39431_, _00808_, _00806_);
  and (_00809_, _39725_, _24895_);
  and (_00810_, _00809_, _25395_);
  not (_00811_, _00810_);
  nor (_00812_, _00811_, _38307_);
  and (_00813_, _00811_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_00814_, _00813_, _00803_);
  or (_00815_, _00814_, _00812_);
  or (_00816_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_00817_, _00816_, _41654_);
  and (_39433_, _00817_, _00815_);
  and (_00818_, _39725_, _30414_);
  and (_00819_, _00818_, _25395_);
  not (_00820_, _00819_);
  nor (_00821_, _00820_, _38307_);
  and (_00822_, _00820_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_00823_, _00822_, _00803_);
  or (_00824_, _00823_, _00821_);
  or (_00825_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_00826_, _00825_, _41654_);
  and (_39434_, _00826_, _00824_);
  nand (_00827_, _00796_, _38285_);
  or (_00828_, _00796_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_00829_, _00828_, _41654_);
  and (_39462_, _00829_, _00827_);
  nand (_00830_, _00796_, _38276_);
  or (_00831_, _00796_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_00832_, _00831_, _41654_);
  and (_39463_, _00832_, _00830_);
  nand (_00833_, _00796_, _38269_);
  or (_00834_, _00796_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_00835_, _00834_, _41654_);
  and (_39464_, _00835_, _00833_);
  nand (_00836_, _00796_, _38261_);
  or (_00837_, _00796_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_00838_, _00837_, _41654_);
  and (_39465_, _00838_, _00836_);
  nand (_00839_, _00796_, _38253_);
  or (_00841_, _00796_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_00842_, _00841_, _41654_);
  and (_39466_, _00842_, _00839_);
  nand (_00843_, _00796_, _38246_);
  or (_00844_, _00796_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_00845_, _00844_, _41654_);
  and (_39467_, _00845_, _00843_);
  nand (_00846_, _00796_, _38239_);
  or (_00847_, _00796_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_00848_, _00847_, _41654_);
  and (_39468_, _00848_, _00846_);
  nor (_00849_, _00801_, _38285_);
  and (_00850_, _00801_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_00851_, _00850_, _00803_);
  or (_00852_, _00851_, _00849_);
  or (_00853_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_00854_, _00853_, _41654_);
  and (_39469_, _00854_, _00852_);
  nor (_00855_, _00801_, _38276_);
  and (_00856_, _00801_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_00857_, _00856_, _00803_);
  or (_00858_, _00857_, _00855_);
  or (_00859_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_00860_, _00859_, _41654_);
  and (_39470_, _00860_, _00858_);
  nor (_00861_, _00801_, _38269_);
  and (_00862_, _00801_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_00863_, _00862_, _00803_);
  or (_00864_, _00863_, _00861_);
  or (_00865_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_00867_, _00865_, _41654_);
  and (_39471_, _00867_, _00864_);
  nor (_00868_, _00801_, _38261_);
  and (_00869_, _00801_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_00870_, _00869_, _00803_);
  or (_00871_, _00870_, _00868_);
  or (_00872_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_00873_, _00872_, _41654_);
  and (_39472_, _00873_, _00871_);
  nor (_00874_, _00801_, _38253_);
  and (_00875_, _00801_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_00876_, _00875_, _00803_);
  or (_00877_, _00876_, _00874_);
  or (_00878_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_00879_, _00878_, _41654_);
  and (_39473_, _00879_, _00877_);
  nor (_00880_, _00801_, _38246_);
  and (_00881_, _00801_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_00882_, _00881_, _00803_);
  or (_00883_, _00882_, _00880_);
  or (_00885_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_00886_, _00885_, _41654_);
  and (_39474_, _00886_, _00883_);
  nor (_00887_, _00801_, _38239_);
  and (_00888_, _00801_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_00889_, _00888_, _00803_);
  or (_00890_, _00889_, _00887_);
  or (_00891_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_00892_, _00891_, _41654_);
  and (_39475_, _00892_, _00890_);
  or (_00893_, _00810_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand (_00894_, _00810_, _38285_);
  and (_00895_, _00894_, _00893_);
  or (_00896_, _00895_, _00803_);
  or (_00897_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_00898_, _00897_, _41654_);
  and (_39476_, _00898_, _00896_);
  nor (_00899_, _00811_, _38276_);
  and (_00900_, _00811_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_00901_, _00900_, _00803_);
  or (_00902_, _00901_, _00899_);
  or (_00903_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_00904_, _00903_, _41654_);
  and (_39478_, _00904_, _00902_);
  and (_00905_, _00810_, _40146_);
  nand (_00906_, _00905_, _38269_);
  or (_00907_, _00905_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_00908_, _00907_, _41654_);
  and (_39479_, _00908_, _00906_);
  nor (_00909_, _00811_, _38261_);
  and (_00910_, _00811_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_00911_, _00910_, _00803_);
  or (_00912_, _00911_, _00909_);
  or (_00913_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_00914_, _00913_, _41654_);
  and (_39480_, _00914_, _00912_);
  nor (_00915_, _00811_, _38253_);
  and (_00916_, _00811_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_00917_, _00916_, _00803_);
  or (_00918_, _00917_, _00915_);
  or (_00919_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_00920_, _00919_, _41654_);
  and (_39481_, _00920_, _00918_);
  nor (_00921_, _00811_, _38246_);
  and (_00922_, _00811_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_00923_, _00922_, _00803_);
  or (_00924_, _00923_, _00921_);
  or (_00925_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_00926_, _00925_, _41654_);
  and (_39482_, _00926_, _00924_);
  nor (_00927_, _00811_, _38239_);
  and (_00928_, _00811_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_00929_, _00928_, _00803_);
  or (_00930_, _00929_, _00927_);
  or (_00931_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_00932_, _00931_, _41654_);
  and (_39483_, _00932_, _00930_);
  and (_00933_, _00820_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_00934_, _00820_, _38285_);
  or (_00935_, _00934_, _00803_);
  or (_00936_, _00935_, _00933_);
  or (_00937_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_00938_, _00937_, _41654_);
  and (_39484_, _00938_, _00936_);
  nor (_00939_, _00820_, _38276_);
  and (_00940_, _00820_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_00941_, _00940_, _00803_);
  or (_00942_, _00941_, _00939_);
  or (_00943_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_00944_, _00943_, _41654_);
  and (_39485_, _00944_, _00942_);
  nor (_00945_, _00820_, _38269_);
  and (_00946_, _00820_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_00947_, _00946_, _00803_);
  or (_00948_, _00947_, _00945_);
  or (_00949_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_00950_, _00949_, _41654_);
  and (_39486_, _00950_, _00948_);
  nor (_00951_, _00820_, _38261_);
  and (_00952_, _00820_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_00953_, _00952_, _00803_);
  or (_00954_, _00953_, _00951_);
  or (_00955_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_00956_, _00955_, _41654_);
  and (_39487_, _00956_, _00954_);
  nor (_00957_, _00820_, _38253_);
  and (_00958_, _00820_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_00959_, _00958_, _00803_);
  or (_00960_, _00959_, _00957_);
  or (_00961_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_00962_, _00961_, _41654_);
  and (_39489_, _00962_, _00960_);
  nor (_00963_, _00820_, _38246_);
  and (_00964_, _00820_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_00965_, _00964_, _00803_);
  or (_00966_, _00965_, _00963_);
  or (_00967_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_00968_, _00967_, _41654_);
  and (_39490_, _00968_, _00966_);
  nor (_00969_, _00820_, _38239_);
  and (_00970_, _00820_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_00971_, _00970_, _00803_);
  or (_00972_, _00971_, _00969_);
  or (_00973_, _40146_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_00974_, _00973_, _41654_);
  and (_39491_, _00974_, _00972_);
  and (_00975_, _40315_, _40466_);
  and (_00976_, _00975_, _40232_);
  nor (_00977_, _40396_, _40176_);
  and (_00978_, _00977_, _00976_);
  not (_00979_, _40271_);
  nor (_00980_, _38954_, _38938_);
  and (_00981_, _38954_, _38938_);
  nor (_00982_, _00981_, _00980_);
  and (_00983_, _38927_, _38915_);
  nor (_00984_, _38927_, _38915_);
  or (_00985_, _00984_, _00983_);
  nor (_00986_, _00985_, _00982_);
  and (_00987_, _00985_, _00982_);
  nor (_00988_, _00987_, _00986_);
  nor (_00989_, _38976_, _38965_);
  and (_00990_, _38976_, _38965_);
  nor (_00991_, _00990_, _00989_);
  not (_00992_, _38904_);
  nor (_00993_, _38987_, _00992_);
  and (_00994_, _38987_, _00992_);
  nor (_00995_, _00994_, _00993_);
  nor (_00996_, _00995_, _00991_);
  and (_00997_, _00995_, _00991_);
  or (_00998_, _00997_, _00996_);
  or (_00999_, _00998_, _00988_);
  nand (_01000_, _00998_, _00988_);
  and (_01001_, _01000_, _00999_);
  or (_01002_, _01001_, _00979_);
  and (_01003_, _40351_, _40548_);
  or (_01004_, _40271_, _38851_);
  and (_01005_, _01004_, _01003_);
  and (_01006_, _01005_, _01002_);
  nor (_01007_, _40351_, _40548_);
  and (_01008_, _01007_, _40271_);
  and (_01009_, _01008_, _38841_);
  or (_01010_, _40271_, _38858_);
  not (_01011_, _40351_);
  and (_01012_, _01011_, _40548_);
  or (_01013_, _00979_, _38768_);
  and (_01014_, _01013_, _01012_);
  and (_01015_, _01014_, _01010_);
  and (_01016_, _01007_, _00979_);
  and (_01017_, _01016_, _38730_);
  or (_01018_, _01017_, _01015_);
  or (_01019_, _01018_, _01009_);
  or (_01020_, _00979_, _38833_);
  nor (_01021_, _01011_, _40548_);
  or (_01022_, _40271_, _38876_);
  and (_01023_, _01022_, _01021_);
  and (_01024_, _01023_, _01020_);
  or (_01025_, _01024_, _01019_);
  or (_01026_, _01025_, _01006_);
  and (_01027_, _01026_, _00978_);
  and (_01028_, _35223_, _42363_);
  not (_01029_, _01028_);
  nor (_01030_, _42364_, _37491_);
  and (_01031_, _01030_, _01029_);
  nor (_01032_, _37590_, _37535_);
  and (_01033_, _01032_, _01031_);
  not (_01034_, _42433_);
  nor (_01035_, _01034_, _42362_);
  and (_01036_, _01035_, _01033_);
  nor (_01037_, _42431_, _36272_);
  and (_01038_, _37036_, _38160_);
  not (_01039_, _01038_);
  and (_01040_, _01039_, _01037_);
  and (_01041_, _01040_, _42734_);
  and (_01042_, _01041_, _01036_);
  and (_01043_, _01042_, _37876_);
  nor (_01044_, _01043_, _34249_);
  and (_01045_, _42912_, p3in_reg[6]);
  and (_01046_, _42908_, p3_in[6]);
  or (_01047_, _01046_, _01045_);
  or (_01048_, _01047_, _01044_);
  not (_01049_, _01044_);
  or (_01050_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_01051_, _01050_, _01048_);
  and (_01052_, _01051_, _01021_);
  or (_01053_, _01052_, _40271_);
  and (_01054_, _42912_, p3in_reg[7]);
  and (_01055_, _42908_, p3_in[7]);
  or (_01056_, _01055_, _01054_);
  or (_01057_, _01056_, _01044_);
  or (_01058_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_01059_, _01058_, _01057_);
  and (_01060_, _01059_, _01007_);
  and (_01061_, _42912_, p3in_reg[5]);
  and (_01062_, _42908_, p3_in[5]);
  or (_01063_, _01062_, _01061_);
  or (_01064_, _01063_, _01044_);
  or (_01065_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01066_, _01065_, _01064_);
  and (_01067_, _01066_, _01012_);
  and (_01068_, _42912_, p3in_reg[4]);
  and (_01069_, _42908_, p3_in[4]);
  or (_01070_, _01069_, _01068_);
  or (_01071_, _01070_, _01044_);
  or (_01072_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_01073_, _01072_, _01071_);
  and (_01074_, _01073_, _01003_);
  or (_01075_, _01074_, _01067_);
  or (_01076_, _01075_, _01060_);
  or (_01077_, _01076_, _01053_);
  and (_01078_, _40396_, _40233_);
  not (_01079_, _40176_);
  and (_01080_, _00975_, _01079_);
  and (_01081_, _01080_, _01078_);
  and (_01082_, _42912_, p3in_reg[2]);
  and (_01083_, _42908_, p3_in[2]);
  or (_01084_, _01083_, _01082_);
  or (_01085_, _01084_, _01044_);
  or (_01086_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_01087_, _01086_, _01085_);
  and (_01088_, _01087_, _01021_);
  or (_01089_, _01088_, _00979_);
  and (_01090_, _42912_, p3in_reg[3]);
  and (_01091_, _42908_, p3_in[3]);
  or (_01092_, _01091_, _01090_);
  or (_01093_, _01092_, _01044_);
  or (_01094_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_01095_, _01094_, _01093_);
  and (_01096_, _01095_, _01007_);
  and (_01097_, _42912_, p3in_reg[1]);
  and (_01098_, _42908_, p3_in[1]);
  or (_01099_, _01098_, _01097_);
  or (_01100_, _01099_, _01044_);
  or (_01101_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_01102_, _01101_, _01100_);
  and (_01103_, _01102_, _01012_);
  and (_01104_, _42912_, p3in_reg[0]);
  and (_01105_, _42908_, p3_in[0]);
  or (_01106_, _01105_, _01104_);
  or (_01107_, _01106_, _01044_);
  or (_01108_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_01109_, _01108_, _01107_);
  and (_01110_, _01109_, _01003_);
  or (_01111_, _01110_, _01103_);
  or (_01112_, _01111_, _01096_);
  or (_01113_, _01112_, _01089_);
  and (_01114_, _01113_, _01081_);
  and (_01115_, _01114_, _01077_);
  and (_01116_, _42912_, p2in_reg[5]);
  and (_01117_, _42908_, p2_in[5]);
  or (_01118_, _01117_, _01116_);
  or (_01119_, _01118_, _01044_);
  or (_01120_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01121_, _01120_, _01119_);
  and (_01122_, _01121_, _01012_);
  or (_01123_, _01122_, _40271_);
  and (_01124_, _42912_, p2in_reg[7]);
  and (_01125_, _42908_, p2_in[7]);
  or (_01126_, _01125_, _01124_);
  or (_01127_, _01126_, _01044_);
  or (_01128_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_01129_, _01128_, _01127_);
  and (_01130_, _01129_, _01007_);
  and (_01131_, _42912_, p2in_reg[4]);
  and (_01132_, _42908_, p2_in[4]);
  or (_01133_, _01132_, _01131_);
  or (_01134_, _01133_, _01044_);
  or (_01135_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_01136_, _01135_, _01134_);
  and (_01137_, _01136_, _01003_);
  and (_01138_, _42912_, p2in_reg[6]);
  and (_01139_, _42908_, p2_in[6]);
  or (_01140_, _01139_, _01138_);
  or (_01141_, _01140_, _01044_);
  or (_01142_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_01143_, _01142_, _01141_);
  and (_01144_, _01143_, _01021_);
  or (_01145_, _01144_, _01137_);
  or (_01146_, _01145_, _01130_);
  or (_01147_, _01146_, _01123_);
  nor (_01148_, _40466_, _40176_);
  and (_01149_, _01148_, _40315_);
  and (_01150_, _01149_, _01078_);
  and (_01151_, _42912_, p2in_reg[1]);
  and (_01152_, _42908_, p2_in[1]);
  or (_01153_, _01152_, _01151_);
  or (_01154_, _01153_, _01044_);
  or (_01155_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_01156_, _01155_, _01154_);
  and (_01157_, _01156_, _01012_);
  or (_01158_, _01157_, _00979_);
  and (_01159_, _42912_, p2in_reg[3]);
  and (_01160_, _42908_, p2_in[3]);
  or (_01161_, _01160_, _01159_);
  or (_01162_, _01161_, _01044_);
  or (_01163_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_01164_, _01163_, _01162_);
  and (_01165_, _01164_, _01007_);
  and (_01166_, _42912_, p2in_reg[0]);
  and (_01167_, _42908_, p2_in[0]);
  or (_01168_, _01167_, _01166_);
  or (_01169_, _01168_, _01044_);
  or (_01170_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_01171_, _01170_, _01169_);
  and (_01172_, _01171_, _01003_);
  and (_01173_, _42912_, p2in_reg[2]);
  and (_01174_, _42908_, p2_in[2]);
  or (_01175_, _01174_, _01173_);
  or (_01176_, _01175_, _01044_);
  or (_01177_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_01178_, _01177_, _01176_);
  and (_01179_, _01178_, _01021_);
  or (_01180_, _01179_, _01172_);
  or (_01181_, _01180_, _01165_);
  or (_01182_, _01181_, _01158_);
  and (_01183_, _01182_, _01150_);
  and (_01184_, _01183_, _01147_);
  or (_01185_, _01184_, _01115_);
  and (_01186_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_01187_, _01186_, _00979_);
  and (_01188_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_01189_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_01190_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_01191_, _01190_, _01189_);
  or (_01192_, _01191_, _01188_);
  or (_01193_, _01192_, _01187_);
  and (_01194_, _01148_, _40316_);
  and (_01195_, _01194_, _01078_);
  and (_01196_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01197_, _01196_, _40271_);
  and (_01198_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_01199_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_01200_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01201_, _01200_, _01199_);
  or (_01202_, _01201_, _01198_);
  or (_01203_, _01202_, _01197_);
  and (_01204_, _01203_, _01195_);
  and (_01205_, _01204_, _01193_);
  and (_01206_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_01207_, _01206_, _00979_);
  and (_01208_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_01209_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_01210_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_01211_, _01210_, _01209_);
  or (_01212_, _01211_, _01208_);
  or (_01213_, _01212_, _01207_);
  and (_01214_, _40396_, _40232_);
  and (_01215_, _01214_, _01194_);
  and (_01216_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_01217_, _01216_, _40271_);
  and (_01218_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_01219_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_01220_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_01221_, _01220_, _01219_);
  or (_01222_, _01221_, _01218_);
  or (_01223_, _01222_, _01217_);
  and (_01224_, _01223_, _01215_);
  and (_01225_, _01224_, _01213_);
  or (_01226_, _01225_, _01205_);
  and (_01227_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_01228_, _01227_, _00979_);
  and (_01229_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_01230_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01231_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_01232_, _01231_, _01230_);
  or (_01233_, _01232_, _01229_);
  or (_01234_, _01233_, _01228_);
  nor (_01235_, _40396_, _40232_);
  and (_01236_, _01235_, _01080_);
  and (_01237_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_01238_, _01237_, _40271_);
  and (_01239_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_01240_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01241_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_01242_, _01241_, _01240_);
  or (_01243_, _01242_, _01239_);
  or (_01244_, _01243_, _01238_);
  and (_01245_, _01244_, _01236_);
  and (_01246_, _01245_, _01234_);
  and (_01247_, _42912_, p0in_reg[0]);
  and (_01248_, _42908_, p0_in[0]);
  or (_01249_, _01248_, _01247_);
  or (_01250_, _01249_, _01044_);
  nand (_01251_, _01044_, _39248_);
  and (_01252_, _01251_, _01250_);
  and (_01253_, _01252_, _01003_);
  or (_01254_, _01253_, _00979_);
  and (_01255_, _42912_, p0in_reg[3]);
  and (_01256_, _42908_, p0_in[3]);
  or (_01257_, _01256_, _01255_);
  or (_01258_, _01257_, _01044_);
  nand (_01259_, _01044_, _39286_);
  and (_01260_, _01259_, _01258_);
  and (_01261_, _01260_, _01007_);
  and (_01262_, _42912_, p0in_reg[2]);
  and (_01263_, _42908_, p0_in[2]);
  or (_01264_, _01263_, _01262_);
  or (_01265_, _01264_, _01044_);
  or (_01266_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_01267_, _01266_, _01265_);
  and (_01268_, _01267_, _01021_);
  and (_01269_, _42912_, p0in_reg[1]);
  and (_01270_, _42908_, p0_in[1]);
  or (_01271_, _01270_, _01269_);
  or (_01272_, _01271_, _01044_);
  or (_01273_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01274_, _01273_, _01272_);
  and (_01275_, _01274_, _01012_);
  or (_01276_, _01275_, _01268_);
  or (_01277_, _01276_, _01261_);
  or (_01278_, _01277_, _01254_);
  and (_01279_, _01214_, _01149_);
  and (_01280_, _42912_, p0in_reg[4]);
  and (_01281_, _42908_, p0_in[4]);
  or (_01282_, _01281_, _01280_);
  or (_01283_, _01282_, _01044_);
  or (_01284_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01285_, _01284_, _01283_);
  and (_01286_, _01285_, _01003_);
  or (_01287_, _01286_, _40271_);
  and (_01288_, _42912_, p0in_reg[7]);
  and (_01289_, _42908_, p0_in[7]);
  or (_01290_, _01289_, _01288_);
  or (_01291_, _01290_, _01044_);
  or (_01292_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_01293_, _01292_, _01291_);
  and (_01294_, _01293_, _01007_);
  and (_01295_, _42912_, p0in_reg[6]);
  and (_01296_, _42908_, p0_in[6]);
  or (_01297_, _01296_, _01295_);
  or (_01298_, _01297_, _01044_);
  or (_01299_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_01300_, _01299_, _01298_);
  and (_01301_, _01300_, _01021_);
  and (_01302_, _42912_, p0in_reg[5]);
  and (_01303_, _42908_, p0_in[5]);
  or (_01304_, _01303_, _01302_);
  or (_01305_, _01304_, _01044_);
  or (_01306_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01307_, _01306_, _01305_);
  and (_01308_, _01307_, _01012_);
  or (_01309_, _01308_, _01301_);
  or (_01310_, _01309_, _01294_);
  or (_01311_, _01310_, _01287_);
  and (_01312_, _01311_, _01279_);
  and (_01313_, _01312_, _01278_);
  or (_01314_, _01313_, _01246_);
  or (_01315_, _01314_, _01226_);
  or (_01316_, _01315_, _01185_);
  nor (_01317_, _40315_, _40176_);
  and (_01318_, _40396_, _40466_);
  and (_01319_, _01318_, _01317_);
  and (_01320_, _01194_, _40396_);
  or (_01321_, _01320_, _01319_);
  nor (_01322_, _01321_, _01236_);
  and (_01323_, _01235_, _01149_);
  not (_01324_, _01323_);
  nor (_01325_, _40316_, _40176_);
  and (_01326_, _01325_, _40396_);
  nor (_01327_, _01326_, _00978_);
  and (_01328_, _01327_, _01324_);
  and (_01329_, _01328_, _01322_);
  nand (_01330_, _43026_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_01331_, _01330_, _01329_);
  and (_01332_, _42912_, p1in_reg[2]);
  and (_01333_, _42908_, p1_in[2]);
  or (_01334_, _01333_, _01332_);
  or (_01335_, _01334_, _01044_);
  or (_01336_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_01337_, _01336_, _01335_);
  and (_01338_, _01337_, _01021_);
  or (_01339_, _01338_, _00979_);
  and (_01340_, _42912_, p1in_reg[3]);
  and (_01341_, _42908_, p1_in[3]);
  or (_01342_, _01341_, _01340_);
  or (_01343_, _01342_, _01044_);
  or (_01344_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_01345_, _01344_, _01343_);
  and (_01346_, _01345_, _01007_);
  and (_01347_, _42912_, p1in_reg[1]);
  and (_01348_, _42908_, p1_in[1]);
  or (_01349_, _01348_, _01347_);
  or (_01350_, _01349_, _01044_);
  or (_01351_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_01352_, _01351_, _01350_);
  and (_01353_, _01352_, _01012_);
  and (_01354_, _42912_, p1in_reg[0]);
  and (_01355_, _42908_, p1_in[0]);
  or (_01356_, _01355_, _01354_);
  or (_01357_, _01356_, _01044_);
  or (_01358_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_01359_, _01358_, _01357_);
  and (_01360_, _01359_, _01003_);
  or (_01361_, _01360_, _01353_);
  or (_01362_, _01361_, _01346_);
  or (_01363_, _01362_, _01339_);
  and (_01365_, _01214_, _01080_);
  and (_01367_, _42912_, p1in_reg[6]);
  and (_01369_, _42908_, p1_in[6]);
  or (_01371_, _01369_, _01367_);
  or (_01373_, _01371_, _01044_);
  or (_01375_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_01377_, _01375_, _01373_);
  and (_01378_, _01377_, _01021_);
  or (_01379_, _01378_, _40271_);
  and (_01380_, _42912_, p1in_reg[7]);
  and (_01381_, _42908_, p1_in[7]);
  or (_01382_, _01381_, _01380_);
  or (_01383_, _01382_, _01044_);
  or (_01385_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_01386_, _01385_, _01383_);
  and (_01388_, _01386_, _01007_);
  and (_01389_, _42912_, p1in_reg[5]);
  and (_01390_, _42908_, p1_in[5]);
  or (_01392_, _01390_, _01389_);
  or (_01393_, _01392_, _01044_);
  or (_01394_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01396_, _01394_, _01393_);
  and (_01397_, _01396_, _01012_);
  and (_01398_, _42912_, p1in_reg[4]);
  and (_01400_, _42908_, p1_in[4]);
  or (_01401_, _01400_, _01398_);
  or (_01402_, _01401_, _01044_);
  or (_01404_, _01049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01405_, _01404_, _01402_);
  and (_01406_, _01405_, _01003_);
  or (_01408_, _01406_, _01397_);
  or (_01409_, _01408_, _01388_);
  or (_01410_, _01409_, _01379_);
  and (_01412_, _01410_, _01365_);
  and (_01413_, _01412_, _01363_);
  and (_01414_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01416_, _01414_, _00979_);
  and (_01417_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_01418_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_01419_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_01420_, _01419_, _01418_);
  or (_01421_, _01420_, _01417_);
  or (_01422_, _01421_, _01416_);
  and (_01423_, _01319_, _40233_);
  and (_01424_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_01425_, _01424_, _40271_);
  and (_01426_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_01427_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01428_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01429_, _01428_, _01427_);
  or (_01430_, _01429_, _01426_);
  or (_01431_, _01430_, _01425_);
  and (_01432_, _01431_, _01423_);
  and (_01433_, _01432_, _01422_);
  and (_01434_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_01435_, _01434_, _00979_);
  and (_01436_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01438_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01439_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_01441_, _01439_, _01438_);
  or (_01442_, _01441_, _01436_);
  or (_01443_, _01442_, _01435_);
  and (_01445_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_01446_, _01445_, _40271_);
  and (_01447_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01449_, _01021_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01450_, _01012_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_01451_, _01450_, _01449_);
  or (_01453_, _01451_, _01447_);
  or (_01454_, _01453_, _01446_);
  and (_01455_, _01454_, _01323_);
  and (_01457_, _01455_, _01443_);
  or (_01458_, _01457_, _01433_);
  nor (_01459_, _01458_, _01413_);
  nand (_01461_, _01459_, _01331_);
  or (_01462_, _01461_, _01316_);
  or (_01463_, _01462_, _01027_);
  and (_01465_, _01323_, _38881_);
  nor (_01466_, _01331_, _29703_);
  nor (_01467_, _01466_, _01465_);
  and (_01469_, _01467_, _01463_);
  and (_01470_, _01016_, _38904_);
  and (_01471_, _01021_, _38987_);
  or (_01472_, _01471_, _40271_);
  and (_01473_, _01003_, _38965_);
  and (_01474_, _01012_, _38976_);
  or (_01475_, _01474_, _01473_);
  or (_01476_, _01475_, _01472_);
  and (_01477_, _01012_, _38927_);
  and (_01478_, _01021_, _38938_);
  or (_01479_, _01478_, _00979_);
  or (_01480_, _01479_, _01477_);
  and (_01481_, _01003_, _38915_);
  not (_01482_, _01007_);
  nor (_01483_, _01482_, _38954_);
  or (_01484_, _01483_, _01481_);
  or (_01485_, _01484_, _01480_);
  and (_01486_, _01485_, _01476_);
  or (_01487_, _01486_, _01470_);
  and (_01488_, _01487_, _01465_);
  not (_01489_, _01329_);
  nand (_01491_, _01326_, _01049_);
  and (_01492_, _01491_, _38701_);
  and (_01494_, _01492_, _42936_);
  and (_01495_, _01494_, _01489_);
  or (_01496_, _01495_, _01488_);
  or (_01498_, _01496_, _01469_);
  or (_01499_, _40271_, _40370_);
  nand (_01500_, _40271_, _38269_);
  and (_01502_, _01500_, _01021_);
  and (_01503_, _01502_, _01499_);
  or (_01504_, _40271_, _40434_);
  nand (_01506_, _40271_, _38285_);
  and (_01507_, _01506_, _01003_);
  and (_01508_, _01507_, _01504_);
  or (_01510_, _01508_, _01503_);
  nand (_01511_, _40271_, _38276_);
  or (_01512_, _40271_, _40226_);
  and (_01514_, _01512_, _01012_);
  and (_01515_, _01514_, _01511_);
  and (_01516_, _01016_, _40169_);
  and (_01518_, _01008_, _40301_);
  or (_01519_, _01518_, _01516_);
  or (_01520_, _01519_, _01515_);
  nor (_01522_, _01520_, _01510_);
  nand (_01523_, _01522_, _01495_);
  and (_01524_, _01523_, _41654_);
  and (_39521_, _01524_, _01498_);
  and (_01525_, _01003_, _40271_);
  and (_01526_, _01525_, _01323_);
  and (_01527_, _01526_, _38878_);
  and (_01528_, _01279_, _01008_);
  and (_01529_, _01528_, _38359_);
  and (_01530_, _01525_, _00978_);
  and (_01531_, _01530_, _38715_);
  or (_01532_, _01531_, _01529_);
  or (_01533_, _01532_, _01527_);
  and (_01534_, _01533_, _16098_);
  not (_01535_, _01016_);
  and (_01536_, _01535_, _38761_);
  and (_01537_, _01536_, _42936_);
  and (_01538_, _01525_, _01465_);
  or (_01539_, _01538_, _43028_);
  or (_01540_, _01539_, _01537_);
  or (_01541_, _01540_, _01534_);
  and (_01543_, _01214_, _01148_);
  and (_01544_, _40315_, _40271_);
  and (_01546_, _01544_, _01021_);
  and (_01547_, _01546_, _01543_);
  and (_01548_, _01547_, _38359_);
  nor (_01550_, _01548_, rst);
  and (_39522_, _01550_, _01541_);
  and (_01551_, _43026_, _25406_);
  and (_01553_, _01551_, _28497_);
  and (_01554_, _01526_, _38881_);
  nor (_01555_, _01554_, _01553_);
  and (_01557_, _01535_, _42936_);
  and (_01558_, _01557_, _38761_);
  nor (_01559_, _01558_, _01534_);
  and (_01561_, _01559_, _01555_);
  or (_01562_, _01561_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  not (_01563_, _01548_);
  and (_01565_, _40396_, _01079_);
  and (_01566_, _40466_, _40233_);
  and (_01567_, _01566_, _01565_);
  and (_01569_, _01525_, _40316_);
  and (_01570_, _01569_, _01567_);
  and (_01571_, _01570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_01573_, _01547_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_01574_, _01573_, _01571_);
  and (_01575_, _01569_, _01543_);
  and (_01576_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_01577_, _01148_, _01078_);
  and (_01578_, _01569_, _01577_);
  and (_01579_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_01580_, _01579_, _01576_);
  or (_01581_, _01580_, _01574_);
  and (_01582_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_01583_, _01544_, _01003_);
  and (_01584_, _01566_, _00977_);
  and (_01585_, _01584_, _01583_);
  and (_01586_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_01587_, _01586_, _01582_);
  and (_01588_, _01567_, _01583_);
  and (_01589_, _01588_, _01059_);
  and (_01590_, _01544_, _01012_);
  and (_01591_, _01590_, _01543_);
  and (_01592_, _01591_, _38309_);
  or (_01593_, _01592_, _01589_);
  or (_01595_, _01593_, _01587_);
  or (_01596_, _01595_, _01581_);
  and (_01598_, _01526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01599_, _01583_, _01577_);
  and (_01600_, _01599_, _01129_);
  and (_01602_, _40466_, _40232_);
  and (_01603_, _01565_, _01602_);
  and (_01604_, _01603_, _01583_);
  and (_01606_, _01604_, _01386_);
  or (_01607_, _01606_, _01600_);
  and (_01608_, _01530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01610_, _01583_, _01543_);
  and (_01611_, _01610_, _01293_);
  or (_01612_, _01611_, _01608_);
  or (_01614_, _01612_, _01607_);
  or (_01615_, _01614_, _01598_);
  nor (_01616_, _01615_, _01596_);
  nand (_01618_, _01561_, _01616_);
  and (_01619_, _01618_, _01563_);
  and (_01620_, _01619_, _01562_);
  nor (_01622_, _01563_, _28465_);
  or (_01623_, _01622_, _01620_);
  and (_39523_, _01623_, _41654_);
  and (_01625_, _01530_, _01001_);
  and (_01626_, _01525_, _01279_);
  and (_01627_, _01626_, _01252_);
  and (_01628_, _01525_, _01195_);
  and (_01629_, _01628_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_01630_, _01525_, _01215_);
  and (_01631_, _01630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_01632_, _01631_, _01629_);
  or (_01633_, _01632_, _01627_);
  and (_01634_, _01599_, _01171_);
  and (_01635_, _01547_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_01636_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_01637_, _01636_, _01635_);
  or (_01638_, _01637_, _01634_);
  and (_01639_, _01588_, _01109_);
  and (_01640_, _01591_, _40336_);
  or (_01641_, _01640_, _01639_);
  and (_01642_, _01570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01643_, _01583_, _01602_);
  and (_01644_, _01643_, _01565_);
  and (_01645_, _01644_, _01359_);
  or (_01647_, _01645_, _01642_);
  or (_01648_, _01647_, _01641_);
  and (_01650_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_01651_, _01526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_01652_, _01651_, _01650_);
  or (_01654_, _01652_, _01648_);
  or (_01655_, _01654_, _01638_);
  or (_01656_, _01655_, _01633_);
  or (_01658_, _01656_, _01541_);
  or (_01659_, _01658_, _01625_);
  or (_01660_, _01561_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_01662_, _01660_, _01659_);
  or (_01663_, _01662_, _01548_);
  nand (_01664_, _01548_, _29615_);
  and (_01666_, _01664_, _41654_);
  and (_39586_, _01666_, _01663_);
  or (_01667_, _01561_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_01669_, _01547_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_01670_, _01570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_01671_, _01670_, _01669_);
  and (_01673_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_01674_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_01675_, _01674_, _01673_);
  or (_01677_, _01675_, _01671_);
  and (_01678_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_01679_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_01680_, _01679_, _01678_);
  and (_01681_, _01588_, _01102_);
  and (_01682_, _01591_, _40529_);
  or (_01683_, _01682_, _01681_);
  or (_01684_, _01683_, _01680_);
  or (_01685_, _01684_, _01677_);
  and (_01686_, _01526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01687_, _01599_, _01156_);
  and (_01688_, _01604_, _01352_);
  or (_01689_, _01688_, _01687_);
  and (_01690_, _01530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_01691_, _01610_, _01274_);
  or (_01692_, _01691_, _01690_);
  or (_01693_, _01692_, _01689_);
  or (_01694_, _01693_, _01686_);
  nor (_01695_, _01694_, _01685_);
  nand (_01696_, _01695_, _01561_);
  and (_01697_, _01696_, _01563_);
  and (_01699_, _01697_, _01667_);
  nor (_01700_, _01563_, _30294_);
  or (_01702_, _01700_, _01699_);
  and (_39587_, _01702_, _41654_);
  or (_01703_, _01561_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_01705_, _01547_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_01706_, _01570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01707_, _01706_, _01705_);
  and (_01709_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_01710_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01711_, _01710_, _01709_);
  or (_01713_, _01711_, _01707_);
  and (_01714_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01715_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_01717_, _01715_, _01714_);
  and (_01718_, _01588_, _01087_);
  and (_01719_, _01591_, _40255_);
  or (_01721_, _01719_, _01718_);
  or (_01722_, _01721_, _01717_);
  or (_01723_, _01722_, _01713_);
  and (_01725_, _01526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01726_, _01599_, _01178_);
  and (_01727_, _01604_, _01337_);
  or (_01729_, _01727_, _01726_);
  and (_01730_, _01530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_01731_, _01610_, _01267_);
  or (_01732_, _01731_, _01730_);
  or (_01733_, _01732_, _01729_);
  or (_01734_, _01733_, _01725_);
  nor (_01735_, _01734_, _01723_);
  nand (_01736_, _01735_, _01561_);
  and (_01737_, _01736_, _01563_);
  and (_01738_, _01737_, _01703_);
  nor (_01739_, _01563_, _30993_);
  or (_01740_, _01739_, _01738_);
  and (_39589_, _01740_, _41654_);
  or (_01741_, _01561_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_01742_, _01570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_01743_, _01547_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_01744_, _01743_, _01742_);
  and (_01745_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_01746_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_01747_, _01746_, _01745_);
  or (_01748_, _01747_, _01744_);
  and (_01750_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_01751_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_01753_, _01751_, _01750_);
  and (_01754_, _01588_, _01095_);
  and (_01755_, _01591_, _40299_);
  or (_01757_, _01755_, _01754_);
  or (_01758_, _01757_, _01753_);
  or (_01759_, _01758_, _01748_);
  and (_01761_, _01526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01762_, _01599_, _01164_);
  and (_01763_, _01604_, _01345_);
  or (_01765_, _01763_, _01762_);
  and (_01766_, _01530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_01767_, _01610_, _01260_);
  or (_01769_, _01767_, _01766_);
  or (_01770_, _01769_, _01765_);
  or (_01771_, _01770_, _01761_);
  nor (_01773_, _01771_, _01759_);
  nand (_01774_, _01773_, _01561_);
  and (_01775_, _01774_, _01563_);
  and (_01777_, _01775_, _01741_);
  nor (_01778_, _01563_, _31724_);
  or (_01779_, _01778_, _01777_);
  and (_39590_, _01779_, _41654_);
  or (_01781_, _01561_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_01782_, _01547_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_01783_, _01570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01784_, _01783_, _01782_);
  and (_01785_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_01786_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01787_, _01786_, _01785_);
  or (_01788_, _01787_, _01784_);
  and (_01789_, _01588_, _01073_);
  and (_01790_, _01591_, _38341_);
  or (_01791_, _01790_, _01789_);
  and (_01792_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01793_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_01794_, _01793_, _01792_);
  or (_01795_, _01794_, _01791_);
  or (_01796_, _01795_, _01788_);
  and (_01797_, _01526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01798_, _01599_, _01136_);
  and (_01799_, _01604_, _01405_);
  or (_01800_, _01799_, _01798_);
  and (_01802_, _01530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01803_, _01610_, _01285_);
  or (_01805_, _01803_, _01802_);
  or (_01806_, _01805_, _01800_);
  or (_01807_, _01806_, _01797_);
  nor (_01809_, _01807_, _01796_);
  nand (_01810_, _01809_, _01561_);
  and (_01811_, _01810_, _01563_);
  and (_01813_, _01811_, _01781_);
  nor (_01814_, _01563_, _32486_);
  or (_01815_, _01814_, _01813_);
  and (_39591_, _01815_, _41654_);
  or (_01817_, _01561_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_01818_, _01570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01820_, _01547_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_01821_, _01820_, _01818_);
  and (_01822_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_01824_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01825_, _01824_, _01822_);
  or (_01826_, _01825_, _01821_);
  and (_01828_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_01829_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_01830_, _01829_, _01828_);
  and (_01832_, _01588_, _01066_);
  and (_01833_, _01591_, _40212_);
  or (_01834_, _01833_, _01832_);
  or (_01835_, _01834_, _01830_);
  or (_01836_, _01835_, _01826_);
  and (_01837_, _01526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01838_, _01599_, _01121_);
  and (_01839_, _01604_, _01396_);
  or (_01840_, _01839_, _01838_);
  and (_01841_, _01530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01842_, _01610_, _01307_);
  or (_01843_, _01842_, _01841_);
  or (_01844_, _01843_, _01840_);
  or (_01845_, _01844_, _01837_);
  nor (_01846_, _01845_, _01836_);
  nand (_01847_, _01846_, _01561_);
  and (_01848_, _01847_, _01563_);
  and (_01849_, _01848_, _01817_);
  nor (_01850_, _01563_, _33314_);
  or (_01851_, _01850_, _01849_);
  and (_39592_, _01851_, _41654_);
  or (_01853_, _01561_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_01854_, _01547_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01856_, _01570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_01857_, _01856_, _01854_);
  and (_01858_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_01860_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_01861_, _01860_, _01858_);
  or (_01862_, _01861_, _01857_);
  and (_01864_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01865_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_01866_, _01865_, _01864_);
  and (_01868_, _01588_, _01051_);
  and (_01869_, _01591_, _40393_);
  or (_01870_, _01869_, _01868_);
  or (_01872_, _01870_, _01866_);
  or (_01873_, _01872_, _01862_);
  and (_01874_, _01526_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01876_, _01599_, _01143_);
  and (_01877_, _01604_, _01377_);
  or (_01878_, _01877_, _01876_);
  and (_01880_, _01530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01881_, _01610_, _01300_);
  or (_01882_, _01881_, _01880_);
  or (_01884_, _01882_, _01878_);
  or (_01885_, _01884_, _01874_);
  nor (_01886_, _01885_, _01873_);
  nand (_01887_, _01886_, _01561_);
  and (_01888_, _01887_, _01563_);
  and (_01889_, _01888_, _01853_);
  nor (_01890_, _01563_, _34032_);
  or (_01891_, _01890_, _01889_);
  and (_39593_, _01891_, _41654_);
  and (_39636_, _40597_, _41654_);
  and (_39638_, _40728_, _41654_);
  nor (_39640_, _40271_, rst);
  and (_39655_, _40745_, _41654_);
  and (_39656_, _40758_, _41654_);
  and (_39657_, _40771_, _41654_);
  and (_39659_, _40781_, _41654_);
  and (_39660_, _40792_, _41654_);
  and (_39661_, _40801_, _41654_);
  and (_39662_, _40814_, _41654_);
  nor (_39663_, _40351_, rst);
  nor (_39664_, _40548_, rst);
  not (_01893_, _41903_);
  nor (_01895_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01896_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01897_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01896_);
  nor (_01899_, _01897_, _01895_);
  nor (_01900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01901_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01896_);
  nor (_01903_, _01901_, _01900_);
  nor (_01904_, _01903_, _01899_);
  not (_01905_, _01904_);
  nor (_01907_, _00149_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01908_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01896_);
  nor (_01909_, _01908_, _01907_);
  and (_01911_, _01909_, _01905_);
  nor (_01912_, _01909_, _01905_);
  nor (_01913_, _01912_, _01911_);
  nor (_01915_, _00170_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01916_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01896_);
  nor (_01917_, _01916_, _01915_);
  not (_01919_, _01917_);
  nor (_01920_, _01919_, _01911_);
  and (_01921_, _01919_, _01911_);
  nor (_01923_, _01921_, _01920_);
  nor (_01924_, _01923_, _01913_);
  not (_01925_, _01903_);
  and (_01926_, _01925_, _01899_);
  and (_01927_, _01926_, _01924_);
  and (_01928_, _01927_, _01893_);
  not (_01929_, _41985_);
  and (_01930_, _01903_, _01899_);
  and (_01931_, _01924_, _01930_);
  and (_01932_, _01931_, _01929_);
  not (_01933_, _41944_);
  nor (_01934_, _01925_, _01899_);
  and (_01935_, _01934_, _01924_);
  and (_01936_, _01935_, _01933_);
  or (_01937_, _01936_, _01932_);
  or (_01938_, _01937_, _01928_);
  not (_01939_, _41821_);
  and (_01940_, _01919_, _01913_);
  and (_01941_, _01940_, _01930_);
  and (_01942_, _01941_, _01939_);
  not (_01943_, _41862_);
  and (_01945_, _01940_, _01904_);
  and (_01946_, _01945_, _01943_);
  not (_01948_, _41780_);
  and (_01949_, _01940_, _01934_);
  and (_01950_, _01949_, _01948_);
  or (_01952_, _01950_, _01946_);
  or (_01953_, _01952_, _01942_);
  not (_01954_, _41560_);
  not (_01956_, _01913_);
  and (_01957_, _01923_, _01956_);
  and (_01958_, _01957_, _01926_);
  and (_01960_, _01958_, _01954_);
  not (_01961_, _41657_);
  and (_01962_, _01957_, _01930_);
  and (_01964_, _01962_, _01961_);
  or (_01965_, _01964_, _01960_);
  not (_01966_, _42149_);
  and (_01968_, _01920_, _01930_);
  and (_01969_, _01968_, _01966_);
  not (_01970_, _42108_);
  and (_01972_, _01934_, _01920_);
  and (_01973_, _01972_, _01970_);
  or (_01974_, _01973_, _01969_);
  not (_01976_, _42067_);
  and (_01977_, _01926_, _01920_);
  and (_01978_, _01977_, _01976_);
  not (_01979_, _41605_);
  and (_01980_, _01917_, _01909_);
  and (_01981_, _01980_, _01934_);
  and (_01982_, _01981_, _01979_);
  or (_01983_, _01982_, _01978_);
  or (_01984_, _01983_, _01974_);
  not (_01985_, _41739_);
  and (_01986_, _01940_, _01926_);
  and (_01987_, _01986_, _01985_);
  not (_01988_, _42190_);
  and (_01989_, _01980_, _01904_);
  and (_01990_, _01989_, _01988_);
  not (_01991_, _42026_);
  and (_01992_, _01917_, _01912_);
  and (_01993_, _01992_, _01991_);
  not (_01994_, _41698_);
  and (_01995_, _01919_, _01912_);
  and (_01996_, _01995_, _01994_);
  or (_01998_, _01996_, _01993_);
  or (_01999_, _01998_, _01990_);
  or (_02001_, _01999_, _01987_);
  or (_02002_, _02001_, _01984_);
  or (_02003_, _02002_, _01965_);
  or (_02005_, _02003_, _01953_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _02005_, _01938_);
  and (_02006_, _01958_, _01966_);
  and (_02008_, _01968_, _01976_);
  and (_02009_, _01972_, _01991_);
  or (_02010_, _02009_, _02008_);
  or (_02012_, _02010_, _02006_);
  and (_02013_, _01935_, _01943_);
  and (_02014_, _01981_, _01988_);
  or (_02016_, _02014_, _02013_);
  or (_02017_, _02016_, _02012_);
  and (_02018_, _01945_, _01948_);
  and (_02020_, _01949_, _01994_);
  and (_02021_, _01941_, _01985_);
  or (_02022_, _02021_, _02020_);
  or (_02024_, _02022_, _02018_);
  and (_02025_, _01927_, _01939_);
  and (_02026_, _01995_, _01979_);
  or (_02028_, _02026_, _02025_);
  or (_02029_, _02028_, _02024_);
  or (_02030_, _02029_, _02017_);
  and (_02031_, _01989_, _01970_);
  and (_02032_, _01962_, _01954_);
  and (_02033_, _01986_, _01961_);
  or (_02034_, _02033_, _02032_);
  and (_02035_, _01931_, _01893_);
  and (_02036_, _01977_, _01929_);
  and (_02037_, _01992_, _01933_);
  or (_02038_, _02037_, _02036_);
  or (_02039_, _02038_, _02035_);
  or (_02040_, _02039_, _02034_);
  or (_02041_, _02040_, _02031_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _02041_, _02030_);
  and (_02042_, _01958_, _01988_);
  and (_02043_, _01931_, _01933_);
  and (_02044_, _01927_, _01943_);
  or (_02045_, _02044_, _02043_);
  or (_02046_, _02045_, _02042_);
  and (_02047_, _01986_, _01994_);
  and (_02049_, _01949_, _01985_);
  or (_02050_, _02049_, _02047_);
  and (_02052_, _01941_, _01948_);
  or (_02053_, _02052_, _02050_);
  and (_02054_, _01972_, _01976_);
  and (_02056_, _01981_, _01954_);
  or (_02057_, _02056_, _02054_);
  and (_02058_, _01977_, _01991_);
  and (_02060_, _01989_, _01966_);
  or (_02061_, _02060_, _02058_);
  or (_02062_, _02061_, _02057_);
  and (_02064_, _01945_, _01939_);
  and (_02065_, _01968_, _01970_);
  and (_02066_, _01992_, _01929_);
  and (_02068_, _01995_, _01961_);
  or (_02069_, _02068_, _02066_);
  or (_02070_, _02069_, _02065_);
  or (_02072_, _02070_, _02064_);
  or (_02073_, _02072_, _02062_);
  and (_02074_, _01935_, _01893_);
  and (_02076_, _01962_, _01979_);
  or (_02077_, _02076_, _02074_);
  or (_02078_, _02077_, _02073_);
  or (_02080_, _02078_, _02053_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _02080_, _02046_);
  and (_02081_, _01935_, _01939_);
  and (_02082_, _01931_, _01943_);
  and (_02083_, _01958_, _01970_);
  or (_02084_, _02083_, _02082_);
  or (_02085_, _02084_, _02081_);
  and (_02086_, _01986_, _01979_);
  and (_02087_, _01941_, _01994_);
  and (_02088_, _01945_, _01985_);
  or (_02089_, _02088_, _02087_);
  or (_02090_, _02089_, _02086_);
  and (_02091_, _01977_, _01933_);
  and (_02092_, _01968_, _01991_);
  or (_02093_, _02092_, _02091_);
  and (_02094_, _01972_, _01929_);
  and (_02095_, _01989_, _01976_);
  or (_02096_, _02095_, _02094_);
  or (_02097_, _02096_, _02093_);
  and (_02098_, _01949_, _01961_);
  and (_02099_, _01981_, _01966_);
  and (_02101_, _01995_, _01954_);
  and (_02102_, _01992_, _01893_);
  or (_02104_, _02102_, _02101_);
  or (_02105_, _02104_, _02099_);
  or (_02106_, _02105_, _02098_);
  or (_02108_, _02106_, _02097_);
  and (_02109_, _01962_, _01988_);
  and (_02110_, _01927_, _01948_);
  or (_02112_, _02110_, _02109_);
  or (_02113_, _02112_, _02108_);
  or (_02114_, _02113_, _02090_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _02114_, _02085_);
  not (_02116_, _41565_);
  and (_02117_, _01962_, _02116_);
  not (_02119_, _41867_);
  and (_02120_, _01935_, _02119_);
  not (_02121_, _41826_);
  and (_02123_, _01927_, _02121_);
  or (_02124_, _02123_, _02120_);
  or (_02125_, _02124_, _02117_);
  not (_02127_, _41662_);
  and (_02128_, _01986_, _02127_);
  not (_02129_, _41703_);
  and (_02131_, _01949_, _02129_);
  not (_02132_, _41785_);
  and (_02133_, _01945_, _02132_);
  or (_02134_, _02133_, _02131_);
  or (_02135_, _02134_, _02128_);
  not (_02136_, _42195_);
  and (_02137_, _01981_, _02136_);
  not (_02138_, _42072_);
  and (_02139_, _01968_, _02138_);
  or (_02140_, _02139_, _02137_);
  not (_02141_, _42031_);
  and (_02142_, _01972_, _02141_);
  not (_02143_, _42113_);
  and (_02144_, _01989_, _02143_);
  or (_02145_, _02144_, _02142_);
  or (_02146_, _02145_, _02140_);
  not (_02147_, _41744_);
  and (_02148_, _01941_, _02147_);
  not (_02149_, _41990_);
  and (_02150_, _01977_, _02149_);
  not (_02151_, _41949_);
  and (_02153_, _01992_, _02151_);
  not (_02154_, _41613_);
  and (_02156_, _01995_, _02154_);
  or (_02157_, _02156_, _02153_);
  or (_02158_, _02157_, _02150_);
  or (_02160_, _02158_, _02148_);
  or (_02161_, _02160_, _02146_);
  not (_02162_, _41908_);
  and (_02164_, _01931_, _02162_);
  not (_02165_, _42154_);
  and (_02166_, _01958_, _02165_);
  or (_02168_, _02166_, _02164_);
  or (_02169_, _02168_, _02161_);
  or (_02170_, _02169_, _02135_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _02170_, _02125_);
  not (_02172_, _41570_);
  and (_02173_, _01962_, _02172_);
  not (_02175_, _41872_);
  and (_02176_, _01935_, _02175_);
  not (_02177_, _42159_);
  and (_02179_, _01958_, _02177_);
  or (_02180_, _02179_, _02176_);
  or (_02181_, _02180_, _02173_);
  not (_02183_, _41749_);
  and (_02184_, _01941_, _02183_);
  not (_02185_, _41667_);
  and (_02186_, _01986_, _02185_);
  not (_02187_, _41708_);
  and (_02188_, _01949_, _02187_);
  or (_02189_, _02188_, _02186_);
  or (_02190_, _02189_, _02184_);
  not (_02191_, _41995_);
  and (_02192_, _01977_, _02191_);
  not (_02193_, _42118_);
  and (_02194_, _01989_, _02193_);
  or (_02195_, _02194_, _02192_);
  not (_02196_, _42200_);
  and (_02197_, _01981_, _02196_);
  not (_02198_, _42036_);
  and (_02199_, _01972_, _02198_);
  or (_02200_, _02199_, _02197_);
  or (_02201_, _02200_, _02195_);
  not (_02202_, _41790_);
  and (_02203_, _01945_, _02202_);
  not (_02204_, _42077_);
  and (_02205_, _01968_, _02204_);
  not (_02206_, _41954_);
  and (_02207_, _01992_, _02206_);
  not (_02208_, _41618_);
  and (_02209_, _01995_, _02208_);
  or (_02210_, _02209_, _02207_);
  or (_02211_, _02210_, _02205_);
  or (_02212_, _02211_, _02203_);
  or (_02213_, _02212_, _02201_);
  not (_02214_, _41913_);
  and (_02215_, _01931_, _02214_);
  not (_02216_, _41831_);
  and (_02217_, _01927_, _02216_);
  or (_02218_, _02217_, _02215_);
  or (_02219_, _02218_, _02213_);
  or (_02220_, _02219_, _02190_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _02220_, _02181_);
  not (_02221_, _42164_);
  and (_02222_, _01958_, _02221_);
  not (_02223_, _42041_);
  and (_02224_, _01972_, _02223_);
  not (_02225_, _42082_);
  and (_02226_, _01968_, _02225_);
  or (_02227_, _02226_, _02224_);
  or (_02228_, _02227_, _02222_);
  not (_02229_, _41877_);
  and (_02230_, _01935_, _02229_);
  not (_02231_, _42205_);
  and (_02232_, _01981_, _02231_);
  or (_02233_, _02232_, _02230_);
  or (_02234_, _02233_, _02228_);
  not (_02235_, _41795_);
  and (_02236_, _01945_, _02235_);
  not (_02237_, _41713_);
  and (_02238_, _01949_, _02237_);
  not (_02239_, _41754_);
  and (_02240_, _01941_, _02239_);
  or (_02241_, _02240_, _02238_);
  or (_02242_, _02241_, _02236_);
  not (_02243_, _41836_);
  and (_02244_, _01927_, _02243_);
  not (_02245_, _41623_);
  and (_02246_, _01995_, _02245_);
  or (_02247_, _02246_, _02244_);
  or (_02248_, _02247_, _02242_);
  or (_02249_, _02248_, _02234_);
  not (_02250_, _42123_);
  and (_02251_, _01989_, _02250_);
  not (_02252_, _41575_);
  and (_02253_, _01962_, _02252_);
  not (_02254_, _41672_);
  and (_02255_, _01986_, _02254_);
  or (_02256_, _02255_, _02253_);
  not (_02257_, _41918_);
  and (_02258_, _01931_, _02257_);
  not (_02259_, _42000_);
  and (_02260_, _01977_, _02259_);
  not (_02261_, _41959_);
  and (_02262_, _01992_, _02261_);
  or (_02263_, _02262_, _02260_);
  or (_02264_, _02263_, _02258_);
  or (_02265_, _02264_, _02256_);
  or (_02266_, _02265_, _02251_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _02266_, _02249_);
  not (_02267_, _42169_);
  and (_02268_, _01958_, _02267_);
  not (_02269_, _42046_);
  and (_02270_, _01972_, _02269_);
  not (_02271_, _42087_);
  and (_02272_, _01968_, _02271_);
  or (_02273_, _02272_, _02270_);
  or (_02274_, _02273_, _02268_);
  not (_02275_, _41923_);
  and (_02276_, _01931_, _02275_);
  not (_02277_, _42210_);
  and (_02278_, _01981_, _02277_);
  or (_02279_, _02278_, _02276_);
  or (_02280_, _02279_, _02274_);
  not (_02281_, _41800_);
  and (_02282_, _01945_, _02281_);
  not (_02283_, _41759_);
  and (_02284_, _01941_, _02283_);
  not (_02285_, _41718_);
  and (_02286_, _01949_, _02285_);
  or (_02287_, _02286_, _02284_);
  or (_02288_, _02287_, _02282_);
  not (_02289_, _41841_);
  and (_02290_, _01927_, _02289_);
  not (_02291_, _41628_);
  and (_02292_, _01995_, _02291_);
  or (_02293_, _02292_, _02290_);
  or (_02294_, _02293_, _02288_);
  or (_02295_, _02294_, _02280_);
  not (_02296_, _42128_);
  and (_02297_, _01989_, _02296_);
  not (_02298_, _41677_);
  and (_02299_, _01986_, _02298_);
  not (_02300_, _41580_);
  and (_02301_, _01962_, _02300_);
  or (_02302_, _02301_, _02299_);
  not (_02303_, _41882_);
  and (_02304_, _01935_, _02303_);
  not (_02305_, _42005_);
  and (_02306_, _01977_, _02305_);
  not (_02307_, _41964_);
  and (_02308_, _01992_, _02307_);
  or (_02309_, _02308_, _02306_);
  or (_02310_, _02309_, _02304_);
  or (_02311_, _02310_, _02302_);
  or (_02312_, _02311_, _02297_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _02312_, _02295_);
  not (_02313_, _42174_);
  and (_02314_, _01958_, _02313_);
  not (_02315_, _42051_);
  and (_02316_, _01972_, _02315_);
  not (_02317_, _42092_);
  and (_02318_, _01968_, _02317_);
  or (_02319_, _02318_, _02316_);
  or (_02320_, _02319_, _02314_);
  not (_02321_, _41928_);
  and (_02322_, _01931_, _02321_);
  not (_02323_, _42215_);
  and (_02324_, _01981_, _02323_);
  or (_02325_, _02324_, _02322_);
  or (_02326_, _02325_, _02320_);
  not (_02327_, _41805_);
  and (_02328_, _01945_, _02327_);
  not (_02329_, _41764_);
  and (_02330_, _01941_, _02329_);
  not (_02331_, _41723_);
  and (_02332_, _01949_, _02331_);
  or (_02333_, _02332_, _02330_);
  or (_02334_, _02333_, _02328_);
  not (_02335_, _41846_);
  and (_02336_, _01927_, _02335_);
  not (_02337_, _41633_);
  and (_02338_, _01995_, _02337_);
  or (_02339_, _02338_, _02336_);
  or (_02340_, _02339_, _02334_);
  or (_02341_, _02340_, _02326_);
  not (_02342_, _42133_);
  and (_02343_, _01989_, _02342_);
  not (_02344_, _41682_);
  and (_02345_, _01986_, _02344_);
  not (_02346_, _41585_);
  and (_02347_, _01962_, _02346_);
  or (_02348_, _02347_, _02345_);
  not (_02349_, _41887_);
  and (_02350_, _01935_, _02349_);
  not (_02351_, _42010_);
  and (_02352_, _01977_, _02351_);
  not (_02353_, _41969_);
  and (_02354_, _01992_, _02353_);
  or (_02355_, _02354_, _02352_);
  or (_02356_, _02355_, _02350_);
  or (_02357_, _02356_, _02348_);
  or (_02358_, _02357_, _02343_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _02358_, _02341_);
  not (_02359_, _42179_);
  and (_02360_, _01958_, _02359_);
  not (_02361_, _42056_);
  and (_02362_, _01972_, _02361_);
  not (_02363_, _42097_);
  and (_02364_, _01968_, _02363_);
  or (_02365_, _02364_, _02362_);
  or (_02366_, _02365_, _02360_);
  not (_02367_, _41933_);
  and (_02368_, _01931_, _02367_);
  not (_02369_, _42220_);
  and (_02370_, _01981_, _02369_);
  or (_02371_, _02370_, _02368_);
  or (_02372_, _02371_, _02366_);
  not (_02373_, _41810_);
  and (_02374_, _01945_, _02373_);
  not (_02375_, _41769_);
  and (_02376_, _01941_, _02375_);
  not (_02377_, _41728_);
  and (_02378_, _01949_, _02377_);
  or (_02379_, _02378_, _02376_);
  or (_02380_, _02379_, _02374_);
  not (_02381_, _41851_);
  and (_02382_, _01927_, _02381_);
  not (_02383_, _41638_);
  and (_02384_, _01995_, _02383_);
  or (_02385_, _02384_, _02382_);
  or (_02386_, _02385_, _02380_);
  or (_02387_, _02386_, _02372_);
  not (_02388_, _42138_);
  and (_02389_, _01989_, _02388_);
  not (_02390_, _41687_);
  and (_02391_, _01986_, _02390_);
  not (_02392_, _41590_);
  and (_02393_, _01962_, _02392_);
  or (_02394_, _02393_, _02391_);
  not (_02395_, _41892_);
  and (_02396_, _01935_, _02395_);
  not (_02397_, _42015_);
  and (_02398_, _01977_, _02397_);
  not (_02399_, _41974_);
  and (_02400_, _01992_, _02399_);
  or (_02401_, _02400_, _02398_);
  or (_02402_, _02401_, _02396_);
  or (_02403_, _02402_, _02394_);
  or (_02404_, _02403_, _02389_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _02404_, _02387_);
  not (_02405_, _41938_);
  and (_02406_, _01931_, _02405_);
  not (_02407_, _41897_);
  and (_02408_, _01935_, _02407_);
  not (_02409_, _42184_);
  and (_02410_, _01958_, _02409_);
  or (_02411_, _02410_, _02408_);
  or (_02412_, _02411_, _02406_);
  not (_02413_, _41733_);
  and (_02414_, _01949_, _02413_);
  not (_02415_, _41774_);
  and (_02416_, _01941_, _02415_);
  not (_02417_, _41815_);
  and (_02418_, _01945_, _02417_);
  or (_02419_, _02418_, _02416_);
  or (_02420_, _02419_, _02414_);
  not (_02421_, _42102_);
  and (_02422_, _01968_, _02421_);
  not (_02423_, _42143_);
  and (_02424_, _01989_, _02423_);
  or (_02425_, _02424_, _02422_);
  not (_02426_, _42225_);
  and (_02428_, _01981_, _02426_);
  not (_02429_, _42020_);
  and (_02430_, _01977_, _02429_);
  or (_02431_, _02430_, _02428_);
  or (_02432_, _02431_, _02425_);
  not (_02433_, _41692_);
  and (_02434_, _01986_, _02433_);
  not (_02435_, _42061_);
  and (_02436_, _01972_, _02435_);
  not (_02437_, _41979_);
  and (_02438_, _01992_, _02437_);
  not (_02439_, _41646_);
  and (_02440_, _01995_, _02439_);
  or (_02441_, _02440_, _02438_);
  or (_02442_, _02441_, _02436_);
  or (_02443_, _02442_, _02434_);
  or (_02444_, _02443_, _02432_);
  not (_02445_, _41595_);
  and (_02446_, _01962_, _02445_);
  not (_02447_, _41856_);
  and (_02448_, _01927_, _02447_);
  or (_02449_, _02448_, _02446_);
  or (_02450_, _02449_, _02444_);
  or (_02451_, _02450_, _02420_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _02451_, _02412_);
  and (_02452_, _01931_, _02149_);
  and (_02453_, _01927_, _02162_);
  and (_02454_, _01958_, _02116_);
  or (_02455_, _02454_, _02453_);
  or (_02456_, _02455_, _02452_);
  and (_02457_, _01941_, _02121_);
  and (_02458_, _01945_, _02119_);
  and (_02459_, _01949_, _02132_);
  or (_02460_, _02459_, _02458_);
  or (_02461_, _02460_, _02457_);
  and (_02462_, _01968_, _02165_);
  and (_02463_, _01972_, _02143_);
  or (_02464_, _02463_, _02462_);
  and (_02465_, _01989_, _02136_);
  and (_02466_, _01977_, _02138_);
  or (_02467_, _02466_, _02465_);
  or (_02468_, _02467_, _02464_);
  and (_02469_, _01986_, _02147_);
  and (_02470_, _01981_, _02154_);
  and (_02471_, _01992_, _02141_);
  and (_02472_, _01995_, _02129_);
  or (_02473_, _02472_, _02471_);
  or (_02474_, _02473_, _02470_);
  or (_02475_, _02474_, _02469_);
  or (_02476_, _02475_, _02468_);
  and (_02477_, _01935_, _02151_);
  and (_02478_, _01962_, _02127_);
  or (_02479_, _02478_, _02477_);
  or (_02480_, _02479_, _02476_);
  or (_02481_, _02480_, _02461_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _02481_, _02456_);
  and (_02482_, _01977_, _02204_);
  and (_02483_, _01972_, _02193_);
  and (_02484_, _01968_, _02177_);
  or (_02485_, _02484_, _02483_);
  or (_02486_, _02485_, _02482_);
  and (_02487_, _01945_, _02175_);
  and (_02488_, _01992_, _02198_);
  or (_02489_, _02488_, _02487_);
  or (_02490_, _02489_, _02486_);
  and (_02491_, _01986_, _02183_);
  and (_02492_, _01949_, _02202_);
  and (_02493_, _01941_, _02216_);
  or (_02494_, _02493_, _02492_);
  or (_02495_, _02494_, _02491_);
  and (_02496_, _01981_, _02208_);
  and (_02497_, _01995_, _02187_);
  or (_02498_, _02497_, _02496_);
  or (_02499_, _02498_, _02495_);
  or (_02500_, _02499_, _02490_);
  and (_02501_, _01927_, _02214_);
  and (_02502_, _01931_, _02191_);
  and (_02503_, _01935_, _02206_);
  or (_02504_, _02503_, _02502_);
  or (_02505_, _02504_, _02501_);
  and (_02506_, _01958_, _02172_);
  and (_02507_, _01962_, _02185_);
  or (_02508_, _02507_, _02506_);
  and (_02509_, _01989_, _02196_);
  or (_02510_, _02509_, _02508_);
  or (_02511_, _02510_, _02505_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _02511_, _02500_);
  and (_02512_, _01927_, _02257_);
  and (_02513_, _01931_, _02259_);
  and (_02514_, _01935_, _02261_);
  or (_02515_, _02514_, _02513_);
  or (_02516_, _02515_, _02512_);
  and (_02517_, _01949_, _02235_);
  and (_02518_, _01945_, _02229_);
  and (_02519_, _01941_, _02243_);
  or (_02520_, _02519_, _02518_);
  or (_02521_, _02520_, _02517_);
  and (_02522_, _01958_, _02252_);
  and (_02523_, _01962_, _02254_);
  or (_02524_, _02523_, _02522_);
  and (_02525_, _01968_, _02221_);
  and (_02526_, _01977_, _02225_);
  or (_02527_, _02526_, _02525_);
  and (_02528_, _01972_, _02250_);
  and (_02529_, _01981_, _02245_);
  or (_02530_, _02529_, _02528_);
  or (_02531_, _02530_, _02527_);
  and (_02532_, _01986_, _02239_);
  and (_02533_, _01989_, _02231_);
  and (_02534_, _01992_, _02223_);
  and (_02535_, _01995_, _02237_);
  or (_02536_, _02535_, _02534_);
  or (_02537_, _02536_, _02533_);
  or (_02538_, _02537_, _02532_);
  or (_02539_, _02538_, _02531_);
  or (_02540_, _02539_, _02524_);
  or (_02541_, _02540_, _02521_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _02541_, _02516_);
  and (_02542_, _01968_, _02267_);
  and (_02543_, _01972_, _02296_);
  or (_02544_, _02543_, _02542_);
  and (_02545_, _01977_, _02271_);
  or (_02546_, _02545_, _02544_);
  and (_02547_, _01945_, _02303_);
  and (_02548_, _01992_, _02269_);
  or (_02549_, _02548_, _02547_);
  or (_02550_, _02549_, _02546_);
  and (_02551_, _01986_, _02283_);
  and (_02552_, _01949_, _02281_);
  and (_02553_, _01941_, _02289_);
  or (_02554_, _02553_, _02552_);
  or (_02555_, _02554_, _02551_);
  and (_02556_, _01981_, _02291_);
  and (_02557_, _01995_, _02285_);
  or (_02558_, _02557_, _02556_);
  or (_02559_, _02558_, _02555_);
  or (_02560_, _02559_, _02550_);
  and (_02561_, _01927_, _02275_);
  and (_02562_, _01935_, _02307_);
  and (_02563_, _01931_, _02305_);
  or (_02564_, _02563_, _02562_);
  or (_02565_, _02564_, _02561_);
  and (_02566_, _01989_, _02277_);
  and (_02567_, _01962_, _02298_);
  and (_02568_, _01958_, _02300_);
  or (_02569_, _02568_, _02567_);
  or (_02570_, _02569_, _02566_);
  or (_02571_, _02570_, _02565_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _02571_, _02560_);
  and (_02572_, _01927_, _02321_);
  and (_02573_, _01962_, _02344_);
  and (_02574_, _01931_, _02351_);
  or (_02575_, _02574_, _02573_);
  or (_02576_, _02575_, _02572_);
  and (_02577_, _01986_, _02329_);
  and (_02578_, _01949_, _02327_);
  and (_02579_, _01945_, _02349_);
  or (_02580_, _02579_, _02578_);
  or (_02581_, _02580_, _02577_);
  and (_02582_, _01972_, _02342_);
  and (_02583_, _01977_, _02317_);
  or (_02584_, _02583_, _02582_);
  and (_02585_, _01981_, _02337_);
  and (_02586_, _01968_, _02313_);
  or (_02587_, _02586_, _02585_);
  or (_02588_, _02587_, _02584_);
  and (_02589_, _01941_, _02335_);
  and (_02590_, _01989_, _02323_);
  and (_02591_, _01995_, _02331_);
  and (_02592_, _01992_, _02315_);
  or (_02593_, _02592_, _02591_);
  or (_02594_, _02593_, _02590_);
  or (_02595_, _02594_, _02589_);
  or (_02596_, _02595_, _02588_);
  and (_02597_, _01958_, _02346_);
  and (_02598_, _01935_, _02353_);
  or (_02599_, _02598_, _02597_);
  or (_02600_, _02599_, _02596_);
  or (_02601_, _02600_, _02581_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _02601_, _02576_);
  and (_02602_, _01931_, _02397_);
  and (_02603_, _01935_, _02399_);
  or (_02604_, _02603_, _02602_);
  and (_02605_, _01927_, _02367_);
  and (_02606_, _01945_, _02395_);
  or (_02607_, _02606_, _02605_);
  or (_02608_, _02607_, _02604_);
  and (_02609_, _01995_, _02377_);
  and (_02610_, _01941_, _02381_);
  and (_02611_, _01949_, _02373_);
  or (_02612_, _02611_, _02610_);
  or (_02613_, _02612_, _02609_);
  and (_02614_, _01986_, _02375_);
  and (_02615_, _01981_, _02383_);
  or (_02616_, _02615_, _02614_);
  or (_02617_, _02616_, _02613_);
  or (_02618_, _02617_, _02608_);
  and (_02619_, _01968_, _02359_);
  and (_02620_, _01972_, _02388_);
  or (_02621_, _02620_, _02619_);
  and (_02623_, _01977_, _02363_);
  and (_02624_, _01992_, _02361_);
  or (_02625_, _02624_, _02623_);
  or (_02626_, _02625_, _02621_);
  and (_02627_, _01958_, _02392_);
  and (_02628_, _01962_, _02390_);
  or (_02629_, _02628_, _02627_);
  and (_02630_, _01989_, _02369_);
  or (_02631_, _02630_, _02629_);
  or (_02632_, _02631_, _02626_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _02632_, _02618_);
  and (_02633_, _01935_, _02437_);
  and (_02634_, _01931_, _02429_);
  and (_02635_, _01927_, _02405_);
  or (_02636_, _02635_, _02634_);
  or (_02637_, _02636_, _02633_);
  and (_02638_, _01941_, _02447_);
  and (_02639_, _01945_, _02407_);
  and (_02640_, _01949_, _02417_);
  or (_02641_, _02640_, _02639_);
  or (_02642_, _02641_, _02638_);
  and (_02643_, _01958_, _02445_);
  and (_02644_, _01962_, _02433_);
  or (_02645_, _02644_, _02643_);
  and (_02646_, _01968_, _02409_);
  and (_02647_, _01977_, _02421_);
  or (_02648_, _02647_, _02646_);
  and (_02649_, _01972_, _02423_);
  and (_02650_, _01981_, _02439_);
  or (_02651_, _02650_, _02649_);
  or (_02652_, _02651_, _02648_);
  and (_02653_, _01986_, _02415_);
  and (_02654_, _01989_, _02426_);
  and (_02655_, _01992_, _02435_);
  and (_02656_, _01995_, _02413_);
  or (_02657_, _02656_, _02655_);
  or (_02658_, _02657_, _02654_);
  or (_02659_, _02658_, _02653_);
  or (_02660_, _02659_, _02652_);
  or (_02661_, _02660_, _02645_);
  or (_02662_, _02661_, _02642_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _02662_, _02637_);
  and (_02663_, _01958_, _02143_);
  and (_02664_, _01927_, _02132_);
  and (_02665_, _01935_, _02121_);
  or (_02666_, _02665_, _02664_);
  or (_02667_, _02666_, _02663_);
  and (_02668_, _01941_, _02129_);
  and (_02669_, _01949_, _02127_);
  and (_02670_, _01945_, _02147_);
  or (_02671_, _02670_, _02669_);
  or (_02672_, _02671_, _02668_);
  and (_02673_, _01968_, _02141_);
  and (_02674_, _01989_, _02138_);
  or (_02675_, _02674_, _02673_);
  and (_02676_, _01981_, _02165_);
  and (_02677_, _01972_, _02149_);
  or (_02678_, _02677_, _02676_);
  or (_02679_, _02678_, _02675_);
  and (_02680_, _01986_, _02154_);
  and (_02681_, _01977_, _02151_);
  and (_02682_, _01992_, _02162_);
  and (_02683_, _01995_, _02116_);
  or (_02684_, _02683_, _02682_);
  or (_02685_, _02684_, _02681_);
  or (_02686_, _02685_, _02680_);
  or (_02687_, _02686_, _02679_);
  and (_02688_, _01962_, _02136_);
  and (_02689_, _01931_, _02119_);
  or (_02690_, _02689_, _02688_);
  or (_02691_, _02690_, _02687_);
  or (_02692_, _02691_, _02672_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02692_, _02667_);
  and (_02693_, _01931_, _02175_);
  and (_02694_, _01972_, _02191_);
  and (_02695_, _01977_, _02206_);
  or (_02696_, _02695_, _02694_);
  or (_02697_, _02696_, _02693_);
  and (_02698_, _01968_, _02198_);
  and (_02699_, _01992_, _02214_);
  or (_02700_, _02699_, _02698_);
  or (_02701_, _02700_, _02697_);
  and (_02702_, _01935_, _02216_);
  and (_02703_, _01986_, _02208_);
  and (_02704_, _01949_, _02185_);
  and (_02705_, _01995_, _02172_);
  or (_02706_, _02705_, _02704_);
  or (_02707_, _02706_, _02703_);
  or (_02708_, _02707_, _02702_);
  or (_02709_, _02708_, _02701_);
  and (_02710_, _01958_, _02193_);
  and (_02711_, _01981_, _02177_);
  and (_02712_, _01962_, _02196_);
  or (_02713_, _02712_, _02711_);
  or (_02714_, _02713_, _02710_);
  and (_02715_, _01989_, _02204_);
  and (_02716_, _01927_, _02202_);
  and (_02717_, _01941_, _02187_);
  and (_02718_, _01945_, _02183_);
  or (_02719_, _02718_, _02717_);
  or (_02720_, _02719_, _02716_);
  or (_02721_, _02720_, _02715_);
  or (_02722_, _02721_, _02714_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02722_, _02709_);
  and (_02723_, _01958_, _02250_);
  and (_02724_, _01935_, _02243_);
  and (_02725_, _01931_, _02229_);
  or (_02726_, _02725_, _02724_);
  or (_02727_, _02726_, _02723_);
  and (_02728_, _01945_, _02239_);
  and (_02729_, _01949_, _02254_);
  and (_02730_, _01941_, _02237_);
  or (_02731_, _02730_, _02729_);
  or (_02732_, _02731_, _02728_);
  and (_02733_, _01977_, _02261_);
  and (_02734_, _01968_, _02223_);
  or (_02735_, _02734_, _02733_);
  and (_02736_, _01981_, _02221_);
  and (_02737_, _01989_, _02225_);
  or (_02738_, _02737_, _02736_);
  or (_02739_, _02738_, _02735_);
  and (_02740_, _01986_, _02245_);
  and (_02741_, _01972_, _02259_);
  and (_02742_, _01995_, _02252_);
  and (_02743_, _01992_, _02257_);
  or (_02744_, _02743_, _02742_);
  or (_02745_, _02744_, _02741_);
  or (_02746_, _02745_, _02740_);
  or (_02747_, _02746_, _02739_);
  and (_02748_, _01962_, _02231_);
  and (_02749_, _01927_, _02235_);
  or (_02750_, _02749_, _02748_);
  or (_02751_, _02750_, _02747_);
  or (_02752_, _02751_, _02732_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02752_, _02727_);
  and (_02753_, _01931_, _02303_);
  and (_02754_, _01972_, _02305_);
  and (_02755_, _01977_, _02307_);
  or (_02756_, _02755_, _02754_);
  or (_02757_, _02756_, _02753_);
  and (_02758_, _01968_, _02269_);
  and (_02759_, _01992_, _02275_);
  or (_02760_, _02759_, _02758_);
  or (_02761_, _02760_, _02757_);
  and (_02762_, _01935_, _02289_);
  and (_02763_, _01986_, _02291_);
  and (_02764_, _01949_, _02298_);
  and (_02765_, _01995_, _02300_);
  or (_02766_, _02765_, _02764_);
  or (_02767_, _02766_, _02763_);
  or (_02768_, _02767_, _02762_);
  or (_02769_, _02768_, _02761_);
  and (_02770_, _01958_, _02296_);
  and (_02771_, _01981_, _02267_);
  and (_02772_, _01962_, _02277_);
  or (_02773_, _02772_, _02771_);
  or (_02774_, _02773_, _02770_);
  and (_02775_, _01989_, _02271_);
  and (_02776_, _01927_, _02281_);
  and (_02777_, _01941_, _02285_);
  and (_02778_, _01945_, _02283_);
  or (_02779_, _02778_, _02777_);
  or (_02780_, _02779_, _02776_);
  or (_02781_, _02780_, _02775_);
  or (_02782_, _02781_, _02774_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02782_, _02769_);
  and (_02783_, _01958_, _02342_);
  and (_02784_, _01931_, _02349_);
  and (_02785_, _01935_, _02335_);
  or (_02786_, _02785_, _02784_);
  or (_02787_, _02786_, _02783_);
  and (_02788_, _01949_, _02344_);
  and (_02789_, _01986_, _02337_);
  and (_02790_, _01945_, _02329_);
  or (_02791_, _02790_, _02789_);
  or (_02792_, _02791_, _02788_);
  and (_02793_, _01981_, _02313_);
  and (_02794_, _01977_, _02353_);
  or (_02795_, _02794_, _02793_);
  and (_02796_, _01989_, _02317_);
  and (_02797_, _01972_, _02351_);
  or (_02798_, _02797_, _02796_);
  or (_02799_, _02798_, _02795_);
  and (_02800_, _01941_, _02331_);
  and (_02801_, _01968_, _02315_);
  and (_02802_, _01992_, _02321_);
  and (_02803_, _01995_, _02346_);
  or (_02804_, _02803_, _02802_);
  or (_02805_, _02804_, _02801_);
  or (_02806_, _02805_, _02800_);
  or (_02807_, _02806_, _02799_);
  and (_02808_, _01962_, _02323_);
  and (_02809_, _01927_, _02327_);
  or (_02810_, _02809_, _02808_);
  or (_02811_, _02810_, _02807_);
  or (_02812_, _02811_, _02792_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02812_, _02787_);
  and (_02813_, _01935_, _02381_);
  and (_02814_, _01931_, _02395_);
  and (_02815_, _01958_, _02388_);
  or (_02817_, _02815_, _02814_);
  or (_02818_, _02817_, _02813_);
  and (_02819_, _01986_, _02383_);
  and (_02820_, _01941_, _02377_);
  and (_02821_, _01945_, _02375_);
  or (_02822_, _02821_, _02820_);
  or (_02823_, _02822_, _02819_);
  and (_02824_, _01977_, _02399_);
  and (_02825_, _01968_, _02361_);
  or (_02826_, _02825_, _02824_);
  and (_02827_, _01972_, _02397_);
  and (_02828_, _01989_, _02363_);
  or (_02829_, _02828_, _02827_);
  or (_02830_, _02829_, _02826_);
  and (_02831_, _01949_, _02390_);
  and (_02832_, _01981_, _02359_);
  and (_02833_, _01995_, _02392_);
  and (_02834_, _01992_, _02367_);
  or (_02835_, _02834_, _02833_);
  or (_02836_, _02835_, _02832_);
  or (_02837_, _02836_, _02831_);
  or (_02838_, _02837_, _02830_);
  and (_02839_, _01962_, _02369_);
  and (_02840_, _01927_, _02373_);
  or (_02841_, _02840_, _02839_);
  or (_02842_, _02841_, _02838_);
  or (_02843_, _02842_, _02823_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02843_, _02818_);
  and (_02844_, _01931_, _02407_);
  and (_02845_, _01927_, _02417_);
  and (_02846_, _01958_, _02423_);
  or (_02847_, _02846_, _02845_);
  or (_02848_, _02847_, _02844_);
  and (_02849_, _01949_, _02433_);
  and (_02850_, _01986_, _02439_);
  and (_02851_, _01945_, _02415_);
  or (_02852_, _02851_, _02850_);
  or (_02853_, _02852_, _02849_);
  and (_02854_, _01972_, _02429_);
  and (_02855_, _01981_, _02409_);
  or (_02856_, _02855_, _02854_);
  and (_02857_, _01977_, _02437_);
  and (_02858_, _01968_, _02435_);
  or (_02859_, _02858_, _02857_);
  or (_02860_, _02859_, _02856_);
  and (_02861_, _01941_, _02413_);
  and (_02862_, _01989_, _02421_);
  and (_02863_, _01995_, _02445_);
  and (_02864_, _01992_, _02405_);
  or (_02865_, _02864_, _02863_);
  or (_02866_, _02865_, _02862_);
  or (_02867_, _02866_, _02861_);
  or (_02868_, _02867_, _02860_);
  and (_02869_, _01962_, _02426_);
  and (_02870_, _01935_, _02447_);
  or (_02871_, _02870_, _02869_);
  or (_02872_, _02871_, _02868_);
  or (_02873_, _02872_, _02853_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02873_, _02848_);
  and (_02874_, _01935_, _02162_);
  and (_02875_, _01931_, _02151_);
  and (_02876_, _01927_, _02119_);
  or (_02877_, _02876_, _02875_);
  or (_02878_, _02877_, _02874_);
  and (_02879_, _01949_, _02147_);
  and (_02880_, _01986_, _02129_);
  or (_02881_, _02880_, _02879_);
  and (_02882_, _01941_, _02132_);
  or (_02883_, _02882_, _02881_);
  and (_02884_, _01972_, _02138_);
  and (_02885_, _01977_, _02141_);
  or (_02886_, _02885_, _02884_);
  and (_02887_, _01968_, _02143_);
  and (_02888_, _01981_, _02116_);
  or (_02889_, _02888_, _02887_);
  or (_02890_, _02889_, _02886_);
  and (_02891_, _01945_, _02121_);
  and (_02892_, _01989_, _02165_);
  and (_02893_, _01992_, _02149_);
  and (_02894_, _01995_, _02127_);
  or (_02895_, _02894_, _02893_);
  or (_02896_, _02895_, _02892_);
  or (_02897_, _02896_, _02891_);
  or (_02898_, _02897_, _02890_);
  and (_02899_, _01958_, _02136_);
  and (_02900_, _01962_, _02154_);
  or (_02901_, _02900_, _02899_);
  or (_02902_, _02901_, _02898_);
  or (_02903_, _02902_, _02883_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _02903_, _02878_);
  and (_02904_, _01931_, _02206_);
  and (_02905_, _01992_, _02191_);
  or (_02906_, _02905_, _02904_);
  and (_02907_, _01935_, _02214_);
  and (_02908_, _01927_, _02175_);
  or (_02909_, _02908_, _02907_);
  or (_02910_, _02909_, _02906_);
  and (_02911_, _01958_, _02196_);
  and (_02912_, _01972_, _02204_);
  and (_02913_, _01977_, _02198_);
  or (_02914_, _02913_, _02912_);
  and (_02915_, _01968_, _02193_);
  or (_02916_, _02915_, _02914_);
  or (_02917_, _02916_, _02911_);
  or (_02918_, _02917_, _02910_);
  and (_02919_, _01962_, _02208_);
  and (_02920_, _01945_, _02216_);
  and (_02921_, _01941_, _02202_);
  or (_02922_, _02921_, _02920_);
  and (_02923_, _01949_, _02183_);
  and (_02924_, _01986_, _02187_);
  or (_02925_, _02924_, _02923_);
  or (_02926_, _02925_, _02922_);
  or (_02927_, _02926_, _02919_);
  and (_02928_, _01989_, _02177_);
  and (_02929_, _01981_, _02172_);
  and (_02930_, _01995_, _02185_);
  or (_02931_, _02930_, _02929_);
  or (_02932_, _02931_, _02928_);
  or (_02933_, _02932_, _02927_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _02933_, _02918_);
  and (_02934_, _01935_, _02257_);
  and (_02935_, _01958_, _02231_);
  and (_02936_, _01927_, _02229_);
  or (_02937_, _02936_, _02935_);
  or (_02938_, _02937_, _02934_);
  and (_02939_, _01945_, _02243_);
  and (_02940_, _01941_, _02235_);
  and (_02941_, _01986_, _02237_);
  or (_02942_, _02941_, _02940_);
  or (_02943_, _02942_, _02939_);
  and (_02944_, _01972_, _02225_);
  and (_02945_, _01977_, _02223_);
  or (_02946_, _02945_, _02944_);
  and (_02947_, _01968_, _02250_);
  and (_02948_, _01989_, _02221_);
  or (_02949_, _02948_, _02947_);
  or (_02950_, _02949_, _02946_);
  and (_02951_, _01949_, _02239_);
  and (_02952_, _01981_, _02252_);
  and (_02953_, _01995_, _02254_);
  and (_02954_, _01992_, _02259_);
  or (_02955_, _02954_, _02953_);
  or (_02956_, _02955_, _02952_);
  or (_02957_, _02956_, _02951_);
  or (_02958_, _02957_, _02950_);
  and (_02959_, _01962_, _02245_);
  and (_02960_, _01931_, _02261_);
  or (_02961_, _02960_, _02959_);
  or (_02962_, _02961_, _02958_);
  or (_02963_, _02962_, _02943_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _02963_, _02938_);
  and (_02964_, _01935_, _02275_);
  and (_02965_, _01962_, _02291_);
  and (_02966_, _01927_, _02303_);
  or (_02967_, _02966_, _02965_);
  or (_02968_, _02967_, _02964_);
  and (_02969_, _01941_, _02281_);
  and (_02970_, _01945_, _02289_);
  or (_02971_, _02970_, _02969_);
  and (_02973_, _01986_, _02285_);
  or (_02974_, _02973_, _02971_);
  and (_02975_, _01981_, _02300_);
  and (_02976_, _01968_, _02296_);
  or (_02977_, _02976_, _02975_);
  and (_02978_, _01977_, _02269_);
  and (_02979_, _01989_, _02267_);
  or (_02980_, _02979_, _02978_);
  or (_02981_, _02980_, _02977_);
  and (_02982_, _01949_, _02283_);
  and (_02984_, _01972_, _02271_);
  and (_02985_, _01995_, _02298_);
  and (_02986_, _01992_, _02305_);
  or (_02987_, _02986_, _02985_);
  or (_02988_, _02987_, _02984_);
  or (_02989_, _02988_, _02982_);
  or (_02990_, _02989_, _02981_);
  and (_02991_, _01958_, _02277_);
  and (_02992_, _01931_, _02307_);
  or (_02993_, _02992_, _02991_);
  or (_02994_, _02993_, _02990_);
  or (_02995_, _02994_, _02974_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02995_, _02968_);
  and (_02996_, _01935_, _02321_);
  and (_02997_, _01962_, _02337_);
  and (_02998_, _01927_, _02349_);
  or (_02999_, _02998_, _02997_);
  or (_03000_, _02999_, _02996_);
  and (_03001_, _01941_, _02327_);
  and (_03002_, _01945_, _02335_);
  or (_03004_, _03002_, _03001_);
  and (_03005_, _01986_, _02331_);
  or (_03006_, _03005_, _03004_);
  and (_03007_, _01981_, _02346_);
  and (_03008_, _01968_, _02342_);
  or (_03009_, _03008_, _03007_);
  and (_03010_, _01977_, _02315_);
  and (_03011_, _01989_, _02313_);
  or (_03012_, _03011_, _03010_);
  or (_03013_, _03012_, _03009_);
  and (_03015_, _01949_, _02329_);
  and (_03016_, _01972_, _02317_);
  and (_03017_, _01995_, _02344_);
  and (_03018_, _01992_, _02351_);
  or (_03019_, _03018_, _03017_);
  or (_03020_, _03019_, _03016_);
  or (_03021_, _03020_, _03015_);
  or (_03022_, _03021_, _03013_);
  and (_03023_, _01958_, _02323_);
  and (_03024_, _01931_, _02353_);
  or (_03026_, _03024_, _03023_);
  or (_03027_, _03026_, _03022_);
  or (_03028_, _03027_, _03006_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _03028_, _03000_);
  and (_03029_, _01935_, _02367_);
  and (_03030_, _01931_, _02399_);
  and (_03031_, _01927_, _02395_);
  or (_03032_, _03031_, _03030_);
  or (_03033_, _03032_, _03029_);
  and (_03034_, _01949_, _02375_);
  and (_03035_, _01986_, _02377_);
  or (_03036_, _03035_, _03034_);
  and (_03037_, _01941_, _02373_);
  or (_03038_, _03037_, _03036_);
  and (_03039_, _01972_, _02363_);
  and (_03040_, _01977_, _02361_);
  or (_03041_, _03040_, _03039_);
  and (_03042_, _01968_, _02388_);
  and (_03043_, _01981_, _02392_);
  or (_03044_, _03043_, _03042_);
  or (_03046_, _03044_, _03041_);
  and (_03047_, _01945_, _02381_);
  and (_03048_, _01989_, _02359_);
  and (_03049_, _01992_, _02397_);
  and (_03050_, _01995_, _02390_);
  or (_03051_, _03050_, _03049_);
  or (_03052_, _03051_, _03048_);
  or (_03053_, _03052_, _03047_);
  or (_03054_, _03053_, _03046_);
  and (_03055_, _01958_, _02369_);
  and (_03057_, _01962_, _02383_);
  or (_03058_, _03057_, _03055_);
  or (_03059_, _03058_, _03054_);
  or (_03060_, _03059_, _03038_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _03060_, _03033_);
  and (_03061_, _01935_, _02405_);
  and (_03062_, _01931_, _02437_);
  and (_03063_, _01927_, _02407_);
  or (_03064_, _03063_, _03062_);
  or (_03065_, _03064_, _03061_);
  and (_03067_, _01949_, _02415_);
  and (_03068_, _01986_, _02413_);
  or (_03069_, _03068_, _03067_);
  and (_03070_, _01941_, _02417_);
  or (_03071_, _03070_, _03069_);
  and (_03072_, _01972_, _02421_);
  and (_03073_, _01977_, _02435_);
  or (_03074_, _03073_, _03072_);
  and (_03075_, _01968_, _02423_);
  and (_03076_, _01981_, _02445_);
  or (_03078_, _03076_, _03075_);
  or (_03079_, _03078_, _03074_);
  and (_03080_, _01945_, _02447_);
  and (_03081_, _01989_, _02409_);
  and (_03082_, _01992_, _02429_);
  and (_03083_, _01995_, _02433_);
  or (_03084_, _03083_, _03082_);
  or (_03085_, _03084_, _03081_);
  or (_03086_, _03085_, _03080_);
  or (_03087_, _03086_, _03079_);
  and (_03089_, _01958_, _02426_);
  and (_03090_, _01962_, _02439_);
  or (_03091_, _03090_, _03089_);
  or (_03092_, _03091_, _03087_);
  or (_03093_, _03092_, _03071_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _03093_, _03065_);
  nand (_03094_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_03095_, \oc8051_golden_model_1.PC [3]);
  or (_03096_, \oc8051_golden_model_1.PC [2], _03095_);
  or (_03097_, _03096_, _03094_);
  or (_03099_, _03097_, _42061_);
  not (_03100_, \oc8051_golden_model_1.PC [1]);
  or (_03101_, _03100_, \oc8051_golden_model_1.PC [0]);
  or (_03102_, _03101_, _03096_);
  or (_03103_, _03102_, _42020_);
  and (_03104_, _03103_, _03099_);
  not (_03105_, \oc8051_golden_model_1.PC [2]);
  or (_03106_, _03105_, \oc8051_golden_model_1.PC [3]);
  or (_03107_, _03106_, _03094_);
  or (_03108_, _03107_, _41897_);
  or (_03110_, _03106_, _03101_);
  or (_03111_, _03110_, _41856_);
  and (_03112_, _03111_, _03108_);
  and (_03113_, _03112_, _03104_);
  nand (_03114_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_03115_, _03114_, _03094_);
  or (_03116_, _03115_, _42225_);
  or (_03117_, _03114_, _03101_);
  or (_03118_, _03117_, _42184_);
  and (_03119_, _03118_, _03116_);
  or (_03121_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_03122_, _03121_, _03094_);
  or (_03123_, _03122_, _41733_);
  or (_03124_, _03121_, _03101_);
  or (_03125_, _03124_, _41692_);
  and (_03126_, _03125_, _03123_);
  and (_03127_, _03126_, _03119_);
  and (_03128_, _03127_, _03113_);
  not (_03129_, \oc8051_golden_model_1.PC [0]);
  or (_03130_, \oc8051_golden_model_1.PC [1], _03129_);
  or (_03132_, _03130_, _03114_);
  or (_03133_, _03132_, _42143_);
  or (_03134_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_03135_, _03134_, _03114_);
  or (_03136_, _03135_, _42102_);
  and (_03137_, _03136_, _03133_);
  or (_03138_, _03121_, _03134_);
  or (_03139_, _03138_, _41595_);
  or (_03140_, _03121_, _03130_);
  or (_03141_, _03140_, _41646_);
  and (_03142_, _03141_, _03139_);
  and (_03143_, _03142_, _03137_);
  or (_03144_, _03130_, _03096_);
  or (_03145_, _03144_, _41979_);
  or (_03146_, _03134_, _03096_);
  or (_03147_, _03146_, _41938_);
  and (_03148_, _03147_, _03145_);
  or (_03149_, _03130_, _03106_);
  or (_03150_, _03149_, _41815_);
  or (_03151_, _03134_, _03106_);
  or (_03152_, _03151_, _41774_);
  and (_03153_, _03152_, _03150_);
  and (_03154_, _03153_, _03148_);
  and (_03155_, _03154_, _03143_);
  and (_03156_, _03155_, _03128_);
  or (_03157_, _03097_, _42026_);
  or (_03158_, _03102_, _41985_);
  and (_03159_, _03158_, _03157_);
  or (_03160_, _03107_, _41862_);
  or (_03161_, _03110_, _41821_);
  and (_03162_, _03161_, _03160_);
  and (_03163_, _03162_, _03159_);
  or (_03164_, _03115_, _42190_);
  or (_03165_, _03117_, _42149_);
  and (_03166_, _03165_, _03164_);
  or (_03167_, _03122_, _41698_);
  or (_03168_, _03124_, _41657_);
  and (_03169_, _03168_, _03167_);
  and (_03170_, _03169_, _03166_);
  and (_03171_, _03170_, _03163_);
  or (_03172_, _03132_, _42108_);
  or (_03173_, _03135_, _42067_);
  and (_03174_, _03173_, _03172_);
  or (_03175_, _03138_, _41560_);
  or (_03176_, _03140_, _41605_);
  and (_03177_, _03176_, _03175_);
  and (_03178_, _03177_, _03174_);
  or (_03179_, _03144_, _41944_);
  or (_03180_, _03146_, _41903_);
  and (_03181_, _03180_, _03179_);
  or (_03182_, _03149_, _41780_);
  or (_03183_, _03151_, _41739_);
  and (_03184_, _03183_, _03182_);
  and (_03185_, _03184_, _03181_);
  and (_03186_, _03185_, _03178_);
  and (_03187_, _03186_, _03171_);
  and (_03188_, _03187_, _03156_);
  or (_03189_, _03097_, _42051_);
  or (_03190_, _03102_, _42010_);
  and (_03191_, _03190_, _03189_);
  or (_03192_, _03107_, _41887_);
  or (_03193_, _03110_, _41846_);
  and (_03194_, _03193_, _03192_);
  and (_03195_, _03194_, _03191_);
  or (_03196_, _03115_, _42215_);
  or (_03197_, _03117_, _42174_);
  and (_03198_, _03197_, _03196_);
  or (_03199_, _03122_, _41723_);
  or (_03200_, _03124_, _41682_);
  and (_03201_, _03200_, _03199_);
  and (_03202_, _03201_, _03198_);
  and (_03203_, _03202_, _03195_);
  or (_03204_, _03132_, _42133_);
  or (_03205_, _03135_, _42092_);
  and (_03206_, _03205_, _03204_);
  or (_03207_, _03138_, _41585_);
  or (_03208_, _03140_, _41633_);
  and (_03209_, _03208_, _03207_);
  and (_03210_, _03209_, _03206_);
  or (_03211_, _03144_, _41969_);
  or (_03212_, _03146_, _41928_);
  and (_03213_, _03212_, _03211_);
  or (_03214_, _03149_, _41805_);
  or (_03215_, _03151_, _41764_);
  and (_03216_, _03215_, _03214_);
  and (_03217_, _03216_, _03213_);
  and (_03218_, _03217_, _03210_);
  and (_03219_, _03218_, _03203_);
  or (_03220_, _03097_, _42056_);
  or (_03221_, _03102_, _42015_);
  and (_03223_, _03221_, _03220_);
  or (_03224_, _03107_, _41892_);
  or (_03225_, _03110_, _41851_);
  and (_03226_, _03225_, _03224_);
  and (_03227_, _03226_, _03223_);
  or (_03228_, _03115_, _42220_);
  or (_03229_, _03117_, _42179_);
  and (_03230_, _03229_, _03228_);
  or (_03231_, _03122_, _41728_);
  or (_03232_, _03124_, _41687_);
  and (_03233_, _03232_, _03231_);
  and (_03234_, _03233_, _03230_);
  and (_03235_, _03234_, _03227_);
  or (_03236_, _03132_, _42138_);
  or (_03237_, _03135_, _42097_);
  and (_03238_, _03237_, _03236_);
  or (_03239_, _03138_, _41590_);
  or (_03240_, _03140_, _41638_);
  and (_03241_, _03240_, _03239_);
  and (_03242_, _03241_, _03238_);
  or (_03243_, _03144_, _41974_);
  or (_03244_, _03146_, _41933_);
  and (_03245_, _03244_, _03243_);
  or (_03246_, _03149_, _41810_);
  or (_03247_, _03151_, _41769_);
  and (_03248_, _03247_, _03246_);
  and (_03249_, _03248_, _03245_);
  and (_03250_, _03249_, _03242_);
  nand (_03251_, _03250_, _03235_);
  or (_03252_, _03251_, _03219_);
  not (_03253_, _03252_);
  and (_03254_, _03253_, _03188_);
  or (_03255_, _03097_, _42041_);
  or (_03256_, _03102_, _42000_);
  and (_03257_, _03256_, _03255_);
  or (_03258_, _03107_, _41877_);
  or (_03259_, _03110_, _41836_);
  and (_03260_, _03259_, _03258_);
  and (_03261_, _03260_, _03257_);
  or (_03262_, _03115_, _42205_);
  or (_03263_, _03117_, _42164_);
  and (_03264_, _03263_, _03262_);
  or (_03265_, _03122_, _41713_);
  or (_03266_, _03124_, _41672_);
  and (_03267_, _03266_, _03265_);
  and (_03268_, _03267_, _03264_);
  and (_03269_, _03268_, _03261_);
  or (_03270_, _03132_, _42123_);
  or (_03271_, _03135_, _42082_);
  and (_03272_, _03271_, _03270_);
  or (_03273_, _03138_, _41575_);
  or (_03274_, _03140_, _41623_);
  and (_03275_, _03274_, _03273_);
  and (_03276_, _03275_, _03272_);
  or (_03277_, _03144_, _41959_);
  or (_03278_, _03146_, _41918_);
  and (_03279_, _03278_, _03277_);
  or (_03280_, _03149_, _41795_);
  or (_03281_, _03151_, _41754_);
  and (_03282_, _03281_, _03280_);
  and (_03283_, _03282_, _03279_);
  and (_03284_, _03283_, _03276_);
  nand (_03285_, _03284_, _03269_);
  or (_03286_, _03097_, _42046_);
  or (_03287_, _03102_, _42005_);
  and (_03288_, _03287_, _03286_);
  or (_03289_, _03107_, _41882_);
  or (_03290_, _03110_, _41841_);
  and (_03291_, _03290_, _03289_);
  and (_03292_, _03291_, _03288_);
  or (_03293_, _03115_, _42210_);
  or (_03294_, _03117_, _42169_);
  and (_03295_, _03294_, _03293_);
  or (_03296_, _03122_, _41718_);
  or (_03297_, _03124_, _41677_);
  and (_03298_, _03297_, _03296_);
  and (_03299_, _03298_, _03295_);
  and (_03300_, _03299_, _03292_);
  or (_03301_, _03132_, _42128_);
  or (_03302_, _03135_, _42087_);
  and (_03303_, _03302_, _03301_);
  or (_03304_, _03138_, _41580_);
  or (_03305_, _03140_, _41628_);
  and (_03306_, _03305_, _03304_);
  and (_03307_, _03306_, _03303_);
  or (_03308_, _03144_, _41964_);
  or (_03309_, _03146_, _41923_);
  and (_03310_, _03309_, _03308_);
  or (_03311_, _03149_, _41800_);
  or (_03312_, _03151_, _41759_);
  and (_03313_, _03312_, _03311_);
  and (_03314_, _03313_, _03310_);
  and (_03315_, _03314_, _03307_);
  nand (_03316_, _03315_, _03300_);
  or (_03317_, _03316_, _03285_);
  not (_03318_, _03317_);
  or (_03319_, _03097_, _42031_);
  or (_03320_, _03102_, _41990_);
  and (_03321_, _03320_, _03319_);
  or (_03322_, _03107_, _41867_);
  or (_03323_, _03110_, _41826_);
  and (_03324_, _03323_, _03322_);
  and (_03325_, _03324_, _03321_);
  or (_03326_, _03115_, _42195_);
  or (_03327_, _03117_, _42154_);
  and (_03328_, _03327_, _03326_);
  or (_03329_, _03122_, _41703_);
  or (_03330_, _03124_, _41662_);
  and (_03331_, _03330_, _03329_);
  and (_03332_, _03331_, _03328_);
  and (_03333_, _03332_, _03325_);
  or (_03334_, _03132_, _42113_);
  or (_03335_, _03135_, _42072_);
  and (_03336_, _03335_, _03334_);
  or (_03337_, _03138_, _41565_);
  or (_03338_, _03140_, _41613_);
  and (_03339_, _03338_, _03337_);
  and (_03340_, _03339_, _03336_);
  or (_03341_, _03144_, _41949_);
  or (_03342_, _03146_, _41908_);
  and (_03343_, _03342_, _03341_);
  or (_03344_, _03149_, _41785_);
  or (_03345_, _03151_, _41744_);
  and (_03346_, _03345_, _03344_);
  and (_03347_, _03346_, _03343_);
  and (_03348_, _03347_, _03340_);
  and (_03349_, _03348_, _03333_);
  or (_03350_, _03097_, _42036_);
  or (_03351_, _03102_, _41995_);
  and (_03352_, _03351_, _03350_);
  or (_03353_, _03107_, _41872_);
  or (_03354_, _03110_, _41831_);
  and (_03355_, _03354_, _03353_);
  and (_03356_, _03355_, _03352_);
  or (_03357_, _03115_, _42200_);
  or (_03358_, _03117_, _42159_);
  and (_03359_, _03358_, _03357_);
  or (_03360_, _03122_, _41708_);
  or (_03361_, _03124_, _41667_);
  and (_03362_, _03361_, _03360_);
  and (_03363_, _03362_, _03359_);
  and (_03364_, _03363_, _03356_);
  or (_03365_, _03132_, _42118_);
  or (_03366_, _03135_, _42077_);
  and (_03367_, _03366_, _03365_);
  or (_03368_, _03138_, _41570_);
  or (_03369_, _03140_, _41618_);
  and (_03370_, _03369_, _03368_);
  and (_03371_, _03370_, _03367_);
  or (_03372_, _03144_, _41954_);
  or (_03373_, _03146_, _41913_);
  and (_03374_, _03373_, _03372_);
  or (_03375_, _03149_, _41790_);
  or (_03376_, _03151_, _41749_);
  and (_03377_, _03376_, _03375_);
  and (_03378_, _03377_, _03374_);
  and (_03379_, _03378_, _03371_);
  nand (_03380_, _03379_, _03364_);
  not (_03381_, _03380_);
  and (_03382_, _03381_, _03349_);
  and (_03383_, _03382_, _03318_);
  and (_03384_, _03383_, _03254_);
  not (_03385_, _03384_);
  or (_03386_, _03380_, _03349_);
  or (_03387_, _03386_, _03317_);
  not (_03388_, _03387_);
  nand (_03389_, _03218_, _03203_);
  and (_03390_, _03250_, _03235_);
  or (_03391_, _03390_, _03389_);
  not (_03392_, _03391_);
  and (_03393_, _03392_, _03188_);
  and (_03394_, _03393_, _03388_);
  not (_03395_, _03394_);
  or (_03396_, _03251_, _03389_);
  not (_03397_, _03396_);
  and (_03398_, _03397_, _03188_);
  and (_03399_, _03398_, _03388_);
  and (_03400_, _03388_, _03254_);
  nor (_03401_, _03400_, _03399_);
  nand (_03402_, _03401_, _03395_);
  and (_03403_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03404_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03405_, _03404_, _03403_);
  and (_03406_, _03405_, _03402_);
  not (_03407_, _03406_);
  nand (_03408_, _03155_, _03128_);
  or (_03409_, _03187_, _03408_);
  nor (_03410_, _03409_, _03396_);
  not (_03411_, _03410_);
  not (_03412_, _03285_);
  or (_03413_, _03316_, _03412_);
  or (_03414_, _03413_, _03386_);
  or (_03415_, _03414_, _03411_);
  nor (_03416_, _03409_, _03252_);
  not (_03417_, _03416_);
  or (_03418_, _03417_, _03387_);
  and (_03419_, _03418_, _03415_);
  or (_03420_, _03381_, _03349_);
  or (_03421_, _03420_, _03317_);
  or (_03422_, _03421_, _03417_);
  and (_03424_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_03425_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03426_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_03427_, _03426_, _03424_);
  and (_03428_, _03427_, _03425_);
  nor (_03429_, _03428_, _03424_);
  and (_03430_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_03431_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_03432_, _03431_, _03430_);
  not (_03433_, _03432_);
  nor (_03434_, _03433_, _03429_);
  and (_03435_, _03433_, _03429_);
  nor (_03436_, _03435_, _03434_);
  not (_03437_, _03436_);
  or (_03438_, _03437_, _03422_);
  and (_03439_, _03438_, _03419_);
  or (_03440_, _03390_, _03219_);
  or (_03441_, _03440_, _03409_);
  or (_03442_, _03441_, _03387_);
  or (_03443_, _03187_, _03156_);
  or (_03444_, _03443_, _03252_);
  or (_03445_, _03444_, _03387_);
  and (_03446_, _03445_, _03442_);
  or (_03447_, _03443_, _03396_);
  or (_03448_, _03447_, _03387_);
  or (_03449_, _03443_, _03391_);
  or (_03450_, _03449_, _03387_);
  and (_03451_, _03450_, _03448_);
  or (_03452_, _03409_, _03391_);
  or (_03453_, _03452_, _03387_);
  or (_03454_, _03443_, _03440_);
  or (_03455_, _03454_, _03387_);
  and (_03456_, _03455_, _03453_);
  and (_03457_, _03456_, _03451_);
  and (_03458_, _03457_, _03446_);
  nor (_03459_, _03094_, _03105_);
  and (_03460_, _03094_, _03105_);
  nor (_03461_, _03460_, _03459_);
  not (_03462_, _03461_);
  nand (_03463_, _03462_, _03458_);
  nand (_03464_, _03463_, _03422_);
  nand (_03465_, _03464_, _03439_);
  nor (_03466_, _03421_, _03411_);
  not (_03467_, _03466_);
  and (_03468_, _03458_, _03419_);
  or (_03469_, _03468_, _03405_);
  and (_03470_, _03469_, _03467_);
  nand (_03471_, _03470_, _03465_);
  not (_03472_, _03440_);
  and (_03473_, _03472_, _03188_);
  and (_03474_, _03473_, _03388_);
  and (_03475_, _03187_, _03408_);
  and (_03476_, _03475_, _03253_);
  and (_03477_, _03476_, _03388_);
  nor (_03478_, _03477_, _03474_);
  not (_03479_, _03478_);
  and (_03480_, _03475_, _03397_);
  and (_03481_, _03480_, _03388_);
  and (_03482_, _03475_, _03472_);
  and (_03483_, _03482_, _03388_);
  or (_03484_, _03483_, _03481_);
  and (_03485_, _03475_, _03392_);
  and (_03486_, _03485_, _03388_);
  and (_03487_, _03410_, _03388_);
  or (_03488_, _03487_, _03486_);
  or (_03489_, _03488_, _03484_);
  or (_03490_, _03489_, _03479_);
  not (_03491_, \oc8051_golden_model_1.ACC [1]);
  and (_03492_, _03130_, _03101_);
  nor (_03493_, _03492_, _03491_);
  and (_03494_, \oc8051_golden_model_1.ACC [0], _03129_);
  and (_03495_, _03492_, _03491_);
  nor (_03496_, _03495_, _03493_);
  and (_03497_, _03496_, _03494_);
  nor (_03498_, _03497_, _03493_);
  and (_03499_, _03461_, \oc8051_golden_model_1.ACC [2]);
  nor (_03500_, _03461_, \oc8051_golden_model_1.ACC [2]);
  nor (_03501_, _03500_, _03499_);
  not (_03502_, _03501_);
  nor (_03503_, _03502_, _03498_);
  and (_03504_, _03502_, _03498_);
  nor (_03505_, _03504_, _03503_);
  and (_03506_, _03505_, _03466_);
  nor (_03507_, _03506_, _03490_);
  nand (_03508_, _03507_, _03471_);
  nor (_03509_, _03490_, _03402_);
  or (_03510_, _03509_, _03405_);
  nand (_03511_, _03510_, _03508_);
  and (_03512_, _03511_, _03407_);
  and (_03513_, _03509_, _03468_);
  nor (_03514_, _03114_, _03100_);
  nor (_03515_, _03403_, \oc8051_golden_model_1.PC [3]);
  nor (_03516_, _03515_, _03514_);
  or (_03517_, _03516_, _03513_);
  and (_03518_, _03467_, _03419_);
  nor (_03519_, _03434_, _03430_);
  and (_03520_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03521_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03522_, _03521_, _03520_);
  not (_03523_, _03522_);
  nor (_03524_, _03523_, _03519_);
  and (_03525_, _03523_, _03519_);
  nor (_03526_, _03525_, _03524_);
  or (_03527_, _03526_, _03422_);
  not (_03528_, _03107_);
  nor (_03529_, _03459_, _03095_);
  nor (_03530_, _03529_, _03528_);
  and (_03531_, _03422_, _03530_);
  nand (_03532_, _03531_, _03458_);
  nand (_03533_, _03532_, _03527_);
  and (_03534_, _03533_, _03518_);
  nor (_03535_, _03503_, _03499_);
  nor (_03536_, _03530_, \oc8051_golden_model_1.ACC [3]);
  and (_03537_, _03530_, \oc8051_golden_model_1.ACC [3]);
  nor (_03538_, _03537_, _03536_);
  and (_03539_, _03538_, _03535_);
  nor (_03540_, _03538_, _03535_);
  nor (_03541_, _03540_, _03539_);
  nor (_03542_, _03541_, _03467_);
  or (_03543_, _03542_, _03534_);
  nand (_03544_, _03543_, _03509_);
  nand (_03545_, _03544_, _03517_);
  or (_03546_, _03545_, _03512_);
  not (_03547_, _03422_);
  nor (_03548_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03549_, _03548_, _03425_);
  nand (_03550_, _03549_, _03547_);
  and (_03551_, _03422_, _03129_);
  nand (_03552_, _03551_, _03458_);
  nand (_03553_, _03552_, _03550_);
  nand (_03554_, _03553_, _03419_);
  or (_03555_, _03468_, _03129_);
  nand (_03556_, _03555_, _03554_);
  nand (_03557_, _03556_, _03467_);
  not (_03558_, \oc8051_golden_model_1.ACC [0]);
  and (_03559_, _03558_, \oc8051_golden_model_1.PC [0]);
  or (_03560_, _03494_, _03467_);
  or (_03561_, _03560_, _03559_);
  and (_03562_, _03561_, _03509_);
  nand (_03563_, _03562_, _03557_);
  or (_03564_, _03509_, \oc8051_golden_model_1.PC [0]);
  nand (_03565_, _03564_, _03563_);
  or (_03566_, _03513_, _03100_);
  nor (_03567_, _03427_, _03425_);
  nor (_03568_, _03567_, _03428_);
  or (_03569_, _03568_, _03422_);
  and (_03570_, _03492_, _03422_);
  nand (_03571_, _03570_, _03458_);
  nand (_03572_, _03571_, _03569_);
  and (_03573_, _03572_, _03518_);
  nor (_03574_, _03496_, _03494_);
  nor (_03575_, _03574_, _03497_);
  nor (_03576_, _03575_, _03467_);
  or (_03577_, _03576_, _03573_);
  nand (_03578_, _03577_, _03509_);
  nand (_03579_, _03578_, _03566_);
  or (_03580_, _03579_, _03565_);
  or (_03581_, _03580_, _03546_);
  or (_03582_, _03581_, _42190_);
  nand (_03583_, _03511_, _03407_);
  or (_03584_, _03545_, _03583_);
  or (_03585_, _03584_, _03580_);
  or (_03586_, _03585_, _42026_);
  and (_03587_, _03586_, _03582_);
  and (_03588_, _03578_, _03566_);
  or (_03589_, _03588_, _03565_);
  and (_03590_, _03544_, _03517_);
  or (_03591_, _03590_, _03512_);
  or (_03592_, _03591_, _03589_);
  or (_03593_, _03592_, _41780_);
  and (_03594_, _03564_, _03563_);
  or (_03595_, _03579_, _03594_);
  or (_03596_, _03590_, _03583_);
  or (_03597_, _03596_, _03595_);
  or (_03598_, _03597_, _41657_);
  and (_03599_, _03598_, _03593_);
  and (_03600_, _03599_, _03587_);
  or (_03601_, _03595_, _03546_);
  or (_03602_, _03601_, _42149_);
  or (_03603_, _03589_, _03546_);
  or (_03604_, _03603_, _42108_);
  and (_03605_, _03604_, _03602_);
  or (_03606_, _03584_, _03595_);
  or (_03607_, _03606_, _41985_);
  or (_03608_, _03584_, _03589_);
  or (_03609_, _03608_, _41944_);
  and (_03610_, _03609_, _03607_);
  and (_03611_, _03610_, _03605_);
  and (_03612_, _03611_, _03600_);
  or (_03613_, _03588_, _03594_);
  or (_03614_, _03591_, _03613_);
  or (_03615_, _03614_, _41739_);
  or (_03616_, _03596_, _03580_);
  or (_03617_, _03616_, _41698_);
  and (_03618_, _03617_, _03615_);
  or (_03619_, _03591_, _03580_);
  or (_03620_, _03619_, _41862_);
  or (_03621_, _03596_, _03613_);
  or (_03622_, _03621_, _41560_);
  and (_03623_, _03622_, _03620_);
  and (_03625_, _03623_, _03618_);
  or (_03626_, _03613_, _03546_);
  or (_03627_, _03626_, _42067_);
  or (_03628_, _03613_, _03584_);
  or (_03629_, _03628_, _41903_);
  and (_03630_, _03629_, _03627_);
  or (_03631_, _03591_, _03595_);
  or (_03632_, _03631_, _41821_);
  or (_03633_, _03596_, _03589_);
  or (_03634_, _03633_, _41605_);
  and (_03635_, _03634_, _03632_);
  and (_03636_, _03635_, _03630_);
  and (_03637_, _03636_, _03625_);
  nand (_03638_, _03637_, _03612_);
  or (_03639_, _03603_, _42128_);
  or (_03640_, _03619_, _41882_);
  and (_03641_, _03640_, _03639_);
  or (_03642_, _03631_, _41841_);
  or (_03643_, _03621_, _41580_);
  and (_03644_, _03643_, _03642_);
  and (_03645_, _03644_, _03641_);
  or (_03646_, _03585_, _42046_);
  or (_03647_, _03616_, _41718_);
  and (_03648_, _03647_, _03646_);
  or (_03649_, _03606_, _42005_);
  or (_03650_, _03628_, _41923_);
  and (_03651_, _03650_, _03649_);
  and (_03652_, _03651_, _03648_);
  and (_03653_, _03652_, _03645_);
  or (_03654_, _03592_, _41800_);
  or (_03655_, _03614_, _41759_);
  and (_03656_, _03655_, _03654_);
  or (_03657_, _03581_, _42210_);
  or (_03658_, _03633_, _41628_);
  and (_03659_, _03658_, _03657_);
  and (_03660_, _03659_, _03656_);
  or (_03661_, _03601_, _42169_);
  or (_03662_, _03597_, _41677_);
  and (_03663_, _03662_, _03661_);
  or (_03664_, _03626_, _42087_);
  or (_03665_, _03608_, _41964_);
  and (_03666_, _03665_, _03664_);
  and (_03667_, _03666_, _03663_);
  and (_03668_, _03667_, _03660_);
  and (_03669_, _03668_, _03653_);
  or (_03670_, _03669_, _03638_);
  nor (_03671_, _03670_, _03385_);
  nor (_03672_, _03638_, _03385_);
  not (_03673_, _03672_);
  not (_03674_, \oc8051_golden_model_1.SP [0]);
  and (_03675_, _03474_, _03674_);
  not (_03676_, _03418_);
  and (_03677_, _03380_, _03349_);
  and (_03678_, _03677_, _03318_);
  and (_03679_, _03678_, _03416_);
  not (_03680_, _03679_);
  nor (_03681_, _03680_, _03670_);
  nor (_03682_, _03442_, _03674_);
  not (_03683_, _03441_);
  and (_03684_, _03678_, _03683_);
  not (_03685_, _03684_);
  nor (_03686_, _03685_, _03670_);
  nor (_03687_, _03685_, _03638_);
  not (_03688_, _03687_);
  not (_03689_, _03447_);
  and (_03690_, _03689_, _03383_);
  and (_03691_, _03678_, _03689_);
  not (_03692_, _03691_);
  nor (_03693_, _03692_, _03670_);
  nor (_03694_, _03692_, _03638_);
  not (_03695_, _03444_);
  and (_03696_, _03678_, _03695_);
  not (_03697_, _03696_);
  or (_03698_, _03697_, _03670_);
  not (_03699_, _03455_);
  not (_03700_, _03414_);
  and (_03701_, _03700_, _03398_);
  not (_03702_, _03701_);
  and (_03703_, _03700_, _03254_);
  not (_03704_, _03703_);
  and (_03705_, _03393_, _03383_);
  not (_03706_, _03705_);
  and (_03707_, _03678_, _03393_);
  not (_03708_, _03707_);
  and (_03709_, _03700_, _03393_);
  nor (_03710_, _03619_, _41897_);
  nor (_03711_, _03616_, _41733_);
  nor (_03712_, _03711_, _03710_);
  nor (_03713_, _03601_, _42184_);
  nor (_03714_, _03628_, _41938_);
  nor (_03715_, _03714_, _03713_);
  and (_03716_, _03715_, _03712_);
  nor (_03717_, _03631_, _41856_);
  nor (_03718_, _03592_, _41815_);
  nor (_03719_, _03718_, _03717_);
  nor (_03720_, _03597_, _41692_);
  nor (_03721_, _03633_, _41646_);
  nor (_03722_, _03721_, _03720_);
  and (_03723_, _03722_, _03719_);
  and (_03724_, _03723_, _03716_);
  nor (_03725_, _03603_, _42143_);
  nor (_03726_, _03585_, _42061_);
  nor (_03727_, _03726_, _03725_);
  nor (_03728_, _03581_, _42225_);
  nor (_03729_, _03626_, _42102_);
  nor (_03730_, _03729_, _03728_);
  and (_03731_, _03730_, _03727_);
  nor (_03732_, _03606_, _42020_);
  nor (_03733_, _03608_, _41979_);
  nor (_03734_, _03733_, _03732_);
  nor (_03735_, _03614_, _41774_);
  nor (_03736_, _03621_, _41595_);
  nor (_03737_, _03736_, _03735_);
  and (_03738_, _03737_, _03734_);
  and (_03739_, _03738_, _03731_);
  and (_03740_, _03739_, _03724_);
  nor (_03741_, _03740_, _03638_);
  not (_03742_, _03669_);
  and (_03743_, _03742_, _03638_);
  nor (_03744_, _03743_, _03741_);
  and (_03745_, _03678_, _03482_);
  and (_03746_, _03678_, _03410_);
  nor (_03747_, _03746_, _03745_);
  not (_03748_, _03747_);
  and (_03749_, _03748_, _03744_);
  nor (_03750_, _03447_, _03414_);
  not (_03751_, _03750_);
  nor (_03752_, _03751_, _03669_);
  nand (_03753_, _03696_, _03744_);
  not (_03754_, \oc8051_golden_model_1.SP [3]);
  and (_03755_, _03695_, _03383_);
  nand (_03756_, _03755_, _03754_);
  nor (_03757_, _03444_, _03414_);
  nor (_03758_, _03449_, _03414_);
  nor (_03759_, _03758_, _03757_);
  nor (_03760_, _03759_, _03669_);
  nor (_03761_, _03755_, _03696_);
  not (_03762_, _03761_);
  and (_03763_, _03759_, \oc8051_golden_model_1.PSW [3]);
  or (_03764_, _03763_, _03762_);
  and (_03765_, _03764_, _03751_);
  or (_03766_, _03765_, _03760_);
  and (_03767_, _03766_, _03756_);
  or (_03768_, _03767_, _03691_);
  and (_03769_, _03768_, _03753_);
  or (_03770_, _03769_, _03752_);
  nand (_03771_, _03744_, _03691_);
  nand (_03772_, _03771_, _03770_);
  nor (_03773_, _03441_, _03414_);
  nor (_03774_, _03773_, _03690_);
  nand (_03775_, _03774_, _03772_);
  or (_03776_, _03774_, _03742_);
  and (_03777_, _03683_, _03383_);
  nor (_03778_, _03684_, _03777_);
  and (_03779_, _03778_, _03776_);
  and (_03780_, _03779_, _03775_);
  nor (_03781_, _03778_, _03744_);
  nor (_03782_, _03781_, _03780_);
  not (_03783_, _03452_);
  not (_03784_, _03386_);
  and (_03785_, _03316_, _03412_);
  and (_03786_, _03785_, _03784_);
  and (_03787_, _03786_, _03783_);
  not (_03788_, _03787_);
  and (_03789_, _03785_, _03382_);
  and (_03790_, _03789_, _03783_);
  and (_03791_, _03785_, _03677_);
  and (_03792_, _03791_, _03783_);
  nor (_03793_, _03792_, _03790_);
  nand (_03794_, _03793_, _03788_);
  not (_03795_, _03794_);
  not (_03796_, _03420_);
  and (_03797_, _03785_, _03796_);
  and (_03798_, _03797_, _03783_);
  and (_03799_, _03316_, _03285_);
  and (_03800_, _03799_, _03381_);
  and (_03801_, _03800_, _03783_);
  nor (_03802_, _03801_, _03798_);
  and (_03803_, _03799_, _03380_);
  and (_03804_, _03803_, _03783_);
  not (_03805_, _03804_);
  and (_03806_, _03805_, _03802_);
  and (_03807_, _03806_, _03795_);
  not (_03808_, _03807_);
  nor (_03809_, _03808_, _03782_);
  and (_03810_, _03783_, _03383_);
  and (_03811_, _03678_, _03783_);
  nor (_03812_, _03811_, _03810_);
  not (_03813_, _03812_);
  nor (_03814_, _03807_, _03669_);
  nor (_03815_, _03814_, _03813_);
  not (_03816_, _03815_);
  nor (_03817_, _03816_, _03809_);
  nor (_03818_, _03417_, _03414_);
  and (_03819_, _03813_, _03744_);
  nor (_03820_, _03819_, _03818_);
  not (_03821_, _03820_);
  nor (_03822_, _03821_, _03817_);
  not (_03823_, _03818_);
  nor (_03824_, _03823_, _03669_);
  or (_03826_, _03824_, _03822_);
  and (_03827_, _03826_, _03680_);
  nor (_03828_, _03744_, _03680_);
  or (_03829_, _03828_, _03827_);
  and (_03830_, _03829_, _03415_);
  and (_03831_, _03473_, _03383_);
  nor (_03832_, _03705_, _03831_);
  and (_03833_, _03678_, _03254_);
  not (_03834_, _03421_);
  and (_03835_, _03480_, _03834_);
  nor (_03836_, _03835_, _03833_);
  and (_03837_, _03836_, _03832_);
  and (_03838_, _03485_, _03834_);
  and (_03839_, _03482_, _03700_);
  nor (_03840_, _03839_, _03838_);
  and (_03841_, _03678_, _03398_);
  nor (_03842_, _03841_, _03384_);
  and (_03843_, _03842_, _03840_);
  and (_03844_, _03843_, _03837_);
  not (_03845_, _03413_);
  and (_03846_, _03845_, _03382_);
  and (_03847_, _03846_, _03683_);
  nor (_03848_, _03847_, _03773_);
  not (_03849_, _03799_);
  nor (_03850_, _03849_, _03420_);
  and (_03851_, _03850_, _03683_);
  nor (_03852_, _03851_, _03757_);
  nor (_03853_, _03413_, _03381_);
  and (_03854_, _03853_, _03683_);
  not (_03855_, _03854_);
  and (_03856_, _03855_, _03852_);
  and (_03857_, _03856_, _03848_);
  and (_03858_, _03785_, _03381_);
  and (_03859_, _03858_, _03683_);
  not (_03860_, _03859_);
  and (_03861_, _03416_, _03383_);
  and (_03862_, _03799_, _03677_);
  and (_03863_, _03862_, _03683_);
  nor (_03864_, _03863_, _03861_);
  and (_03865_, _03864_, _03860_);
  and (_03866_, _03476_, _03834_);
  and (_03867_, _03785_, _03380_);
  and (_03868_, _03867_, _03683_);
  nor (_03869_, _03868_, _03866_);
  and (_03870_, _03800_, _03683_);
  not (_03871_, _03870_);
  and (_03872_, _03871_, _03869_);
  and (_03873_, _03872_, _03865_);
  and (_03874_, _03873_, _03857_);
  and (_03875_, _03874_, _03844_);
  nor (_03876_, _03875_, _03405_);
  and (_03877_, _03875_, _03462_);
  nor (_03878_, _03877_, _03876_);
  not (_03879_, _03516_);
  nor (_03880_, _03875_, _03879_);
  not (_03881_, _03530_);
  and (_03882_, _03875_, _03881_);
  nor (_03883_, _03882_, _03880_);
  not (_03884_, _03883_);
  and (_03885_, _03884_, _03878_);
  nor (_03886_, _03875_, _03129_);
  and (_03887_, _03875_, _03129_);
  nor (_03888_, _03887_, _03886_);
  not (_03889_, _03888_);
  nor (_03890_, _03887_, _03100_);
  and (_03891_, _03887_, _03100_);
  nor (_03892_, _03891_, _03890_);
  nor (_03893_, _03892_, _03889_);
  and (_03894_, _03893_, _03885_);
  and (_03895_, _03894_, _02271_);
  nor (_03896_, _03883_, _03878_);
  and (_03897_, _03892_, _03889_);
  and (_03898_, _03897_, _03896_);
  and (_03899_, _03898_, _02269_);
  nor (_03900_, _03899_, _03895_);
  and (_03901_, _03892_, _03888_);
  and (_03902_, _03883_, _03878_);
  and (_03903_, _03902_, _03901_);
  and (_03904_, _03903_, _02289_);
  nor (_03905_, _03892_, _03888_);
  nor (_03906_, _03884_, _03878_);
  and (_03907_, _03906_, _03905_);
  and (_03908_, _03907_, _02291_);
  nor (_03909_, _03908_, _03904_);
  and (_03910_, _03909_, _03900_);
  and (_03911_, _03901_, _03885_);
  and (_03912_, _03911_, _02267_);
  and (_03913_, _03905_, _03885_);
  and (_03914_, _03913_, _02296_);
  nor (_03915_, _03914_, _03912_);
  and (_03916_, _03901_, _03896_);
  and (_03917_, _03916_, _02305_);
  and (_03918_, _03905_, _03896_);
  and (_03919_, _03918_, _02307_);
  nor (_03920_, _03919_, _03917_);
  and (_03921_, _03920_, _03915_);
  and (_03922_, _03921_, _03910_);
  and (_03923_, _03902_, _03893_);
  and (_03924_, _03923_, _02283_);
  and (_03925_, _03906_, _03897_);
  and (_03926_, _03925_, _02285_);
  nor (_03927_, _03926_, _03924_);
  and (_03928_, _03902_, _03897_);
  and (_03929_, _03928_, _02303_);
  and (_03930_, _03905_, _03902_);
  and (_03931_, _03930_, _02281_);
  nor (_03932_, _03931_, _03929_);
  and (_03933_, _03932_, _03927_);
  and (_03934_, _03897_, _03885_);
  and (_03935_, _03934_, _02277_);
  and (_03936_, _03896_, _03893_);
  and (_03937_, _03936_, _02275_);
  nor (_03938_, _03937_, _03935_);
  and (_03939_, _03906_, _03893_);
  and (_03940_, _03939_, _02300_);
  and (_03941_, _03906_, _03901_);
  and (_03942_, _03941_, _02298_);
  nor (_03943_, _03942_, _03940_);
  and (_03944_, _03943_, _03938_);
  and (_03945_, _03944_, _03933_);
  and (_03946_, _03945_, _03922_);
  nor (_03947_, _03946_, _03415_);
  nor (_03948_, _03947_, _03748_);
  not (_03949_, _03948_);
  nor (_03950_, _03949_, _03830_);
  nor (_03951_, _03950_, _03749_);
  and (_03952_, _03480_, _03700_);
  not (_03953_, _03952_);
  and (_03954_, _03678_, _03480_);
  nor (_03955_, _03954_, _03835_);
  and (_03956_, _03955_, _03953_);
  and (_03957_, _03485_, _03700_);
  not (_03958_, _03957_);
  and (_03959_, _03678_, _03485_);
  nor (_03960_, _03959_, _03838_);
  and (_03961_, _03960_, _03958_);
  and (_03962_, _03961_, _03956_);
  and (_03963_, _03473_, _03700_);
  not (_03964_, _03963_);
  and (_03965_, _03476_, _03700_);
  not (_03966_, _03965_);
  and (_03967_, _03678_, _03476_);
  nor (_03968_, _03967_, _03866_);
  and (_03969_, _03968_, _03966_);
  and (_03970_, _03969_, _03964_);
  and (_03971_, _03970_, _03962_);
  not (_03972_, _03971_);
  nor (_03973_, _03972_, _03951_);
  and (_03974_, _03678_, _03473_);
  and (_03975_, _03972_, _03669_);
  nor (_03976_, _03975_, _03974_);
  not (_03977_, _03976_);
  nor (_03978_, _03977_, _03973_);
  and (_03979_, _03974_, \oc8051_golden_model_1.SP [3]);
  or (_03980_, _03979_, _03831_);
  or (_03981_, _03980_, _03978_);
  nand (_03982_, _03744_, _03831_);
  and (_03983_, _03982_, _03981_);
  nor (_03984_, _03983_, _03709_);
  and (_03985_, _03709_, _03669_);
  nor (_03986_, _03985_, _03984_);
  and (_03987_, _03986_, _03708_);
  and (_03988_, _03707_, \oc8051_golden_model_1.SP [3]);
  or (_03989_, _03988_, _03987_);
  and (_03990_, _03989_, _03706_);
  nor (_03991_, _03706_, _03744_);
  or (_03992_, _03991_, _03990_);
  and (_03993_, _03992_, _03704_);
  nor (_03994_, _03704_, _03669_);
  or (_03995_, _03994_, _03993_);
  and (_03996_, _03995_, _03385_);
  nor (_03997_, _03744_, _03385_);
  or (_03998_, _03997_, _03996_);
  nand (_03999_, _03998_, _03702_);
  nor (_04000_, _03702_, _03669_);
  not (_04001_, _04000_);
  and (_04002_, _04001_, _03999_);
  nor (_04003_, _03581_, _42220_);
  nor (_04004_, _03585_, _42056_);
  nor (_04005_, _04004_, _04003_);
  nor (_04006_, _03631_, _41851_);
  nor (_04007_, _03614_, _41769_);
  nor (_04008_, _04007_, _04006_);
  and (_04009_, _04008_, _04005_);
  nor (_04010_, _03601_, _42179_);
  nor (_04011_, _03603_, _42138_);
  nor (_04012_, _04011_, _04010_);
  nor (_04013_, _03606_, _42015_);
  nor (_04014_, _03628_, _41933_);
  nor (_04015_, _04014_, _04013_);
  and (_04016_, _04015_, _04012_);
  and (_04017_, _04016_, _04009_);
  nor (_04018_, _03621_, _41590_);
  nor (_04019_, _03597_, _41687_);
  nor (_04020_, _04019_, _04018_);
  nor (_04021_, _03619_, _41892_);
  nor (_04022_, _03592_, _41810_);
  nor (_04023_, _04022_, _04021_);
  and (_04024_, _04023_, _04020_);
  nor (_04025_, _03626_, _42097_);
  nor (_04027_, _03608_, _41974_);
  nor (_04028_, _04027_, _04025_);
  nor (_04029_, _03616_, _41728_);
  nor (_04030_, _03633_, _41638_);
  nor (_04031_, _04030_, _04029_);
  and (_04032_, _04031_, _04028_);
  and (_04033_, _04032_, _04024_);
  and (_04034_, _04033_, _04017_);
  nor (_04035_, _04034_, _03638_);
  nor (_04036_, _03696_, _03679_);
  and (_04037_, _04036_, _03692_);
  and (_04038_, _03778_, _03747_);
  and (_04039_, _03832_, _03812_);
  and (_04040_, _04039_, _04038_);
  and (_04041_, _04040_, _04037_);
  not (_04042_, _04041_);
  and (_04043_, _04042_, _04035_);
  not (_04044_, _04043_);
  and (_04045_, _04035_, _03384_);
  not (_04046_, _04045_);
  and (_04047_, _03918_, _02261_);
  and (_04048_, _03930_, _02235_);
  nor (_04049_, _04048_, _04047_);
  and (_04050_, _03934_, _02231_);
  and (_04051_, _03928_, _02229_);
  nor (_04052_, _04051_, _04050_);
  and (_04053_, _04052_, _04049_);
  and (_04054_, _03936_, _02257_);
  and (_04055_, _03923_, _02239_);
  nor (_04056_, _04055_, _04054_);
  and (_04057_, _03925_, _02237_);
  and (_04058_, _03907_, _02245_);
  nor (_04059_, _04058_, _04057_);
  and (_04060_, _04059_, _04056_);
  and (_04061_, _04060_, _04053_);
  and (_04062_, _03913_, _02250_);
  and (_04063_, _03916_, _02259_);
  nor (_04064_, _04063_, _04062_);
  and (_04065_, _03903_, _02243_);
  and (_04066_, _03941_, _02254_);
  nor (_04067_, _04066_, _04065_);
  and (_04068_, _04067_, _04064_);
  and (_04069_, _03898_, _02223_);
  and (_04070_, _03894_, _02225_);
  nor (_04071_, _04070_, _04069_);
  and (_04072_, _03911_, _02221_);
  and (_04073_, _03939_, _02252_);
  nor (_04074_, _04073_, _04072_);
  and (_04075_, _04074_, _04071_);
  and (_04076_, _04075_, _04068_);
  and (_04077_, _04076_, _04061_);
  nor (_04078_, _04077_, _03415_);
  not (_04079_, _03398_);
  nor (_04080_, _03480_, _03410_);
  and (_04081_, _04080_, _04079_);
  and (_04082_, _03441_, _03417_);
  not (_04083_, _03349_);
  nor (_04084_, _03449_, _04083_);
  not (_04085_, _04084_);
  and (_04086_, _04085_, _04082_);
  and (_04087_, _04086_, _04081_);
  nor (_04088_, _04087_, _03380_);
  and (_04089_, _03473_, _03380_);
  nor (_04090_, _04089_, _03485_);
  not (_04091_, _04090_);
  nor (_04092_, _04091_, _04088_);
  nor (_04093_, _04092_, _03849_);
  not (_04094_, _04093_);
  and (_04095_, _03803_, _03476_);
  and (_04096_, _03803_, _03410_);
  nor (_04097_, _04096_, _04095_);
  not (_04098_, _04097_);
  not (_04099_, _03803_);
  and (_04100_, _03390_, _03188_);
  not (_04101_, _04100_);
  and (_04102_, _04101_, _04082_);
  nor (_04103_, _04102_, _04099_);
  nor (_04104_, _04103_, _04098_);
  and (_04105_, _03800_, _03473_);
  and (_04106_, _03799_, _03393_);
  nor (_04107_, _04106_, _04105_);
  not (_04108_, _03449_);
  and (_04109_, _03803_, _04108_);
  and (_04110_, _03799_, _03784_);
  and (_04111_, _04110_, _04108_);
  or (_04112_, _04111_, _04109_);
  nor (_04113_, _03443_, _03251_);
  and (_04114_, _04113_, _03799_);
  nor (_04115_, _04114_, _04112_);
  and (_04116_, _04115_, _04107_);
  and (_04117_, _03755_, \oc8051_golden_model_1.SP [2]);
  not (_04118_, _04117_);
  and (_04119_, _03803_, _03480_);
  and (_04120_, _03800_, _03254_);
  nor (_04121_, _04120_, _04119_);
  and (_04122_, _04121_, _04118_);
  and (_04123_, _04122_, _04116_);
  and (_04124_, _03800_, _03476_);
  not (_04125_, \oc8051_golden_model_1.SP [2]);
  nor (_04126_, _03974_, _03707_);
  nor (_04128_, _04126_, _04125_);
  nor (_04129_, _04128_, _04124_);
  and (_04130_, _04129_, _04123_);
  and (_04131_, _04130_, _04104_);
  and (_04132_, _04131_, _04094_);
  not (_04133_, _04132_);
  nor (_04134_, _04133_, _04078_);
  nor (_04135_, _03581_, _42205_);
  nor (_04136_, _03621_, _41575_);
  nor (_04137_, _04136_, _04135_);
  nor (_04138_, _03585_, _42041_);
  nor (_04139_, _03616_, _41713_);
  nor (_04140_, _04139_, _04138_);
  and (_04141_, _04140_, _04137_);
  nor (_04142_, _03628_, _41918_);
  nor (_04143_, _03597_, _41672_);
  nor (_04144_, _04143_, _04142_);
  nor (_04145_, _03619_, _41877_);
  nor (_04146_, _03614_, _41754_);
  nor (_04147_, _04146_, _04145_);
  and (_04148_, _04147_, _04144_);
  and (_04149_, _04148_, _04141_);
  nor (_04150_, _03592_, _41795_);
  nor (_04151_, _03633_, _41623_);
  nor (_04152_, _04151_, _04150_);
  nor (_04153_, _03601_, _42164_);
  nor (_04154_, _03606_, _42000_);
  nor (_04155_, _04154_, _04153_);
  and (_04156_, _04155_, _04152_);
  nor (_04157_, _03626_, _42082_);
  nor (_04158_, _03608_, _41959_);
  nor (_04159_, _04158_, _04157_);
  nor (_04160_, _03603_, _42123_);
  nor (_04161_, _03631_, _41836_);
  nor (_04162_, _04161_, _04160_);
  and (_04163_, _04162_, _04159_);
  and (_04164_, _04163_, _04156_);
  and (_04165_, _04164_, _04149_);
  not (_04166_, _03709_);
  nor (_04167_, _03818_, _03750_);
  and (_04168_, _04167_, _04166_);
  and (_04169_, _03774_, _03759_);
  nor (_04170_, _03703_, _03701_);
  and (_04171_, _04170_, _04169_);
  and (_04172_, _04171_, _04168_);
  and (_04173_, _04172_, _03971_);
  and (_04174_, _04173_, _03807_);
  nor (_04175_, _04174_, _04165_);
  not (_04176_, _04175_);
  and (_04177_, _04176_, _04134_);
  and (_04178_, _04177_, _04046_);
  and (_04179_, _04178_, _04044_);
  not (_04180_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_04181_, _03616_, _41703_);
  or (_04182_, _03597_, _41662_);
  and (_04183_, _04182_, _04181_);
  or (_04184_, _03631_, _41826_);
  or (_04185_, _03614_, _41744_);
  and (_04186_, _04185_, _04184_);
  and (_04187_, _04186_, _04183_);
  or (_04188_, _03603_, _42113_);
  or (_04189_, _03608_, _41949_);
  and (_04190_, _04189_, _04188_);
  or (_04191_, _03585_, _42031_);
  or (_04192_, _03628_, _41908_);
  and (_04193_, _04192_, _04191_);
  and (_04194_, _04193_, _04190_);
  and (_04195_, _04194_, _04187_);
  or (_04196_, _03621_, _41565_);
  or (_04197_, _03633_, _41613_);
  and (_04198_, _04197_, _04196_);
  or (_04199_, _03619_, _41867_);
  or (_04200_, _03592_, _41785_);
  and (_04201_, _04200_, _04199_);
  and (_04202_, _04201_, _04198_);
  or (_04203_, _03581_, _42195_);
  or (_04204_, _03601_, _42154_);
  and (_04205_, _04204_, _04203_);
  or (_04206_, _03626_, _42072_);
  or (_04207_, _03606_, _41990_);
  and (_04208_, _04207_, _04206_);
  and (_04209_, _04208_, _04205_);
  and (_04210_, _04209_, _04202_);
  and (_04211_, _04210_, _04195_);
  nor (_04212_, _04211_, _03702_);
  not (_04213_, _04212_);
  nor (_04214_, _04211_, _03823_);
  nor (_04215_, _03812_, _03670_);
  not (_04216_, _03773_);
  nor (_04217_, _04211_, _04216_);
  or (_04218_, _04211_, _03751_);
  nor (_04219_, _04211_, _03759_);
  and (_04220_, _03799_, _03382_);
  nor (_04221_, _04220_, _03700_);
  not (_04222_, _03789_);
  and (_04223_, _03677_, _03845_);
  nor (_04224_, _04223_, _03791_);
  and (_04225_, _04224_, _04222_);
  and (_04226_, _04225_, _04221_);
  nor (_04227_, _04226_, _03449_);
  not (_04229_, _04227_);
  and (_04230_, _04223_, _03695_);
  nand (_04231_, _03349_, _03316_);
  nor (_04232_, _04231_, _03444_);
  nor (_04233_, _04232_, _04230_);
  and (_04234_, _03862_, _04108_);
  not (_04235_, _04234_);
  not (_04236_, _03454_);
  and (_04237_, _04223_, _04236_);
  nor (_04238_, _04237_, _03757_);
  and (_04239_, _04238_, _04235_);
  and (_04240_, _04239_, _04233_);
  and (_04241_, _04240_, _04229_);
  or (_04242_, _04241_, _04219_);
  nand (_04243_, _04242_, _03697_);
  nand (_04244_, _03698_, _04243_);
  and (_04245_, _03755_, _03674_);
  or (_04246_, _04245_, _03750_);
  and (_04247_, _04223_, _03689_);
  nor (_04248_, _04231_, _03447_);
  or (_04249_, _04248_, _04247_);
  nor (_04250_, _04249_, _04246_);
  nand (_04251_, _04250_, _04244_);
  nand (_04252_, _04251_, _04218_);
  and (_04253_, _04252_, _03692_);
  or (_04254_, _03693_, _04253_);
  and (_04255_, _04211_, _03690_);
  and (_04256_, _03799_, _03349_);
  nor (_04257_, _04256_, _03700_);
  and (_04258_, _04257_, _04222_);
  and (_04259_, _04258_, _04224_);
  nor (_04260_, _04259_, _03441_);
  nor (_04261_, _04260_, _04255_);
  and (_04262_, _04261_, _04254_);
  or (_04263_, _04262_, _04217_);
  nand (_04264_, _04263_, _03778_);
  nor (_04265_, _03778_, _03670_);
  nor (_04266_, _04265_, _03808_);
  nand (_04267_, _04266_, _04264_);
  and (_04268_, _04211_, _03808_);
  and (_04269_, _03853_, _03783_);
  and (_04270_, _04269_, _03349_);
  nor (_04271_, _04270_, _03813_);
  not (_04272_, _04271_);
  nor (_04273_, _04272_, _04268_);
  and (_04274_, _04273_, _04267_);
  or (_04275_, _04274_, _04215_);
  and (_04276_, _03789_, _03416_);
  nor (_04277_, _04223_, _04220_);
  nand (_04278_, _03677_, _03316_);
  and (_04279_, _04278_, _03414_);
  nand (_04280_, _04279_, _04277_);
  and (_04281_, _04280_, _03416_);
  nor (_04282_, _04281_, _04276_);
  and (_04283_, _04282_, _04275_);
  or (_04284_, _04283_, _04214_);
  and (_04285_, _04284_, _03680_);
  or (_04286_, _04285_, _03681_);
  and (_04287_, _03789_, _03410_);
  and (_04288_, _04223_, _03410_);
  nor (_04289_, _04288_, _04287_);
  not (_04290_, _04289_);
  not (_04291_, _03791_);
  and (_04292_, _04257_, _04291_);
  nor (_04293_, _04292_, _03411_);
  nor (_04294_, _04293_, _04290_);
  and (_04295_, _04294_, _04286_);
  and (_04296_, _03934_, _02136_);
  and (_04297_, _03907_, _02154_);
  nor (_04298_, _04297_, _04296_);
  and (_04299_, _03916_, _02149_);
  and (_04300_, _03939_, _02116_);
  nor (_04301_, _04300_, _04299_);
  and (_04302_, _04301_, _04298_);
  and (_04303_, _03936_, _02162_);
  and (_04304_, _03941_, _02127_);
  nor (_04305_, _04304_, _04303_);
  and (_04306_, _03928_, _02119_);
  and (_04307_, _03930_, _02132_);
  nor (_04308_, _04307_, _04306_);
  and (_04309_, _04308_, _04305_);
  and (_04310_, _04309_, _04302_);
  and (_04311_, _03925_, _02129_);
  and (_04312_, _03923_, _02147_);
  nor (_04313_, _04312_, _04311_);
  and (_04314_, _03913_, _02143_);
  and (_04315_, _03898_, _02141_);
  nor (_04316_, _04315_, _04314_);
  and (_04317_, _04316_, _04313_);
  and (_04318_, _03911_, _02165_);
  and (_04319_, _03918_, _02151_);
  nor (_04320_, _04319_, _04318_);
  and (_04321_, _03894_, _02138_);
  and (_04322_, _03903_, _02121_);
  nor (_04323_, _04322_, _04321_);
  and (_04324_, _04323_, _04320_);
  and (_04325_, _04324_, _04317_);
  and (_04326_, _04325_, _04310_);
  nor (_04327_, _04326_, _03415_);
  or (_04328_, _04327_, _04295_);
  and (_04330_, _03746_, _03670_);
  and (_04331_, _04223_, _03482_);
  nor (_04332_, _04331_, _03745_);
  not (_04333_, _04332_);
  nor (_04334_, _04333_, _04330_);
  and (_04335_, _04334_, _04328_);
  not (_04336_, _03745_);
  nor (_04337_, _04336_, _03670_);
  or (_04338_, _04337_, _04335_);
  and (_04339_, _04223_, _03485_);
  not (_04340_, _04231_);
  and (_04341_, _04340_, _03485_);
  nor (_04342_, _04341_, _04339_);
  and (_04343_, _04342_, _04338_);
  not (_04344_, _04211_);
  nor (_04345_, _04344_, _03961_);
  not (_04346_, _03476_);
  nor (_04347_, _04256_, _03789_);
  and (_04348_, _04347_, _04224_);
  nor (_04349_, _04348_, _04346_);
  nor (_04350_, _04349_, _04345_);
  and (_04351_, _04350_, _04343_);
  nor (_04352_, _04344_, _03969_);
  not (_04353_, _03480_);
  not (_04354_, _04220_);
  nor (_04355_, _04223_, _03789_);
  and (_04356_, _04355_, _04354_);
  or (_04357_, _04356_, _04353_);
  and (_04358_, _03862_, _03480_);
  and (_04359_, _03791_, _03480_);
  nor (_04360_, _04359_, _04358_);
  and (_04361_, _04360_, _04357_);
  not (_04362_, _04361_);
  nor (_04363_, _04362_, _04352_);
  and (_04364_, _04363_, _04351_);
  nor (_04365_, _04344_, _03956_);
  and (_04366_, _03791_, _03473_);
  not (_04367_, _04366_);
  and (_04368_, _03862_, _03473_);
  nor (_04369_, _04368_, _03963_);
  and (_04370_, _04369_, _04367_);
  and (_04371_, _04223_, _03473_);
  not (_04372_, _04371_);
  and (_04373_, _04220_, _03473_);
  and (_04374_, _03789_, _03473_);
  nor (_04375_, _04374_, _04373_);
  and (_04376_, _04375_, _04372_);
  and (_04377_, _04376_, _04370_);
  not (_04378_, _04377_);
  nor (_04379_, _04378_, _04365_);
  and (_04380_, _04379_, _04364_);
  nor (_04381_, _04211_, _03964_);
  or (_04382_, _04381_, _04380_);
  and (_04383_, _03974_, _03674_);
  nor (_04384_, _04383_, _03831_);
  and (_04385_, _04384_, _04382_);
  not (_04386_, _03831_);
  nor (_04387_, _04386_, _03670_);
  or (_04388_, _04387_, _04385_);
  not (_04389_, _03393_);
  and (_04390_, _04277_, _04278_);
  nor (_04391_, _04390_, _04389_);
  and (_04392_, _03789_, _03393_);
  nor (_04393_, _04392_, _03709_);
  not (_04394_, _04393_);
  nor (_04395_, _04394_, _04391_);
  and (_04396_, _04395_, _04388_);
  nor (_04397_, _04211_, _04166_);
  or (_04398_, _04397_, _04396_);
  and (_04399_, _03707_, _03674_);
  nor (_04400_, _04399_, _03705_);
  and (_04401_, _04400_, _04398_);
  nor (_04402_, _03706_, _03670_);
  nor (_04403_, _04402_, _04401_);
  not (_04404_, _03254_);
  nor (_04405_, _04259_, _04404_);
  nor (_04406_, _04405_, _04403_);
  nor (_04407_, _04211_, _03704_);
  or (_04408_, _04407_, _04406_);
  and (_04409_, _04408_, _03385_);
  nor (_04410_, _04409_, _03671_);
  nor (_04411_, _04259_, _04079_);
  or (_04412_, _04411_, _04410_);
  nand (_04413_, _04412_, _04213_);
  or (_04414_, _04413_, _04180_);
  nor (_04415_, _03592_, _41805_);
  nor (_04416_, _03616_, _41723_);
  nor (_04417_, _04416_, _04415_);
  nor (_04418_, _03603_, _42133_);
  nor (_04419_, _03628_, _41928_);
  nor (_04420_, _04419_, _04418_);
  and (_04421_, _04420_, _04417_);
  nor (_04422_, _03597_, _41682_);
  nor (_04423_, _03633_, _41633_);
  nor (_04424_, _04423_, _04422_);
  nor (_04425_, _03619_, _41887_);
  nor (_04426_, _03614_, _41764_);
  nor (_04427_, _04426_, _04425_);
  and (_04428_, _04427_, _04424_);
  and (_04429_, _04428_, _04421_);
  nor (_04431_, _03626_, _42092_);
  nor (_04432_, _03585_, _42051_);
  nor (_04433_, _04432_, _04431_);
  nor (_04434_, _03581_, _42215_);
  nor (_04435_, _03601_, _42174_);
  nor (_04436_, _04435_, _04434_);
  and (_04437_, _04436_, _04433_);
  nor (_04438_, _03606_, _42010_);
  nor (_04439_, _03608_, _41969_);
  nor (_04440_, _04439_, _04438_);
  nor (_04441_, _03631_, _41846_);
  nor (_04442_, _03621_, _41585_);
  nor (_04443_, _04442_, _04441_);
  and (_04444_, _04443_, _04440_);
  and (_04445_, _04444_, _04437_);
  and (_04446_, _04445_, _04429_);
  nor (_04447_, _04446_, _03638_);
  and (_04448_, _04447_, _04042_);
  not (_04449_, _04448_);
  and (_04450_, _04447_, _03384_);
  not (_04451_, _04450_);
  nor (_04452_, _03619_, _41872_);
  nor (_04453_, _03633_, _41618_);
  nor (_04454_, _04453_, _04452_);
  nor (_04455_, _03608_, _41954_);
  nor (_04456_, _03597_, _41667_);
  nor (_04457_, _04456_, _04455_);
  and (_04458_, _04457_, _04454_);
  nor (_04459_, _03585_, _42036_);
  nor (_04460_, _03621_, _41570_);
  nor (_04461_, _04460_, _04459_);
  nor (_04462_, _03581_, _42200_);
  nor (_04463_, _03603_, _42118_);
  nor (_04464_, _04463_, _04462_);
  and (_04465_, _04464_, _04461_);
  and (_04466_, _04465_, _04458_);
  nor (_04467_, _03601_, _42159_);
  nor (_04468_, _03616_, _41708_);
  nor (_04469_, _04468_, _04467_);
  nor (_04470_, _03628_, _41913_);
  nor (_04471_, _03631_, _41831_);
  nor (_04472_, _04471_, _04470_);
  and (_04473_, _04472_, _04469_);
  nor (_04474_, _03606_, _41995_);
  nor (_04475_, _03614_, _41749_);
  nor (_04476_, _04475_, _04474_);
  nor (_04477_, _03626_, _42077_);
  nor (_04478_, _03592_, _41790_);
  nor (_04479_, _04478_, _04477_);
  and (_04480_, _04479_, _04476_);
  and (_04481_, _04480_, _04473_);
  and (_04482_, _04481_, _04466_);
  nor (_04483_, _04482_, _04174_);
  not (_04484_, _04483_);
  and (_04485_, _03903_, _02216_);
  and (_04486_, _03930_, _02202_);
  nor (_04487_, _04486_, _04485_);
  and (_04488_, _03934_, _02196_);
  and (_04489_, _03898_, _02198_);
  nor (_04490_, _04489_, _04488_);
  and (_04491_, _04490_, _04487_);
  and (_04492_, _03911_, _02177_);
  and (_04493_, _03913_, _02193_);
  nor (_04494_, _04493_, _04492_);
  and (_04495_, _03916_, _02191_);
  and (_04496_, _03936_, _02214_);
  nor (_04497_, _04496_, _04495_);
  and (_04498_, _04497_, _04494_);
  and (_04499_, _04498_, _04491_);
  and (_04500_, _03939_, _02172_);
  and (_04501_, _03941_, _02185_);
  nor (_04502_, _04501_, _04500_);
  and (_04503_, _03928_, _02175_);
  and (_04504_, _03923_, _02183_);
  nor (_04505_, _04504_, _04503_);
  and (_04506_, _04505_, _04502_);
  and (_04507_, _03894_, _02204_);
  and (_04508_, _03918_, _02206_);
  nor (_04509_, _04508_, _04507_);
  and (_04510_, _03925_, _02187_);
  and (_04511_, _03907_, _02208_);
  nor (_04512_, _04511_, _04510_);
  and (_04513_, _04512_, _04509_);
  and (_04514_, _04513_, _04506_);
  and (_04515_, _04514_, _04499_);
  nor (_04516_, _04515_, _03415_);
  nor (_04517_, _03867_, _03803_);
  nor (_04518_, _03480_, _03695_);
  and (_04519_, _04518_, _04389_);
  nor (_04520_, _04519_, _04517_);
  not (_04521_, _04520_);
  and (_04522_, _03803_, _03485_);
  not (_04523_, _04522_);
  and (_04524_, _03803_, _03473_);
  and (_04525_, _03867_, _03476_);
  nor (_04526_, _04525_, _04524_);
  and (_04527_, _04526_, _04523_);
  and (_04528_, _03449_, _03447_);
  nor (_04529_, _04528_, _04099_);
  or (_04530_, _03683_, _03254_);
  and (_04532_, _04530_, _03867_);
  nor (_04533_, _04532_, _04529_);
  and (_04534_, _04533_, _04527_);
  and (_04535_, _04534_, _04521_);
  not (_04536_, \oc8051_golden_model_1.SP [1]);
  not (_04537_, _03755_);
  and (_04538_, _04126_, _04537_);
  nor (_04539_, _04538_, _04536_);
  or (_04540_, _03485_, _03410_);
  or (_04541_, _04540_, _03398_);
  nor (_04542_, _03473_, _03416_);
  nand (_04543_, _04542_, _04528_);
  or (_04544_, _04543_, _04541_);
  and (_04545_, _04544_, _03867_);
  nor (_04546_, _04545_, _04539_);
  and (_04547_, _04546_, _04535_);
  and (_04548_, _04547_, _04104_);
  not (_04549_, _04548_);
  nor (_04550_, _04549_, _04516_);
  and (_04551_, _04550_, _04484_);
  and (_04552_, _04551_, _04451_);
  and (_04553_, _04552_, _04449_);
  not (_04554_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_04555_, _04412_, _04213_);
  or (_04556_, _04555_, _04554_);
  and (_04557_, _04556_, _04553_);
  nand (_04558_, _04557_, _04414_);
  not (_04559_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_04560_, _04555_, _04559_);
  not (_04561_, _04553_);
  not (_04562_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_04563_, _04413_, _04562_);
  and (_04564_, _04563_, _04561_);
  nand (_04565_, _04564_, _04560_);
  nand (_04566_, _04565_, _04558_);
  nand (_04567_, _04566_, _04179_);
  not (_04568_, _04179_);
  not (_04569_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_04570_, _04555_, _04569_);
  not (_04571_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_04572_, _04413_, _04571_);
  and (_04573_, _04572_, _04561_);
  nand (_04574_, _04573_, _04570_);
  not (_04575_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_04576_, _04413_, _04575_);
  not (_04577_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_04578_, _04555_, _04577_);
  and (_04579_, _04578_, _04553_);
  nand (_04580_, _04579_, _04576_);
  nand (_04581_, _04580_, _04574_);
  nand (_04582_, _04581_, _04568_);
  nand (_04583_, _04582_, _04567_);
  nand (_04584_, _04583_, _04002_);
  not (_04585_, _04002_);
  nand (_04586_, _04413_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_04587_, _04555_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_04588_, _04587_, _04561_);
  nand (_04589_, _04588_, _04586_);
  nand (_04590_, _04555_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_04591_, _04413_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_04592_, _04591_, _04553_);
  nand (_04593_, _04592_, _04590_);
  nand (_04594_, _04593_, _04589_);
  nand (_04595_, _04594_, _04179_);
  nand (_04596_, _04413_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_04597_, _04555_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_04598_, _04597_, _04561_);
  nand (_04599_, _04598_, _04596_);
  nand (_04600_, _04555_, \oc8051_golden_model_1.IRAM[12] [0]);
  nand (_04601_, _04413_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_04602_, _04601_, _04553_);
  nand (_04603_, _04602_, _04600_);
  nand (_04604_, _04603_, _04599_);
  nand (_04605_, _04604_, _04568_);
  nand (_04606_, _04605_, _04595_);
  nand (_04607_, _04606_, _04585_);
  and (_04608_, _04607_, _04584_);
  and (_04609_, _04608_, _03699_);
  nor (_04610_, _03846_, _03388_);
  and (_04611_, _04610_, _04355_);
  nor (_04612_, _04611_, _03454_);
  not (_04613_, _04612_);
  nor (_04614_, _04613_, _04609_);
  and (_04615_, _03850_, _04108_);
  not (_04616_, _04615_);
  nor (_04617_, _04616_, _03638_);
  and (_04618_, _04211_, _04617_);
  or (_04619_, _04618_, _04614_);
  and (_04620_, _04111_, \oc8051_golden_model_1.SP [0]);
  nor (_04621_, _04620_, _04232_);
  not (_04622_, _04621_);
  nor (_04623_, _04622_, _04619_);
  and (_04624_, _03853_, _03695_);
  not (_04625_, _04624_);
  nor (_04626_, _04625_, _04608_);
  not (_04627_, _04626_);
  and (_04628_, _04627_, _04623_);
  nor (_04629_, _03697_, _03638_);
  not (_04630_, _03757_);
  nor (_04631_, _04630_, _03638_);
  and (_04633_, _04631_, _04211_);
  nor (_04634_, _04633_, _04629_);
  and (_04635_, _04634_, _04628_);
  not (_04636_, _04635_);
  and (_04637_, _04636_, _03698_);
  nor (_04638_, _03445_, _03674_);
  nor (_04639_, _04638_, _04637_);
  nor (_04640_, _04537_, _03638_);
  and (_04641_, _04640_, _04211_);
  nor (_04642_, _04641_, _04248_);
  and (_04643_, _04642_, _04639_);
  nor (_04644_, _03751_, _03638_);
  and (_04645_, _03853_, _03689_);
  not (_04646_, _04645_);
  nor (_04647_, _04646_, _04608_);
  nor (_04648_, _04647_, _04644_);
  and (_04649_, _04648_, _04643_);
  and (_04650_, _04644_, _04344_);
  nor (_04651_, _04650_, _04649_);
  nor (_04652_, _04651_, _03694_);
  nor (_04653_, _04652_, _03693_);
  or (_04654_, _04653_, _03690_);
  nand (_04655_, _03690_, _03674_);
  nand (_04656_, _04655_, _04654_);
  and (_04657_, _04656_, _03688_);
  nor (_04658_, _04657_, _03686_);
  nor (_04659_, _04231_, _03452_);
  or (_04660_, _04659_, _04658_);
  nor (_04661_, _04660_, _03682_);
  nor (_04662_, _03680_, _03638_);
  not (_04663_, _04269_);
  nor (_04664_, _04608_, _04663_);
  nor (_04665_, _04664_, _04662_);
  and (_04666_, _04665_, _04661_);
  nor (_04667_, _04666_, _03681_);
  nor (_04668_, _04667_, _03676_);
  nor (_04669_, _03418_, \oc8051_golden_model_1.SP [0]);
  nor (_04670_, _04669_, _04668_);
  or (_04671_, _04110_, _03803_);
  nor (_04672_, _03638_, _03411_);
  and (_04673_, _04672_, _04671_);
  nor (_04674_, _04220_, _03785_);
  not (_04675_, _04674_);
  and (_04676_, _04675_, _04672_);
  nor (_04677_, _04676_, _04673_);
  and (_04678_, _03853_, _03410_);
  not (_04679_, _04678_);
  nor (_04680_, _04679_, _03638_);
  and (_04681_, _04672_, _03700_);
  nor (_04682_, _04681_, _04680_);
  and (_04683_, _04682_, _04677_);
  nor (_04684_, _04683_, _04344_);
  and (_04685_, _04340_, _03482_);
  nor (_04686_, _04685_, _04684_);
  not (_04687_, _04686_);
  nor (_04688_, _04687_, _04670_);
  and (_04689_, _03853_, _03482_);
  not (_04690_, _04689_);
  nor (_04691_, _04690_, _04608_);
  not (_04692_, _04691_);
  and (_04693_, _04692_, _04688_);
  not (_04694_, _03839_);
  nor (_04695_, _04694_, _03638_);
  and (_04696_, _04695_, _04211_);
  nor (_04697_, _04696_, _03483_);
  and (_04698_, _04697_, _04693_);
  and (_04699_, _03483_, _03674_);
  nor (_04700_, _04699_, _04698_);
  not (_04701_, _03959_);
  nor (_04702_, _04701_, _03638_);
  not (_04703_, _03838_);
  nor (_04704_, _04703_, _03638_);
  nor (_04705_, _04704_, _04702_);
  not (_04706_, _03967_);
  nor (_04707_, _04706_, _03638_);
  not (_04708_, _03866_);
  nor (_04709_, _04708_, _03638_);
  nor (_04710_, _04709_, _04707_);
  and (_04711_, _04710_, _04705_);
  nor (_04712_, _04711_, _04344_);
  nor (_04713_, _04712_, _03477_);
  not (_04714_, _04713_);
  nor (_04715_, _04714_, _04700_);
  and (_04716_, _03477_, _03674_);
  nor (_04717_, _04716_, _04715_);
  nor (_04718_, _03955_, _03638_);
  and (_04719_, _04718_, _04211_);
  nor (_04720_, _04719_, _03474_);
  not (_04721_, _04720_);
  nor (_04722_, _04721_, _04717_);
  nor (_04723_, _04722_, _03675_);
  and (_04724_, _04340_, _03254_);
  nor (_04725_, _04724_, _04723_);
  nor (_04726_, _03704_, _03638_);
  and (_04727_, _03853_, _03254_);
  not (_04728_, _04727_);
  nor (_04729_, _04728_, _04608_);
  nor (_04730_, _04729_, _04726_);
  and (_04731_, _04730_, _04725_);
  and (_04732_, _04726_, _04344_);
  nor (_04734_, _04732_, _04731_);
  nor (_04735_, _03833_, _03400_);
  nor (_04736_, _04735_, _03674_);
  nor (_04737_, _04736_, _04734_);
  and (_04738_, _04737_, _03673_);
  nor (_04739_, _04738_, _03671_);
  and (_04740_, _04340_, _03398_);
  nor (_04741_, _04740_, _04739_);
  nor (_04742_, _03702_, _03638_);
  and (_04743_, _03853_, _03398_);
  not (_04744_, _04743_);
  nor (_04745_, _04744_, _04608_);
  nor (_04746_, _04745_, _04742_);
  and (_04747_, _04746_, _04741_);
  and (_04748_, _04742_, _04344_);
  nor (_04749_, _04748_, _04747_);
  not (_04750_, _04482_);
  and (_04751_, _04742_, _04750_);
  and (_04752_, _04536_, \oc8051_golden_model_1.SP [0]);
  and (_04753_, \oc8051_golden_model_1.SP [1], _03674_);
  nor (_04754_, _04753_, _04752_);
  not (_04755_, _04754_);
  and (_04756_, _04755_, _03474_);
  and (_04757_, _04695_, _04750_);
  and (_04758_, _04447_, _03679_);
  not (_04759_, _03690_);
  and (_04760_, _04631_, _04750_);
  not (_04761_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_04762_, _04413_, _04761_);
  not (_04763_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_04764_, _04555_, _04763_);
  and (_04765_, _04764_, _04553_);
  nand (_04766_, _04765_, _04762_);
  not (_04767_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_04768_, _04555_, _04767_);
  not (_04769_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_04770_, _04413_, _04769_);
  and (_04771_, _04770_, _04561_);
  nand (_04772_, _04771_, _04768_);
  nand (_04773_, _04772_, _04766_);
  nand (_04774_, _04773_, _04179_);
  not (_04775_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_04776_, _04555_, _04775_);
  not (_04777_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_04778_, _04413_, _04777_);
  and (_04779_, _04778_, _04561_);
  nand (_04780_, _04779_, _04776_);
  not (_04781_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_04782_, _04413_, _04781_);
  not (_04783_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_04784_, _04555_, _04783_);
  and (_04785_, _04784_, _04553_);
  nand (_04786_, _04785_, _04782_);
  nand (_04787_, _04786_, _04780_);
  nand (_04788_, _04787_, _04568_);
  nand (_04789_, _04788_, _04774_);
  nand (_04790_, _04789_, _04002_);
  nand (_04791_, _04413_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_04792_, _04555_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_04793_, _04792_, _04561_);
  nand (_04794_, _04793_, _04791_);
  nand (_04795_, _04555_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_04796_, _04413_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_04797_, _04796_, _04553_);
  nand (_04798_, _04797_, _04795_);
  nand (_04799_, _04798_, _04794_);
  nand (_04800_, _04799_, _04179_);
  nand (_04801_, _04413_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_04802_, _04555_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_04803_, _04802_, _04561_);
  nand (_04804_, _04803_, _04801_);
  nand (_04805_, _04555_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_04806_, _04413_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_04807_, _04806_, _04553_);
  nand (_04808_, _04807_, _04805_);
  nand (_04809_, _04808_, _04804_);
  nand (_04810_, _04809_, _04568_);
  nand (_04811_, _04810_, _04800_);
  nand (_04812_, _04811_, _04585_);
  and (_04813_, _04812_, _04790_);
  nor (_04814_, _04624_, _03699_);
  or (_04815_, _04814_, _04813_);
  not (_04816_, _04631_);
  and (_04817_, _04754_, _04111_);
  nor (_04818_, _03444_, _03380_);
  and (_04819_, _04818_, _03316_);
  nor (_04820_, _04819_, _04817_);
  and (_04821_, _04750_, _04617_);
  or (_04822_, _04821_, _04111_);
  and (_04823_, _03853_, _04236_);
  nor (_04824_, _04823_, _04617_);
  or (_04825_, _04824_, _04822_);
  and (_04826_, _04825_, _04820_);
  and (_04827_, _04826_, _04816_);
  and (_04828_, _04827_, _04815_);
  nor (_04829_, _04828_, _04760_);
  and (_04830_, _04446_, _04629_);
  or (_04831_, _04830_, _04829_);
  nor (_04832_, _04755_, _03445_);
  nor (_04833_, _04832_, _04640_);
  not (_04834_, _04833_);
  nor (_04835_, _04834_, _04831_);
  and (_04836_, _04640_, _04750_);
  nor (_04837_, _04836_, _04835_);
  not (_04838_, _03316_);
  nor (_04839_, _03447_, _04838_);
  and (_04840_, _04839_, _03381_);
  nor (_04841_, _04840_, _04837_);
  nand (_04842_, _04812_, _04790_);
  and (_04843_, _04842_, _04645_);
  nor (_04844_, _04843_, _04644_);
  and (_04845_, _04844_, _04841_);
  and (_04846_, _04644_, _04750_);
  nor (_04847_, _04846_, _04845_);
  and (_04848_, _04446_, _03694_);
  nor (_04849_, _04848_, _04847_);
  and (_04850_, _04849_, _04759_);
  and (_04851_, _04755_, _03690_);
  nor (_04852_, _04851_, _04850_);
  and (_04853_, _03687_, _04446_);
  nor (_04854_, _04853_, _04852_);
  nor (_04855_, _04755_, _03442_);
  nor (_04856_, _03452_, _03380_);
  and (_04857_, _04856_, _03316_);
  nor (_04858_, _04857_, _04855_);
  and (_04859_, _04858_, _04854_);
  and (_04860_, _04842_, _04269_);
  nor (_04861_, _04860_, _04662_);
  and (_04862_, _04861_, _04859_);
  nor (_04863_, _04862_, _04758_);
  nor (_04864_, _04863_, _03676_);
  nor (_04865_, _04754_, _03418_);
  nor (_04866_, _04865_, _04864_);
  nor (_04867_, _04683_, _04750_);
  and (_04868_, _03482_, _03381_);
  and (_04869_, _04868_, _03316_);
  nor (_04870_, _04869_, _04867_);
  not (_04871_, _04870_);
  nor (_04872_, _04871_, _04866_);
  nor (_04873_, _04813_, _04690_);
  nor (_04874_, _04873_, _04695_);
  and (_04875_, _04874_, _04872_);
  nor (_04876_, _04875_, _04757_);
  nor (_04877_, _04876_, _03483_);
  and (_04878_, _04755_, _03483_);
  nor (_04879_, _04878_, _04877_);
  nor (_04880_, _04711_, _04750_);
  nor (_04881_, _04880_, _03477_);
  not (_04882_, _04881_);
  nor (_04883_, _04882_, _04879_);
  and (_04884_, _04755_, _03477_);
  nor (_04885_, _04884_, _04883_);
  and (_04886_, _04718_, _04482_);
  nor (_04887_, _04886_, _03474_);
  not (_04888_, _04887_);
  nor (_04889_, _04888_, _04885_);
  nor (_04890_, _04889_, _04756_);
  and (_04891_, _03858_, _03254_);
  nor (_04892_, _04891_, _04120_);
  not (_04893_, _04892_);
  nor (_04894_, _04893_, _04890_);
  and (_04895_, _04842_, _04727_);
  nor (_04896_, _04895_, _04726_);
  and (_04897_, _04896_, _04894_);
  and (_04898_, _04726_, _04750_);
  nor (_04899_, _04898_, _04897_);
  nor (_04900_, _04755_, _04735_);
  nor (_04901_, _04900_, _04899_);
  and (_04902_, _04901_, _03673_);
  nor (_04903_, _04902_, _04450_);
  and (_04904_, _03800_, _03398_);
  and (_04905_, _03789_, _03398_);
  and (_04906_, _03786_, _03398_);
  or (_04907_, _04906_, _04905_);
  nor (_04908_, _04907_, _04904_);
  not (_04909_, _04908_);
  nor (_04910_, _04909_, _04903_);
  and (_04911_, _04842_, _04743_);
  nor (_04912_, _04911_, _04742_);
  and (_04913_, _04912_, _04910_);
  nor (_04914_, _04913_, _04751_);
  not (_04915_, _00000_);
  not (_04916_, _04676_);
  nor (_04917_, _04681_, _04673_);
  and (_04918_, _04917_, _04916_);
  nor (_04919_, _04640_, _04631_);
  nor (_04920_, _03687_, _04617_);
  and (_04921_, _04920_, _04919_);
  not (_04922_, _04742_);
  and (_04923_, _03789_, _03689_);
  not (_04924_, _04923_);
  not (_04925_, _04906_);
  and (_04926_, _03785_, _03254_);
  nor (_04927_, _04926_, _04120_);
  and (_04928_, _04927_, _04925_);
  and (_04929_, _04928_, _04924_);
  nor (_04930_, _04624_, _04269_);
  nor (_04931_, _04114_, _03690_);
  and (_04932_, _04931_, _04930_);
  not (_04933_, _03445_);
  nor (_04934_, _03483_, _04933_);
  nor (_04935_, _04727_, _04689_);
  and (_04936_, _04935_, _04934_);
  and (_04937_, _04936_, _04932_);
  and (_04938_, _04937_, _04929_);
  and (_04939_, _03858_, _04236_);
  nor (_04940_, _04939_, _04823_);
  nand (_04941_, _04610_, _03414_);
  and (_04942_, _04941_, _04236_);
  not (_04943_, _04942_);
  and (_04944_, _04943_, _04940_);
  and (_04945_, _04944_, _03795_);
  and (_04946_, _04945_, _04938_);
  nor (_04947_, _04743_, _04905_);
  not (_04948_, _04111_);
  and (_04949_, _04948_, _03478_);
  and (_04950_, _04949_, _03806_);
  and (_04951_, _04950_, _04947_);
  and (_04952_, _03867_, _03695_);
  and (_04953_, _03867_, _03482_);
  nor (_04954_, _04953_, _04952_);
  and (_04955_, _04100_, _03803_);
  not (_04956_, _03382_);
  and (_04957_, _03785_, _04956_);
  and (_04958_, _04957_, _03689_);
  nor (_04959_, _04958_, _04955_);
  and (_04960_, _04959_, _04954_);
  and (_04961_, _03858_, _03482_);
  nor (_04962_, _04961_, _04645_);
  and (_04963_, _03858_, _03695_);
  and (_04964_, _03850_, _03482_);
  nor (_04965_, _04964_, _04963_);
  and (_04966_, _04965_, _04962_);
  and (_04967_, _04966_, _04960_);
  and (_04968_, _03442_, _03418_);
  and (_04969_, _04968_, _04735_);
  and (_04970_, _03799_, _03420_);
  and (_04971_, _04970_, _03482_);
  not (_04972_, _04971_);
  and (_04973_, _03867_, _03398_);
  nor (_04974_, _04973_, _04904_);
  and (_04975_, _04974_, _04972_);
  and (_04976_, _04975_, _04969_);
  and (_04977_, _04976_, _04967_);
  and (_04978_, _04977_, _04951_);
  and (_04979_, _04978_, _04946_);
  and (_04980_, _04979_, _04922_);
  nor (_04981_, _04695_, _04644_);
  and (_04982_, _04981_, _04980_);
  and (_04983_, _04982_, _04921_);
  nor (_04984_, _03703_, _03384_);
  and (_04985_, _04984_, _04037_);
  nor (_04986_, _04985_, _03638_);
  not (_04987_, _04986_);
  nor (_04988_, _04718_, _04680_);
  and (_04989_, _04988_, _04987_);
  and (_04990_, _04989_, _04711_);
  and (_04991_, _04990_, _04983_);
  and (_04992_, _04991_, _04918_);
  nor (_04993_, _04992_, _04915_);
  not (_04994_, _04993_);
  nor (_04995_, _04994_, _04914_);
  not (_04996_, _04995_);
  nor (_04997_, _04996_, _04749_);
  not (_04998_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_04999_, _04413_, _04998_);
  not (_05000_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_05001_, _04555_, _05000_);
  and (_05002_, _05001_, _04553_);
  nand (_05003_, _05002_, _04999_);
  not (_05004_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_05005_, _04555_, _05004_);
  not (_05006_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_05007_, _04413_, _05006_);
  and (_05008_, _05007_, _04561_);
  nand (_05009_, _05008_, _05005_);
  nand (_05010_, _05009_, _05003_);
  nand (_05011_, _05010_, _04179_);
  not (_05012_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_05013_, _04555_, _05012_);
  not (_05014_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_05015_, _04413_, _05014_);
  and (_05016_, _05015_, _04561_);
  nand (_05017_, _05016_, _05013_);
  not (_05018_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_05019_, _04413_, _05018_);
  not (_05020_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_05021_, _04555_, _05020_);
  and (_05022_, _05021_, _04553_);
  nand (_05023_, _05022_, _05019_);
  nand (_05024_, _05023_, _05017_);
  nand (_05025_, _05024_, _04568_);
  nand (_05026_, _05025_, _05011_);
  nand (_05027_, _05026_, _04002_);
  nand (_05028_, _04413_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_05029_, _04555_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_05030_, _05029_, _04561_);
  nand (_05031_, _05030_, _05028_);
  nand (_05032_, _04555_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_05033_, _04413_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_05034_, _05033_, _04553_);
  nand (_05035_, _05034_, _05032_);
  nand (_05036_, _05035_, _05031_);
  nand (_05037_, _05036_, _04179_);
  nand (_05038_, _04413_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_05039_, _04555_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_05040_, _05039_, _04561_);
  nand (_05041_, _05040_, _05038_);
  nand (_05042_, _04555_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_05043_, _04413_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_05044_, _05043_, _04553_);
  nand (_05045_, _05044_, _05042_);
  nand (_05046_, _05045_, _05041_);
  nand (_05047_, _05046_, _04568_);
  nand (_05048_, _05047_, _05037_);
  nand (_05049_, _05048_, _04585_);
  nand (_05050_, _05049_, _05027_);
  and (_05051_, _05050_, _04743_);
  and (_05052_, _05050_, _04689_);
  and (_05053_, _04629_, _03740_);
  and (_05054_, _05050_, _04624_);
  and (_05055_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_05056_, _05055_, \oc8051_golden_model_1.SP [2]);
  nor (_05057_, _05056_, \oc8051_golden_model_1.SP [3]);
  and (_05058_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_05059_, _05058_, \oc8051_golden_model_1.SP [3]);
  and (_05060_, _05059_, \oc8051_golden_model_1.SP [0]);
  nor (_05061_, _05060_, _05057_);
  and (_05062_, _05061_, _04111_);
  and (_05063_, _05050_, _03699_);
  not (_05064_, \oc8051_golden_model_1.PSW [3]);
  and (_05065_, _03455_, _05064_);
  nor (_05066_, _05065_, _05063_);
  nor (_05067_, _05066_, _04617_);
  and (_05068_, _04617_, _03669_);
  nor (_05069_, _05068_, _04111_);
  not (_05070_, _05069_);
  nor (_05071_, _05070_, _05067_);
  or (_05072_, _05071_, _04624_);
  nor (_05073_, _05072_, _05062_);
  or (_05074_, _05073_, _04631_);
  nor (_05075_, _05074_, _05054_);
  and (_05076_, _04631_, _03742_);
  or (_05077_, _05076_, _04629_);
  nor (_05078_, _05077_, _05075_);
  nor (_05079_, _05078_, _05053_);
  nor (_05080_, _05079_, _04933_);
  nor (_05081_, _05061_, _03445_);
  nor (_05082_, _05081_, _04640_);
  not (_05083_, _05082_);
  nor (_05084_, _05083_, _05080_);
  and (_05085_, _04640_, _03742_);
  nor (_05086_, _05085_, _04645_);
  not (_05087_, _05086_);
  nor (_05088_, _05087_, _05084_);
  and (_05089_, _05050_, _04645_);
  nor (_05090_, _05089_, _04644_);
  not (_05091_, _05090_);
  nor (_05092_, _05091_, _05088_);
  and (_05093_, _04644_, _03742_);
  or (_05094_, _05093_, _03694_);
  nor (_05095_, _05094_, _05092_);
  and (_05096_, _03740_, _03694_);
  nor (_05097_, _05096_, _05095_);
  and (_05098_, _05097_, _04759_);
  and (_05099_, _05061_, _03690_);
  nor (_05100_, _05099_, _05098_);
  nor (_05101_, _05100_, _03687_);
  nor (_05102_, _03688_, _03744_);
  or (_05103_, _05102_, _05101_);
  and (_05104_, _05103_, _03442_);
  not (_05105_, _03442_);
  nor (_05106_, _04269_, _05105_);
  nor (_05107_, _05061_, _04269_);
  nor (_05108_, _05107_, _05106_);
  nor (_05109_, _05108_, _05104_);
  and (_05110_, _05050_, _04269_);
  nor (_05111_, _05110_, _04662_);
  not (_05112_, _05111_);
  nor (_05113_, _05112_, _05109_);
  not (_05114_, _04662_);
  nor (_05115_, _05114_, _03744_);
  nor (_05116_, _05115_, _05113_);
  nor (_05117_, _05116_, _03676_);
  and (_05118_, _05061_, _03676_);
  not (_05119_, _05118_);
  and (_05120_, _05119_, _04683_);
  not (_05121_, _05120_);
  nor (_05122_, _05121_, _05117_);
  nor (_05123_, _04683_, _03742_);
  nor (_05124_, _05123_, _05122_);
  nor (_05125_, _05124_, _04689_);
  or (_05126_, _05125_, _04695_);
  nor (_05127_, _05126_, _05052_);
  and (_05128_, _04695_, _03742_);
  nor (_05129_, _05128_, _05127_);
  nor (_05130_, _05129_, _03483_);
  and (_05131_, _05061_, _03483_);
  not (_05132_, _05131_);
  and (_05133_, _05132_, _04711_);
  not (_05134_, _05133_);
  nor (_05135_, _05134_, _05130_);
  nor (_05136_, _04711_, _03742_);
  nor (_05137_, _05136_, _03477_);
  not (_05138_, _05137_);
  nor (_05139_, _05138_, _05135_);
  and (_05140_, _05061_, _03477_);
  nor (_05141_, _05140_, _04718_);
  not (_05142_, _05141_);
  nor (_05143_, _05142_, _05139_);
  and (_05144_, _04718_, _03669_);
  nor (_05145_, _05144_, _03474_);
  not (_05146_, _05145_);
  nor (_05147_, _05146_, _05143_);
  and (_05148_, _05061_, _03474_);
  nor (_05149_, _05148_, _04727_);
  not (_05150_, _05149_);
  nor (_05151_, _05150_, _05147_);
  and (_05152_, _05050_, _04727_);
  nor (_05153_, _05152_, _04726_);
  not (_05154_, _05153_);
  nor (_05155_, _05154_, _05151_);
  not (_05156_, _04735_);
  and (_05157_, _04726_, _03742_);
  nor (_05158_, _05157_, _05156_);
  not (_05159_, _05158_);
  nor (_05160_, _05159_, _05155_);
  nor (_05161_, _05061_, _04735_);
  nor (_05162_, _05161_, _03672_);
  not (_05163_, _05162_);
  nor (_05164_, _05163_, _05160_);
  not (_05165_, _03740_);
  and (_05166_, _03672_, _05165_);
  nor (_05167_, _05166_, _04743_);
  not (_05168_, _05167_);
  nor (_05169_, _05168_, _05164_);
  or (_05170_, _05169_, _04742_);
  nor (_05171_, _05170_, _05051_);
  and (_05172_, _04742_, _03742_);
  nor (_05173_, _05172_, _05171_);
  not (_05174_, _04165_);
  and (_05175_, _04742_, _05174_);
  nor (_05176_, _05055_, \oc8051_golden_model_1.SP [2]);
  nor (_05177_, _05176_, _05056_);
  and (_05178_, _05177_, _03474_);
  and (_05179_, _04695_, _05174_);
  and (_05180_, _04035_, _03679_);
  nor (_05181_, _05177_, _03442_);
  or (_05182_, _05181_, _03798_);
  nor (_05183_, _05182_, _03794_);
  not (_05184_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_05185_, _04413_, _05184_);
  not (_05186_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_05187_, _04555_, _05186_);
  and (_05188_, _05187_, _04553_);
  nand (_05189_, _05188_, _05185_);
  not (_05190_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_05191_, _04555_, _05190_);
  not (_05192_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_05193_, _04413_, _05192_);
  and (_05194_, _05193_, _04561_);
  nand (_05195_, _05194_, _05191_);
  nand (_05196_, _05195_, _05189_);
  nand (_05197_, _05196_, _04179_);
  not (_05198_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_05199_, _04555_, _05198_);
  not (_05200_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_05201_, _04413_, _05200_);
  and (_05202_, _05201_, _04561_);
  nand (_05203_, _05202_, _05199_);
  not (_05204_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_05205_, _04413_, _05204_);
  not (_05206_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_05207_, _04555_, _05206_);
  and (_05208_, _05207_, _04553_);
  nand (_05209_, _05208_, _05205_);
  nand (_05210_, _05209_, _05203_);
  nand (_05211_, _05210_, _04568_);
  nand (_05212_, _05211_, _05197_);
  nand (_05213_, _05212_, _04002_);
  nand (_05214_, _04413_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_05215_, _04555_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_05216_, _05215_, _04561_);
  nand (_05217_, _05216_, _05214_);
  nand (_05218_, _04555_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_05219_, _04413_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_05220_, _05219_, _04553_);
  nand (_05221_, _05220_, _05218_);
  nand (_05222_, _05221_, _05217_);
  nand (_05223_, _05222_, _04179_);
  nand (_05224_, _04413_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_05225_, _04555_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_05226_, _05225_, _04561_);
  nand (_05227_, _05226_, _05224_);
  nand (_05228_, _04555_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_05229_, _04413_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_05230_, _05229_, _04553_);
  nand (_05231_, _05230_, _05228_);
  nand (_05232_, _05231_, _05227_);
  nand (_05233_, _05232_, _04568_);
  nand (_05234_, _05233_, _05223_);
  nand (_05235_, _05234_, _04585_);
  nand (_05236_, _05235_, _05213_);
  nor (_05237_, _05236_, _03455_);
  nor (_05238_, _05237_, _04943_);
  and (_05239_, _04165_, _04617_);
  nor (_05240_, _05239_, _05238_);
  not (_05241_, _05177_);
  and (_05242_, _05241_, _04111_);
  and (_05243_, _03785_, _03695_);
  nor (_05244_, _05243_, _05242_);
  and (_05245_, _05244_, _05240_);
  and (_05246_, _05236_, _04624_);
  nor (_05247_, _05246_, _04631_);
  and (_05248_, _05247_, _05245_);
  and (_05249_, _04631_, _05174_);
  nor (_05250_, _05249_, _05248_);
  and (_05251_, _04629_, _04034_);
  nor (_05252_, _05251_, _05250_);
  or (_05253_, _05177_, _03445_);
  nand (_05254_, _05253_, _05252_);
  and (_05255_, _03785_, _03689_);
  and (_05256_, _04640_, _04165_);
  nor (_05257_, _05256_, _05255_);
  not (_05258_, _05257_);
  nor (_05259_, _05258_, _05254_);
  and (_05260_, _05236_, _04645_);
  nor (_05261_, _05260_, _04644_);
  and (_05262_, _05261_, _05259_);
  and (_05263_, _04644_, _05174_);
  nor (_05264_, _05263_, _05262_);
  and (_05265_, _04034_, _03694_);
  nor (_05266_, _05265_, _05264_);
  and (_05267_, _05266_, _04759_);
  and (_05268_, _05177_, _03690_);
  nor (_05269_, _05268_, _05267_);
  and (_05270_, _03687_, _04034_);
  nor (_05271_, _05270_, _05269_);
  and (_05272_, _05271_, _05183_);
  and (_05273_, _05236_, _04269_);
  nor (_05274_, _05273_, _04662_);
  and (_05275_, _05274_, _05272_);
  nor (_05276_, _05275_, _05180_);
  nor (_05277_, _05276_, _03676_);
  nor (_05278_, _05241_, _03418_);
  nor (_05279_, _05278_, _05277_);
  nor (_05280_, _04683_, _05174_);
  and (_05281_, _03785_, _03482_);
  nor (_05282_, _05281_, _05280_);
  not (_05283_, _05282_);
  nor (_05284_, _05283_, _05279_);
  and (_05285_, _05236_, _04689_);
  nor (_05286_, _05285_, _04695_);
  and (_05287_, _05286_, _05284_);
  nor (_05288_, _05287_, _05179_);
  nor (_05289_, _05288_, _03483_);
  and (_05290_, _05177_, _03483_);
  nor (_05291_, _05290_, _05289_);
  nor (_05292_, _04711_, _05174_);
  nor (_05293_, _05292_, _03477_);
  not (_05294_, _05293_);
  nor (_05295_, _05294_, _05291_);
  and (_05296_, _05177_, _03477_);
  nor (_05297_, _05296_, _05295_);
  and (_05298_, _04718_, _04165_);
  nor (_05299_, _05298_, _03474_);
  not (_05300_, _05299_);
  nor (_05301_, _05300_, _05297_);
  nor (_05302_, _05301_, _05178_);
  nor (_05303_, _05302_, _04926_);
  and (_05304_, _05236_, _04727_);
  nor (_05305_, _05304_, _04726_);
  and (_05306_, _05305_, _05303_);
  and (_05307_, _04726_, _05174_);
  nor (_05308_, _05307_, _05306_);
  nor (_05309_, _05177_, _04735_);
  nor (_05310_, _05309_, _05308_);
  and (_05311_, _05310_, _03673_);
  nor (_05312_, _05311_, _04045_);
  and (_05313_, _03785_, _03398_);
  nor (_05314_, _05313_, _05312_);
  and (_05315_, _05236_, _04743_);
  nor (_05316_, _05315_, _04742_);
  and (_05317_, _05316_, _05314_);
  nor (_05318_, _05317_, _05175_);
  nor (_05319_, _05318_, _04994_);
  not (_05320_, _05319_);
  nor (_05321_, _05320_, _05173_);
  and (_05322_, _05321_, _04997_);
  or (_05323_, _05322_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_05324_, _05058_, _03674_);
  nor (_05325_, _05177_, _04753_);
  nor (_05326_, _05325_, _05324_);
  and (_05327_, _05059_, _03674_);
  nor (_05328_, _05324_, _05061_);
  nor (_05329_, _05328_, _05327_);
  and (_05330_, _43759_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_05331_, _05330_);
  and (_05332_, _04969_, _04934_);
  and (_05333_, _05332_, _04949_);
  nor (_05334_, _05333_, _05331_);
  and (_05335_, _05334_, _05329_);
  and (_05336_, _05335_, _05326_);
  and (_05337_, _05336_, _04752_);
  not (_05338_, _05337_);
  and (_05339_, _05338_, _05323_);
  not (_05340_, _05322_);
  and (_05341_, _04482_, _04211_);
  and (_05342_, _04165_, _03742_);
  and (_05343_, _05342_, _05341_);
  and (_05344_, _03740_, _03638_);
  nor (_05345_, _04446_, _04034_);
  and (_05346_, _05345_, _05344_);
  and (_05347_, _05346_, _05343_);
  and (_05348_, _05347_, \oc8051_golden_model_1.IP [7]);
  and (_05349_, _04165_, _03669_);
  and (_05350_, _05349_, _05341_);
  not (_05351_, _03638_);
  nor (_05352_, _03740_, _05351_);
  and (_05353_, _05352_, _05345_);
  and (_05354_, _05353_, _05350_);
  and (_05355_, _05354_, \oc8051_golden_model_1.B [7]);
  nor (_05356_, _05355_, _05348_);
  not (_05357_, _04446_);
  and (_05358_, _05357_, _04034_);
  and (_05359_, _05358_, _05352_);
  and (_05360_, _05359_, _05350_);
  and (_05361_, _05360_, \oc8051_golden_model_1.PSW [7]);
  not (_05362_, _04034_);
  and (_05363_, _04446_, _05362_);
  and (_05364_, _05363_, _05352_);
  and (_05365_, _05364_, _05350_);
  and (_05366_, _05365_, \oc8051_golden_model_1.ACC [7]);
  nor (_05367_, _05366_, _05361_);
  and (_05368_, _05367_, _05356_);
  not (_05369_, _05350_);
  and (_05370_, _04446_, _04034_);
  nand (_05371_, _05370_, _05344_);
  nor (_05372_, _05371_, _05369_);
  and (_05373_, _05372_, \oc8051_golden_model_1.P0INREG [7]);
  not (_05374_, _05373_);
  and (_05375_, _05358_, _05344_);
  and (_05376_, _05375_, _05350_);
  and (_05377_, _05376_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05378_, _05377_);
  and (_05379_, _05363_, _05344_);
  and (_05380_, _05379_, _05350_);
  and (_05381_, _05380_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05382_, _05350_, _05346_);
  and (_05383_, _05382_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05384_, _05383_, _05381_);
  and (_05385_, _05384_, _05378_);
  and (_05386_, _05385_, _05374_);
  and (_05387_, _05386_, _05368_);
  nor (_05388_, _04482_, _04211_);
  and (_05389_, _05388_, _05174_);
  nand (_05390_, _05389_, _03669_);
  nor (_05391_, _05390_, _05371_);
  and (_05392_, _05391_, \oc8051_golden_model_1.PCON [7]);
  not (_05393_, _05392_);
  and (_05394_, _04482_, _04344_);
  and (_05395_, _05394_, _05342_);
  and (_05396_, _05395_, _05375_);
  and (_05397_, _05396_, \oc8051_golden_model_1.SBUF [7]);
  and (_05398_, _05379_, _05343_);
  and (_05399_, _05398_, \oc8051_golden_model_1.IE [7]);
  nor (_05400_, _05399_, _05397_);
  and (_05401_, _05400_, _05393_);
  nor (_05402_, _04165_, _03669_);
  nand (_05403_, _05402_, _05394_);
  nor (_05404_, _05403_, _05371_);
  and (_05405_, _05404_, \oc8051_golden_model_1.TH1 [7]);
  and (_05406_, _05375_, _05343_);
  and (_05407_, _05406_, \oc8051_golden_model_1.SCON [7]);
  nor (_05408_, _05407_, _05405_);
  nor (_05409_, _04482_, _04344_);
  nand (_05410_, _05409_, _05342_);
  nor (_05411_, _05410_, _05371_);
  and (_05412_, _05411_, \oc8051_golden_model_1.TL0 [7]);
  not (_05413_, _05395_);
  nor (_05414_, _05413_, _05371_);
  and (_05415_, _05414_, \oc8051_golden_model_1.TMOD [7]);
  nor (_05416_, _05415_, _05412_);
  and (_05417_, _05416_, _05408_);
  and (_05418_, _05417_, _05401_);
  and (_05419_, _05418_, _05387_);
  not (_05420_, _05388_);
  nor (_05421_, _05420_, _05371_);
  and (_05422_, _05421_, _05349_);
  and (_05423_, _05422_, \oc8051_golden_model_1.DPH [7]);
  not (_05424_, _05423_);
  nand (_05425_, _05402_, _05341_);
  nor (_05426_, _05425_, _05371_);
  and (_05427_, _05426_, \oc8051_golden_model_1.TH0 [7]);
  and (_05428_, _05421_, _05342_);
  and (_05429_, _05428_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05430_, _05429_, _05427_);
  and (_05431_, _05430_, _05424_);
  not (_05432_, _05349_);
  nor (_05433_, _05371_, _05432_);
  and (_05434_, _05433_, _05394_);
  and (_05435_, _05434_, \oc8051_golden_model_1.SP [7]);
  not (_05436_, _05435_);
  not (_05437_, _05343_);
  nor (_05438_, _05371_, _05437_);
  and (_05439_, _05438_, \oc8051_golden_model_1.TCON [7]);
  and (_05440_, _05433_, _05409_);
  and (_05441_, _05440_, \oc8051_golden_model_1.DPL [7]);
  nor (_05442_, _05441_, _05439_);
  and (_05443_, _05442_, _05436_);
  and (_05444_, _05443_, _05431_);
  and (_05445_, _05444_, _05419_);
  not (_05446_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_05447_, _04413_, _05446_);
  not (_05448_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_05449_, _04555_, _05448_);
  and (_05450_, _05449_, _04553_);
  nand (_05451_, _05450_, _05447_);
  not (_05452_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_05453_, _04555_, _05452_);
  not (_05454_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_05455_, _04413_, _05454_);
  and (_05456_, _05455_, _04561_);
  nand (_05457_, _05456_, _05453_);
  nand (_05458_, _05457_, _05451_);
  nand (_05459_, _05458_, _04179_);
  not (_05460_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_05461_, _04555_, _05460_);
  not (_05462_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_05463_, _04413_, _05462_);
  and (_05464_, _05463_, _04561_);
  nand (_05465_, _05464_, _05461_);
  not (_05466_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_05467_, _04413_, _05466_);
  not (_05468_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_05469_, _04555_, _05468_);
  and (_05470_, _05469_, _04553_);
  nand (_05471_, _05470_, _05467_);
  nand (_05472_, _05471_, _05465_);
  nand (_05473_, _05472_, _04568_);
  nand (_05474_, _05473_, _05459_);
  nand (_05475_, _05474_, _04002_);
  nand (_05476_, _04413_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_05477_, _04555_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_05478_, _05477_, _04561_);
  nand (_05479_, _05478_, _05476_);
  nand (_05480_, _04555_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_05481_, _04413_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_05482_, _05481_, _04553_);
  nand (_05483_, _05482_, _05480_);
  nand (_05484_, _05483_, _05479_);
  nand (_05485_, _05484_, _04179_);
  nand (_05486_, _04413_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_05487_, _04555_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_05488_, _05487_, _04561_);
  nand (_05489_, _05488_, _05486_);
  nand (_05490_, _04555_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_05491_, _04413_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_05492_, _05491_, _04553_);
  nand (_05493_, _05492_, _05490_);
  nand (_05494_, _05493_, _05489_);
  nand (_05495_, _05494_, _04568_);
  nand (_05496_, _05495_, _05485_);
  nand (_05497_, _05496_, _04585_);
  nand (_05498_, _05497_, _05475_);
  or (_05499_, _05498_, _03638_);
  and (_05500_, _05499_, _05445_);
  not (_05501_, _05500_);
  and (_05502_, _05360_, \oc8051_golden_model_1.PSW [3]);
  not (_05503_, _05502_);
  and (_05504_, _05347_, \oc8051_golden_model_1.IP [3]);
  not (_05505_, _05504_);
  and (_05506_, _05365_, \oc8051_golden_model_1.ACC [3]);
  and (_05507_, _05354_, \oc8051_golden_model_1.B [3]);
  nor (_05508_, _05507_, _05506_);
  and (_05509_, _05508_, _05505_);
  and (_05510_, _05509_, _05503_);
  and (_05511_, _05426_, \oc8051_golden_model_1.TH0 [3]);
  and (_05512_, _05438_, \oc8051_golden_model_1.TCON [3]);
  nor (_05513_, _05512_, _05511_);
  and (_05514_, _05376_, \oc8051_golden_model_1.P1INREG [3]);
  nand (_05515_, _05388_, _05342_);
  nor (_05516_, _05515_, _05371_);
  and (_05517_, _05516_, \oc8051_golden_model_1.TL1 [3]);
  nor (_05518_, _05517_, _05514_);
  and (_05519_, _05518_, _05513_);
  and (_05520_, _05406_, \oc8051_golden_model_1.SCON [3]);
  and (_05521_, _05404_, \oc8051_golden_model_1.TH1 [3]);
  nor (_05522_, _05521_, _05520_);
  and (_05523_, _05411_, \oc8051_golden_model_1.TL0 [3]);
  and (_05524_, _05414_, \oc8051_golden_model_1.TMOD [3]);
  nor (_05525_, _05524_, _05523_);
  and (_05526_, _05525_, _05522_);
  and (_05527_, _05526_, _05519_);
  and (_05528_, _05527_, _05510_);
  and (_05529_, _05391_, \oc8051_golden_model_1.PCON [3]);
  not (_05530_, _05529_);
  and (_05531_, _05380_, \oc8051_golden_model_1.P2INREG [3]);
  and (_05532_, _05382_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_05533_, _05532_, _05531_);
  and (_05534_, _05533_, _05530_);
  and (_05535_, _05396_, \oc8051_golden_model_1.SBUF [3]);
  and (_05536_, _05398_, \oc8051_golden_model_1.IE [3]);
  nor (_05537_, _05536_, _05535_);
  and (_05538_, _05537_, _05534_);
  and (_05539_, _05372_, \oc8051_golden_model_1.P0INREG [3]);
  not (_05540_, _05539_);
  and (_05541_, _05422_, \oc8051_golden_model_1.DPH [3]);
  not (_05542_, _05541_);
  and (_05543_, _05434_, \oc8051_golden_model_1.SP [3]);
  nand (_05544_, _05409_, _05349_);
  nor (_05545_, _05544_, _05371_);
  and (_05546_, _05545_, \oc8051_golden_model_1.DPL [3]);
  nor (_05547_, _05546_, _05543_);
  and (_05548_, _05547_, _05542_);
  and (_05549_, _05548_, _05540_);
  and (_05550_, _05549_, _05538_);
  and (_05551_, _05550_, _05528_);
  or (_05552_, _05050_, _03638_);
  and (_05553_, _05552_, _05551_);
  not (_05554_, _05553_);
  and (_05555_, _05347_, \oc8051_golden_model_1.IP [1]);
  and (_05556_, _05365_, \oc8051_golden_model_1.ACC [1]);
  nor (_05557_, _05556_, _05555_);
  and (_05558_, _05360_, \oc8051_golden_model_1.PSW [1]);
  and (_05559_, _05354_, \oc8051_golden_model_1.B [1]);
  nor (_05560_, _05559_, _05558_);
  and (_05561_, _05560_, _05557_);
  and (_05562_, _05372_, \oc8051_golden_model_1.P0INREG [1]);
  not (_05563_, _05562_);
  and (_05564_, _05376_, \oc8051_golden_model_1.P1INREG [1]);
  not (_05565_, _05564_);
  and (_05566_, _05380_, \oc8051_golden_model_1.P2INREG [1]);
  and (_05567_, _05382_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_05568_, _05567_, _05566_);
  and (_05569_, _05568_, _05565_);
  and (_05570_, _05569_, _05563_);
  and (_05571_, _05570_, _05561_);
  and (_05572_, _05391_, \oc8051_golden_model_1.PCON [1]);
  not (_05573_, _05572_);
  and (_05574_, _05396_, \oc8051_golden_model_1.SBUF [1]);
  and (_05575_, _05398_, \oc8051_golden_model_1.IE [1]);
  nor (_05576_, _05575_, _05574_);
  and (_05577_, _05576_, _05573_);
  and (_05578_, _05404_, \oc8051_golden_model_1.TH1 [1]);
  and (_05579_, _05406_, \oc8051_golden_model_1.SCON [1]);
  nor (_05580_, _05579_, _05578_);
  and (_05581_, _05414_, \oc8051_golden_model_1.TMOD [1]);
  and (_05582_, _05411_, \oc8051_golden_model_1.TL0 [1]);
  nor (_05583_, _05582_, _05581_);
  and (_05584_, _05583_, _05580_);
  and (_05585_, _05584_, _05577_);
  and (_05586_, _05585_, _05571_);
  and (_05587_, _05422_, \oc8051_golden_model_1.DPH [1]);
  not (_05588_, _05587_);
  and (_05589_, _05426_, \oc8051_golden_model_1.TH0 [1]);
  and (_05590_, _05428_, \oc8051_golden_model_1.TL1 [1]);
  nor (_05591_, _05590_, _05589_);
  and (_05592_, _05591_, _05588_);
  and (_05593_, _05434_, \oc8051_golden_model_1.SP [1]);
  not (_05594_, _05593_);
  and (_05595_, _05438_, \oc8051_golden_model_1.TCON [1]);
  and (_05596_, _05440_, \oc8051_golden_model_1.DPL [1]);
  nor (_05597_, _05596_, _05595_);
  and (_05598_, _05597_, _05594_);
  and (_05599_, _05598_, _05592_);
  and (_05600_, _05599_, _05586_);
  or (_05601_, _04842_, _03638_);
  and (_05602_, _05601_, _05600_);
  not (_05603_, _05602_);
  and (_05604_, _05347_, \oc8051_golden_model_1.IP [0]);
  not (_05605_, _05604_);
  and (_05606_, _05360_, \oc8051_golden_model_1.PSW [0]);
  not (_05607_, _05606_);
  and (_05608_, _05365_, \oc8051_golden_model_1.ACC [0]);
  and (_05609_, _05354_, \oc8051_golden_model_1.B [0]);
  nor (_05610_, _05609_, _05608_);
  and (_05611_, _05610_, _05607_);
  and (_05612_, _05611_, _05605_);
  and (_05613_, _05426_, \oc8051_golden_model_1.TH0 [0]);
  and (_05614_, _05438_, \oc8051_golden_model_1.TCON [0]);
  nor (_05615_, _05614_, _05613_);
  and (_05616_, _05376_, \oc8051_golden_model_1.P1INREG [0]);
  and (_05617_, _05516_, \oc8051_golden_model_1.TL1 [0]);
  nor (_05618_, _05617_, _05616_);
  and (_05619_, _05618_, _05615_);
  and (_05620_, _05406_, \oc8051_golden_model_1.SCON [0]);
  and (_05621_, _05404_, \oc8051_golden_model_1.TH1 [0]);
  nor (_05622_, _05621_, _05620_);
  and (_05623_, _05414_, \oc8051_golden_model_1.TMOD [0]);
  and (_05624_, _05411_, \oc8051_golden_model_1.TL0 [0]);
  nor (_05625_, _05624_, _05623_);
  and (_05626_, _05625_, _05622_);
  and (_05627_, _05626_, _05619_);
  and (_05628_, _05627_, _05612_);
  and (_05629_, _05391_, \oc8051_golden_model_1.PCON [0]);
  not (_05630_, _05629_);
  and (_05631_, _05380_, \oc8051_golden_model_1.P2INREG [0]);
  and (_05632_, _05382_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_05633_, _05632_, _05631_);
  and (_05634_, _05633_, _05630_);
  and (_05635_, _05396_, \oc8051_golden_model_1.SBUF [0]);
  and (_05636_, _05398_, \oc8051_golden_model_1.IE [0]);
  nor (_05637_, _05636_, _05635_);
  and (_05638_, _05637_, _05634_);
  and (_05639_, _05372_, \oc8051_golden_model_1.P0INREG [0]);
  not (_05640_, _05639_);
  and (_05641_, _05422_, \oc8051_golden_model_1.DPH [0]);
  not (_05642_, _05641_);
  and (_05643_, _05434_, \oc8051_golden_model_1.SP [0]);
  and (_05644_, _05545_, \oc8051_golden_model_1.DPL [0]);
  nor (_05645_, _05644_, _05643_);
  and (_05646_, _05645_, _05642_);
  and (_05647_, _05646_, _05640_);
  and (_05648_, _05647_, _05638_);
  and (_05649_, _05648_, _05628_);
  not (_05650_, _05649_);
  and (_05651_, _04608_, _05351_);
  or (_05652_, _05651_, _05650_);
  and (_05653_, _05652_, _05603_);
  and (_05654_, _05347_, \oc8051_golden_model_1.IP [2]);
  and (_05655_, _05365_, \oc8051_golden_model_1.ACC [2]);
  nor (_05656_, _05655_, _05654_);
  and (_05657_, _05360_, \oc8051_golden_model_1.PSW [2]);
  and (_05658_, _05354_, \oc8051_golden_model_1.B [2]);
  nor (_05659_, _05658_, _05657_);
  and (_05660_, _05659_, _05656_);
  and (_05661_, _05438_, \oc8051_golden_model_1.TCON [2]);
  and (_05662_, _05426_, \oc8051_golden_model_1.TH0 [2]);
  nor (_05663_, _05662_, _05661_);
  and (_05664_, _05376_, \oc8051_golden_model_1.P1INREG [2]);
  and (_05665_, _05516_, \oc8051_golden_model_1.TL1 [2]);
  nor (_05666_, _05665_, _05664_);
  and (_05667_, _05666_, _05663_);
  and (_05668_, _05414_, \oc8051_golden_model_1.TMOD [2]);
  and (_05669_, _05411_, \oc8051_golden_model_1.TL0 [2]);
  nor (_05670_, _05669_, _05668_);
  and (_05671_, _05406_, \oc8051_golden_model_1.SCON [2]);
  and (_05672_, _05404_, \oc8051_golden_model_1.TH1 [2]);
  nor (_05673_, _05672_, _05671_);
  and (_05674_, _05673_, _05670_);
  and (_05675_, _05674_, _05667_);
  and (_05676_, _05675_, _05660_);
  and (_05677_, _05391_, \oc8051_golden_model_1.PCON [2]);
  not (_05678_, _05677_);
  and (_05679_, _05396_, \oc8051_golden_model_1.SBUF [2]);
  and (_05680_, _05398_, \oc8051_golden_model_1.IE [2]);
  nor (_05681_, _05680_, _05679_);
  and (_05682_, _05681_, _05678_);
  and (_05683_, _05380_, \oc8051_golden_model_1.P2INREG [2]);
  and (_05684_, _05382_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_05685_, _05684_, _05683_);
  and (_05686_, _05685_, _05682_);
  and (_05687_, _05372_, \oc8051_golden_model_1.P0INREG [2]);
  not (_05688_, _05687_);
  and (_05689_, _05422_, \oc8051_golden_model_1.DPH [2]);
  not (_05690_, _05689_);
  and (_05691_, _05434_, \oc8051_golden_model_1.SP [2]);
  and (_05692_, _05545_, \oc8051_golden_model_1.DPL [2]);
  nor (_05693_, _05692_, _05691_);
  and (_05694_, _05693_, _05690_);
  and (_05695_, _05694_, _05688_);
  and (_05696_, _05695_, _05686_);
  and (_05697_, _05696_, _05676_);
  or (_05698_, _05236_, _03638_);
  and (_05699_, _05698_, _05697_);
  not (_05700_, _05699_);
  and (_05701_, _05700_, _05653_);
  and (_05702_, _05701_, _05554_);
  and (_05703_, _05360_, \oc8051_golden_model_1.PSW [5]);
  and (_05704_, _05354_, \oc8051_golden_model_1.B [5]);
  nor (_05705_, _05704_, _05703_);
  and (_05706_, _05347_, \oc8051_golden_model_1.IP [5]);
  and (_05707_, _05365_, \oc8051_golden_model_1.ACC [5]);
  nor (_05708_, _05707_, _05706_);
  and (_05709_, _05708_, _05705_);
  and (_05710_, _05438_, \oc8051_golden_model_1.TCON [5]);
  and (_05711_, _05426_, \oc8051_golden_model_1.TH0 [5]);
  nor (_05712_, _05711_, _05710_);
  and (_05713_, _05376_, \oc8051_golden_model_1.P1INREG [5]);
  and (_05714_, _05516_, \oc8051_golden_model_1.TL1 [5]);
  nor (_05715_, _05714_, _05713_);
  and (_05716_, _05715_, _05712_);
  and (_05717_, _05414_, \oc8051_golden_model_1.TMOD [5]);
  and (_05718_, _05411_, \oc8051_golden_model_1.TL0 [5]);
  nor (_05719_, _05718_, _05717_);
  and (_05720_, _05406_, \oc8051_golden_model_1.SCON [5]);
  and (_05721_, _05404_, \oc8051_golden_model_1.TH1 [5]);
  nor (_05722_, _05721_, _05720_);
  and (_05723_, _05722_, _05719_);
  and (_05724_, _05723_, _05716_);
  and (_05725_, _05724_, _05709_);
  and (_05726_, _05391_, \oc8051_golden_model_1.PCON [5]);
  not (_05727_, _05726_);
  and (_05728_, _05396_, \oc8051_golden_model_1.SBUF [5]);
  and (_05729_, _05398_, \oc8051_golden_model_1.IE [5]);
  nor (_05730_, _05729_, _05728_);
  and (_05731_, _05730_, _05727_);
  and (_05732_, _05380_, \oc8051_golden_model_1.P2INREG [5]);
  and (_05733_, _05382_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_05734_, _05733_, _05732_);
  and (_05735_, _05734_, _05731_);
  and (_05736_, _05372_, \oc8051_golden_model_1.P0INREG [5]);
  not (_05737_, _05736_);
  and (_05738_, _05422_, \oc8051_golden_model_1.DPH [5]);
  not (_05739_, _05738_);
  and (_05740_, _05434_, \oc8051_golden_model_1.SP [5]);
  and (_05741_, _05545_, \oc8051_golden_model_1.DPL [5]);
  nor (_05742_, _05741_, _05740_);
  and (_05743_, _05742_, _05739_);
  and (_05744_, _05743_, _05737_);
  and (_05745_, _05744_, _05735_);
  and (_05746_, _05745_, _05725_);
  not (_05747_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_05748_, _04413_, _05747_);
  not (_05749_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_05750_, _04555_, _05749_);
  and (_05751_, _05750_, _04553_);
  nand (_05752_, _05751_, _05748_);
  not (_05753_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_05754_, _04555_, _05753_);
  not (_05755_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_05756_, _04413_, _05755_);
  and (_05757_, _05756_, _04561_);
  nand (_05758_, _05757_, _05754_);
  nand (_05759_, _05758_, _05752_);
  nand (_05760_, _05759_, _04179_);
  not (_05761_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_05762_, _04555_, _05761_);
  not (_05763_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_05764_, _04413_, _05763_);
  and (_05765_, _05764_, _04561_);
  nand (_05766_, _05765_, _05762_);
  not (_05767_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_05768_, _04413_, _05767_);
  not (_05769_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_05770_, _04555_, _05769_);
  and (_05771_, _05770_, _04553_);
  nand (_05772_, _05771_, _05768_);
  nand (_05773_, _05772_, _05766_);
  nand (_05774_, _05773_, _04568_);
  nand (_05775_, _05774_, _05760_);
  nand (_05776_, _05775_, _04002_);
  nand (_05777_, _04413_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_05778_, _04555_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_05779_, _05778_, _04561_);
  nand (_05780_, _05779_, _05777_);
  nand (_05781_, _04555_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_05782_, _04413_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_05783_, _05782_, _04553_);
  nand (_05784_, _05783_, _05781_);
  nand (_05785_, _05784_, _05780_);
  nand (_05786_, _05785_, _04179_);
  nand (_05787_, _04413_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_05788_, _04555_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_05789_, _05788_, _04561_);
  nand (_05790_, _05789_, _05787_);
  nand (_05791_, _04555_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand (_05792_, _04413_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_05793_, _05792_, _04553_);
  nand (_05794_, _05793_, _05791_);
  nand (_05795_, _05794_, _05790_);
  nand (_05796_, _05795_, _04568_);
  nand (_05797_, _05796_, _05786_);
  nand (_05798_, _05797_, _04585_);
  nand (_05799_, _05798_, _05776_);
  or (_05800_, _05799_, _03638_);
  and (_05801_, _05800_, _05746_);
  and (_05802_, _05414_, \oc8051_golden_model_1.TMOD [4]);
  not (_05803_, _05802_);
  and (_05804_, _05406_, \oc8051_golden_model_1.SCON [4]);
  and (_05805_, _05396_, \oc8051_golden_model_1.SBUF [4]);
  nor (_05806_, _05805_, _05804_);
  and (_05807_, _05806_, _05803_);
  and (_05808_, _05411_, \oc8051_golden_model_1.TL0 [4]);
  and (_05809_, _05398_, \oc8051_golden_model_1.IE [4]);
  nor (_05810_, _05809_, _05808_);
  and (_05811_, _05426_, \oc8051_golden_model_1.TH0 [4]);
  and (_05812_, _05404_, \oc8051_golden_model_1.TH1 [4]);
  nor (_05813_, _05812_, _05811_);
  and (_05814_, _05813_, _05810_);
  and (_05815_, _05422_, \oc8051_golden_model_1.DPH [4]);
  and (_05816_, _05428_, \oc8051_golden_model_1.TL1 [4]);
  nor (_05817_, _05816_, _05815_);
  and (_05818_, _05817_, _05814_);
  and (_05819_, _05818_, _05807_);
  and (_05820_, _05434_, \oc8051_golden_model_1.SP [4]);
  and (_05821_, _05545_, \oc8051_golden_model_1.DPL [4]);
  nor (_05822_, _05821_, _05820_);
  and (_05823_, _05376_, \oc8051_golden_model_1.P1INREG [4]);
  not (_05824_, _05823_);
  and (_05825_, _05372_, \oc8051_golden_model_1.P0INREG [4]);
  not (_05826_, _05825_);
  and (_05827_, _05380_, \oc8051_golden_model_1.P2INREG [4]);
  and (_05828_, _05382_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_05829_, _05828_, _05827_);
  and (_05830_, _05829_, _05826_);
  and (_05831_, _05830_, _05824_);
  and (_05832_, _05360_, \oc8051_golden_model_1.PSW [4]);
  and (_05833_, _05365_, \oc8051_golden_model_1.ACC [4]);
  nor (_05834_, _05833_, _05832_);
  and (_05835_, _05347_, \oc8051_golden_model_1.IP [4]);
  and (_05836_, _05354_, \oc8051_golden_model_1.B [4]);
  nor (_05837_, _05836_, _05835_);
  and (_05838_, _05837_, _05834_);
  and (_05839_, _05391_, \oc8051_golden_model_1.PCON [4]);
  and (_05840_, _05438_, \oc8051_golden_model_1.TCON [4]);
  nor (_05841_, _05840_, _05839_);
  and (_05842_, _05841_, _05838_);
  and (_05843_, _05842_, _05831_);
  and (_05844_, _05843_, _05822_);
  and (_05845_, _05844_, _05819_);
  not (_05846_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_05847_, _04413_, _05846_);
  not (_05848_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_05849_, _04555_, _05848_);
  and (_05850_, _05849_, _04553_);
  nand (_05851_, _05850_, _05847_);
  not (_05852_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_05853_, _04555_, _05852_);
  not (_05854_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05855_, _04413_, _05854_);
  and (_05856_, _05855_, _04561_);
  nand (_05857_, _05856_, _05853_);
  nand (_05858_, _05857_, _05851_);
  nand (_05859_, _05858_, _04179_);
  not (_05860_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_05861_, _04555_, _05860_);
  not (_05862_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05863_, _04413_, _05862_);
  and (_05864_, _05863_, _04561_);
  nand (_05865_, _05864_, _05861_);
  not (_05866_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_05867_, _04413_, _05866_);
  not (_05868_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_05869_, _04555_, _05868_);
  and (_05870_, _05869_, _04553_);
  nand (_05871_, _05870_, _05867_);
  nand (_05872_, _05871_, _05865_);
  nand (_05873_, _05872_, _04568_);
  nand (_05874_, _05873_, _05859_);
  nand (_05875_, _05874_, _04002_);
  nand (_05876_, _04413_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_05877_, _04555_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_05878_, _05877_, _04561_);
  nand (_05879_, _05878_, _05876_);
  nand (_05880_, _04555_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_05881_, _04413_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_05882_, _05881_, _04553_);
  nand (_05883_, _05882_, _05880_);
  nand (_05884_, _05883_, _05879_);
  nand (_05885_, _05884_, _04179_);
  nand (_05886_, _04413_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_05887_, _04555_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_05888_, _05887_, _04561_);
  nand (_05889_, _05888_, _05886_);
  nand (_05890_, _04555_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_05891_, _04413_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_05892_, _05891_, _04553_);
  nand (_05893_, _05892_, _05890_);
  nand (_05894_, _05893_, _05889_);
  nand (_05895_, _05894_, _04568_);
  nand (_05896_, _05895_, _05885_);
  nand (_05897_, _05896_, _04585_);
  nand (_05898_, _05897_, _05875_);
  or (_05899_, _05898_, _03638_);
  and (_05900_, _05899_, _05845_);
  nor (_05901_, _05900_, _05801_);
  and (_05902_, _05901_, _05702_);
  nor (_05903_, _05902_, _05501_);
  and (_05904_, _05406_, \oc8051_golden_model_1.SCON [6]);
  not (_05905_, _05904_);
  and (_05906_, _05426_, \oc8051_golden_model_1.TH0 [6]);
  and (_05907_, _05396_, \oc8051_golden_model_1.SBUF [6]);
  nor (_05908_, _05907_, _05906_);
  and (_05909_, _05908_, _05905_);
  and (_05910_, _05414_, \oc8051_golden_model_1.TMOD [6]);
  and (_05911_, _05398_, \oc8051_golden_model_1.IE [6]);
  nor (_05912_, _05911_, _05910_);
  and (_05913_, _05411_, \oc8051_golden_model_1.TL0 [6]);
  and (_05914_, _05404_, \oc8051_golden_model_1.TH1 [6]);
  nor (_05915_, _05914_, _05913_);
  and (_05916_, _05915_, _05912_);
  and (_05917_, _05422_, \oc8051_golden_model_1.DPH [6]);
  and (_05918_, _05428_, \oc8051_golden_model_1.TL1 [6]);
  nor (_05919_, _05918_, _05917_);
  and (_05920_, _05919_, _05916_);
  and (_05921_, _05920_, _05909_);
  and (_05922_, _05434_, \oc8051_golden_model_1.SP [6]);
  and (_05923_, _05545_, \oc8051_golden_model_1.DPL [6]);
  nor (_05924_, _05923_, _05922_);
  and (_05925_, _05376_, \oc8051_golden_model_1.P1INREG [6]);
  not (_05926_, _05925_);
  and (_05927_, _05372_, \oc8051_golden_model_1.P0INREG [6]);
  not (_05928_, _05927_);
  and (_05929_, _05380_, \oc8051_golden_model_1.P2INREG [6]);
  and (_05930_, _05382_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_05931_, _05930_, _05929_);
  and (_05932_, _05931_, _05928_);
  and (_05933_, _05932_, _05926_);
  and (_05934_, _05347_, \oc8051_golden_model_1.IP [6]);
  and (_05935_, _05365_, \oc8051_golden_model_1.ACC [6]);
  nor (_05936_, _05935_, _05934_);
  and (_05937_, _05360_, \oc8051_golden_model_1.PSW [6]);
  and (_05938_, _05354_, \oc8051_golden_model_1.B [6]);
  nor (_05939_, _05938_, _05937_);
  and (_05940_, _05939_, _05936_);
  and (_05941_, _05391_, \oc8051_golden_model_1.PCON [6]);
  and (_05942_, _05438_, \oc8051_golden_model_1.TCON [6]);
  nor (_05943_, _05942_, _05941_);
  and (_05944_, _05943_, _05940_);
  and (_05945_, _05944_, _05933_);
  and (_05946_, _05945_, _05924_);
  and (_05947_, _05946_, _05921_);
  not (_05948_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_05949_, _04413_, _05948_);
  not (_05951_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_05952_, _04555_, _05951_);
  and (_05954_, _05952_, _04553_);
  nand (_05955_, _05954_, _05949_);
  not (_05957_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_05958_, _04555_, _05957_);
  not (_05960_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_05961_, _04413_, _05960_);
  and (_05963_, _05961_, _04561_);
  nand (_05964_, _05963_, _05958_);
  nand (_05966_, _05964_, _05955_);
  nand (_05967_, _05966_, _04179_);
  not (_05969_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_05970_, _04555_, _05969_);
  not (_05972_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_05973_, _04413_, _05972_);
  and (_05975_, _05973_, _04561_);
  nand (_05976_, _05975_, _05970_);
  not (_05978_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_05979_, _04413_, _05978_);
  not (_05981_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_05982_, _04555_, _05981_);
  and (_05984_, _05982_, _04553_);
  nand (_05985_, _05984_, _05979_);
  nand (_05987_, _05985_, _05976_);
  nand (_05988_, _05987_, _04568_);
  nand (_05989_, _05988_, _05967_);
  nand (_05990_, _05989_, _04002_);
  nand (_05991_, _04413_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_05992_, _04555_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_05993_, _05992_, _04561_);
  nand (_05994_, _05993_, _05991_);
  nand (_05995_, _04555_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_05996_, _04413_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_05997_, _05996_, _04553_);
  nand (_05998_, _05997_, _05995_);
  nand (_05999_, _05998_, _05994_);
  nand (_06000_, _05999_, _04179_);
  nand (_06001_, _04413_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_06002_, _04555_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_06003_, _06002_, _04561_);
  nand (_06004_, _06003_, _06001_);
  nand (_06005_, _04555_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_06006_, _04413_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_06007_, _06006_, _04553_);
  nand (_06008_, _06007_, _06005_);
  nand (_06009_, _06008_, _06004_);
  nand (_06010_, _06009_, _04568_);
  nand (_06011_, _06010_, _06000_);
  nand (_06012_, _06011_, _04585_);
  nand (_06013_, _06012_, _05990_);
  or (_06014_, _06013_, _03638_);
  and (_06015_, _06014_, _05947_);
  and (_06016_, _06015_, _05500_);
  nor (_06017_, _06015_, _05500_);
  nor (_06018_, _06017_, _06016_);
  not (_06019_, _06018_);
  and (_06020_, _06019_, _05902_);
  nor (_06021_, _06020_, _05903_);
  and (_06022_, _06021_, _04742_);
  and (_06023_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_06024_, _06023_, \oc8051_golden_model_1.PC [6]);
  and (_06025_, _06024_, _03514_);
  and (_06026_, _06025_, \oc8051_golden_model_1.PC [7]);
  nor (_06027_, _06025_, \oc8051_golden_model_1.PC [7]);
  nor (_06028_, _06027_, _06026_);
  and (_06029_, _06028_, _03474_);
  not (_06030_, _04707_);
  and (_06031_, _03934_, _01988_);
  and (_06032_, _03907_, _01979_);
  nor (_06033_, _06032_, _06031_);
  and (_06034_, _03898_, _01991_);
  and (_06035_, _03939_, _01954_);
  nor (_06036_, _06035_, _06034_);
  and (_06037_, _06036_, _06033_);
  and (_06038_, _03918_, _01933_);
  and (_06039_, _03941_, _01961_);
  nor (_06040_, _06039_, _06038_);
  and (_06041_, _03928_, _01943_);
  and (_06042_, _03930_, _01948_);
  nor (_06043_, _06042_, _06041_);
  and (_06044_, _06043_, _06040_);
  and (_06046_, _06044_, _06037_);
  and (_06048_, _03925_, _01994_);
  and (_06049_, _03923_, _01985_);
  nor (_06051_, _06049_, _06048_);
  and (_06052_, _03911_, _01966_);
  and (_06054_, _03916_, _01929_);
  nor (_06055_, _06054_, _06052_);
  and (_06057_, _06055_, _06051_);
  and (_06058_, _03894_, _01976_);
  and (_06060_, _03936_, _01893_);
  nor (_06061_, _06060_, _06058_);
  and (_06063_, _03913_, _01970_);
  and (_06064_, _03903_, _01939_);
  nor (_06066_, _06064_, _06063_);
  and (_06067_, _06066_, _06061_);
  and (_06069_, _06067_, _06057_);
  and (_06070_, _06069_, _06046_);
  nor (_06072_, _06070_, _05500_);
  and (_06073_, _06072_, _04709_);
  not (_06075_, _03670_);
  nor (_06076_, _04447_, _06075_);
  nor (_06078_, _04035_, _03744_);
  and (_06079_, _06078_, _06076_);
  not (_06080_, _06079_);
  nor (_06081_, _06080_, _05371_);
  and (_06082_, _06081_, \oc8051_golden_model_1.TCON [7]);
  not (_06083_, _04035_);
  and (_06084_, _06083_, _03744_);
  and (_06085_, _06084_, _06076_);
  and (_06086_, _06085_, _05364_);
  and (_06087_, _06086_, \oc8051_golden_model_1.ACC [7]);
  nor (_06088_, _06087_, _06082_);
  and (_06089_, _06079_, _05346_);
  and (_06090_, _06089_, \oc8051_golden_model_1.IP [7]);
  not (_06091_, _06090_);
  and (_06092_, _06085_, _05359_);
  and (_06093_, _06092_, \oc8051_golden_model_1.PSW [7]);
  and (_06094_, _06085_, _05353_);
  and (_06095_, _06094_, \oc8051_golden_model_1.B [7]);
  nor (_06096_, _06095_, _06093_);
  and (_06097_, _06096_, _06091_);
  and (_06098_, _06097_, _06088_);
  and (_06099_, _06079_, _05375_);
  and (_06100_, _06099_, \oc8051_golden_model_1.SCON [7]);
  and (_06101_, _06079_, _05379_);
  and (_06102_, _06101_, \oc8051_golden_model_1.IE [7]);
  nor (_06103_, _06102_, _06100_);
  and (_06104_, _06085_, _05379_);
  and (_06105_, _06104_, \oc8051_golden_model_1.P2INREG [7]);
  and (_06106_, _06085_, _05346_);
  and (_06107_, _06106_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06108_, _06107_, _06105_);
  not (_06109_, _06085_);
  nor (_06110_, _06109_, _05371_);
  and (_06111_, _06110_, \oc8051_golden_model_1.P0INREG [7]);
  and (_06112_, _06085_, _05375_);
  and (_06113_, _06112_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_06114_, _06113_, _06111_);
  and (_06115_, _06114_, _06108_);
  and (_06116_, _06115_, _06103_);
  and (_06117_, _06116_, _06098_);
  and (_06118_, _06117_, _05499_);
  nor (_06119_, _06118_, _05389_);
  and (_06120_, _05389_, \oc8051_golden_model_1.PSW [7]);
  nor (_06121_, _06120_, _06119_);
  nor (_06122_, _06121_, _05114_);
  not (_06123_, _03694_);
  or (_06124_, _06119_, _06123_);
  not (_06125_, _04629_);
  not (_06126_, _05389_);
  nand (_06127_, _06118_, _06126_);
  or (_06128_, _06127_, _06125_);
  not (_06129_, _05498_);
  and (_06130_, _05898_, _05799_);
  nor (_06131_, _04813_, _04608_);
  and (_06132_, _05236_, _05050_);
  and (_06133_, _06132_, _06131_);
  and (_06134_, _06133_, _06130_);
  and (_06135_, _06134_, _06013_);
  or (_06136_, _06135_, _06129_);
  nand (_06137_, _06135_, _06129_);
  and (_06138_, _06137_, _06136_);
  nor (_06139_, _03849_, _03444_);
  nor (_06140_, _06139_, _05243_);
  or (_06141_, _06140_, _06138_);
  not (_06142_, \oc8051_golden_model_1.ACC [7]);
  nor (_06143_, _04111_, _06142_);
  or (_06144_, _06143_, _04963_);
  or (_06145_, _06139_, _04952_);
  and (_06146_, _06028_, _04111_);
  or (_06147_, _06146_, _06145_);
  or (_06148_, _06147_, _06144_);
  and (_06149_, _06148_, _06141_);
  or (_06150_, _06149_, _04624_);
  nor (_06151_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_06152_, _06151_, _04125_);
  nor (_06153_, _06152_, _03754_);
  nor (_06154_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_06155_, _06154_, _03754_);
  and (_06156_, _06155_, _03674_);
  nor (_06157_, _06156_, _06153_);
  nor (_06158_, _06157_, _04126_);
  not (_06159_, _06158_);
  nand (_06160_, _05050_, _04663_);
  not (_06161_, _04126_);
  and (_06162_, _04269_, _03669_);
  nor (_06163_, _06162_, _06161_);
  nand (_06164_, _06163_, _06160_);
  and (_06165_, _06164_, _06159_);
  not (_06166_, _06165_);
  nor (_06167_, _06151_, _04125_);
  nor (_06168_, _06167_, _06152_);
  nor (_06169_, _06168_, _04126_);
  not (_06170_, _06169_);
  nand (_06171_, _05236_, _04663_);
  and (_06172_, _04269_, _04165_);
  nor (_06173_, _06172_, _06161_);
  nand (_06174_, _06173_, _06171_);
  and (_06175_, _06174_, _06170_);
  or (_06176_, _04608_, _04269_);
  and (_06177_, _04269_, _04211_);
  nor (_06178_, _06177_, _06161_);
  nand (_06179_, _06178_, _06176_);
  nor (_06180_, _04126_, \oc8051_golden_model_1.SP [0]);
  not (_06181_, _06180_);
  and (_06182_, _06181_, _06179_);
  or (_06183_, _06182_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor (_06184_, _04754_, _04126_);
  not (_06185_, _06184_);
  and (_06186_, _04813_, _04663_);
  nor (_06187_, _04482_, _04663_);
  or (_06188_, _06187_, _06161_);
  or (_06189_, _06188_, _06186_);
  nand (_06190_, _06189_, _06185_);
  nand (_06191_, _06181_, _06179_);
  or (_06192_, _06191_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_06193_, _06192_, _06190_);
  and (_06194_, _06193_, _06183_);
  or (_06195_, _06191_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_06196_, _06189_, _06185_);
  or (_06197_, _06182_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_06198_, _06197_, _06196_);
  and (_06199_, _06198_, _06195_);
  nor (_06200_, _06199_, _06194_);
  nand (_06201_, _06200_, _06175_);
  not (_06202_, _06175_);
  or (_06203_, _06182_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_06204_, _06191_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_06205_, _06204_, _06190_);
  and (_06206_, _06205_, _06203_);
  or (_06207_, _06191_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_06208_, _06182_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_06209_, _06208_, _06196_);
  and (_06210_, _06209_, _06207_);
  nor (_06211_, _06210_, _06206_);
  nand (_06212_, _06211_, _06202_);
  nand (_06213_, _06212_, _06201_);
  nand (_06214_, _06213_, _06166_);
  or (_06215_, _06182_, _05448_);
  or (_06216_, _06191_, _05446_);
  and (_06217_, _06216_, _06190_);
  nand (_06218_, _06217_, _06215_);
  or (_06219_, _06191_, _05454_);
  or (_06220_, _06182_, _05452_);
  and (_06221_, _06220_, _06196_);
  nand (_06222_, _06221_, _06219_);
  nand (_06223_, _06222_, _06218_);
  nand (_06224_, _06223_, _06175_);
  or (_06225_, _06191_, _05466_);
  or (_06226_, _06182_, _05468_);
  and (_06227_, _06226_, _06190_);
  nand (_06228_, _06227_, _06225_);
  or (_06229_, _06191_, _05462_);
  or (_06230_, _06182_, _05460_);
  and (_06231_, _06230_, _06196_);
  nand (_06232_, _06231_, _06229_);
  nand (_06233_, _06232_, _06228_);
  nand (_06234_, _06233_, _06202_);
  nand (_06235_, _06234_, _06224_);
  nand (_06236_, _06235_, _06165_);
  and (_06237_, _06236_, _06214_);
  or (_06238_, _06237_, _04625_);
  and (_06239_, _06238_, _06150_);
  or (_06240_, _06239_, _04631_);
  and (_06241_, _05900_, _05801_);
  or (_06242_, _05652_, _05603_);
  and (_06243_, _05699_, _05553_);
  not (_06244_, _06243_);
  nor (_06245_, _06244_, _06242_);
  and (_06246_, _06245_, _06241_);
  and (_06247_, _06246_, _06015_);
  or (_06248_, _06247_, _05501_);
  nand (_06249_, _06247_, _05501_);
  and (_06250_, _06249_, _06248_);
  or (_06251_, _06250_, _04816_);
  and (_06252_, _06251_, _06240_);
  or (_06253_, _06252_, _04629_);
  and (_06254_, _06253_, _06128_);
  or (_06255_, _06254_, _04933_);
  nor (_06256_, _06028_, _03445_);
  nor (_06257_, _06256_, _04640_);
  and (_06258_, _06257_, _06255_);
  and (_06259_, _06129_, _04640_);
  or (_06260_, _06259_, _03694_);
  or (_06261_, _06260_, _06258_);
  and (_06262_, _06261_, _06124_);
  or (_06263_, _06262_, _03690_);
  nand (_06264_, _05500_, _03690_);
  and (_06265_, _06264_, _03688_);
  and (_06266_, _06265_, _06263_);
  nor (_06267_, _06118_, _06126_);
  not (_06268_, _06267_);
  and (_06269_, _06268_, _06127_);
  and (_06270_, _06269_, _03687_);
  or (_06271_, _06270_, _06266_);
  and (_06272_, _06271_, _03442_);
  not (_06273_, _06028_);
  or (_06274_, _06273_, _03442_);
  nand (_06275_, _06274_, _03807_);
  or (_06276_, _06275_, _06272_);
  nand (_06277_, _05500_, _03808_);
  and (_06278_, _06277_, _06276_);
  or (_06279_, _06278_, _04269_);
  nand (_06280_, _06236_, _06214_);
  or (_06281_, _06280_, _03638_);
  and (_06282_, _05445_, _04269_);
  nand (_06283_, _06282_, _06281_);
  and (_06284_, _06283_, _05114_);
  and (_06285_, _06284_, _06279_);
  or (_06286_, _06285_, _06122_);
  and (_06287_, _06286_, _03418_);
  or (_06288_, _06273_, _03418_);
  nand (_06289_, _06288_, _04677_);
  or (_06290_, _06289_, _06287_);
  not (_06291_, _04677_);
  nand (_06292_, _05498_, _06291_);
  and (_06293_, _06292_, _06290_);
  or (_06294_, _06293_, _04680_);
  nor (_06295_, _03638_, _03415_);
  not (_06296_, _06295_);
  nand (_06297_, _04672_, _03853_);
  or (_06298_, _06237_, _06297_);
  and (_06299_, _06298_, _06296_);
  and (_06300_, _06299_, _06294_);
  nor (_06301_, _04971_, _04953_);
  not (_06302_, _04964_);
  nor (_06303_, _04961_, _04689_);
  and (_06304_, _06303_, _06302_);
  and (_06305_, _06304_, _06301_);
  not (_06306_, _06305_);
  not (_06307_, _06070_);
  nor (_06308_, _06307_, _05498_);
  and (_06309_, _03898_, _02315_);
  and (_06310_, _03928_, _02349_);
  nor (_06311_, _06310_, _06309_);
  and (_06312_, _03903_, _02335_);
  and (_06313_, _03939_, _02346_);
  nor (_06314_, _06313_, _06312_);
  and (_06315_, _06314_, _06311_);
  and (_06316_, _03934_, _02323_);
  and (_06317_, _03925_, _02331_);
  nor (_06318_, _06317_, _06316_);
  and (_06319_, _03911_, _02313_);
  and (_06320_, _03918_, _02353_);
  nor (_06321_, _06320_, _06319_);
  and (_06322_, _06321_, _06318_);
  and (_06323_, _06322_, _06315_);
  and (_06324_, _03930_, _02327_);
  and (_06325_, _03923_, _02329_);
  nor (_06326_, _06325_, _06324_);
  and (_06327_, _03916_, _02351_);
  and (_06328_, _03907_, _02337_);
  nor (_06329_, _06328_, _06327_);
  and (_06330_, _06329_, _06326_);
  and (_06331_, _03894_, _02317_);
  and (_06332_, _03941_, _02344_);
  nor (_06333_, _06332_, _06331_);
  and (_06334_, _03913_, _02342_);
  and (_06335_, _03936_, _02321_);
  nor (_06336_, _06335_, _06334_);
  and (_06337_, _06336_, _06333_);
  and (_06338_, _06337_, _06330_);
  and (_06339_, _06338_, _06323_);
  and (_06340_, _03918_, _02399_);
  and (_06341_, _03930_, _02373_);
  nor (_06342_, _06341_, _06340_);
  and (_06343_, _03934_, _02369_);
  and (_06344_, _03928_, _02395_);
  nor (_06345_, _06344_, _06343_);
  and (_06346_, _06345_, _06342_);
  and (_06347_, _03936_, _02367_);
  and (_06348_, _03923_, _02375_);
  nor (_06349_, _06348_, _06347_);
  and (_06350_, _03939_, _02392_);
  and (_06351_, _03907_, _02383_);
  nor (_06352_, _06351_, _06350_);
  and (_06353_, _06352_, _06349_);
  and (_06354_, _06353_, _06346_);
  and (_06355_, _03913_, _02388_);
  and (_06356_, _03916_, _02397_);
  nor (_06357_, _06356_, _06355_);
  and (_06358_, _03903_, _02381_);
  and (_06359_, _03941_, _02390_);
  nor (_06360_, _06359_, _06358_);
  and (_06361_, _06360_, _06357_);
  and (_06362_, _03898_, _02361_);
  and (_06363_, _03894_, _02363_);
  nor (_06364_, _06363_, _06362_);
  and (_06365_, _03911_, _02359_);
  and (_06366_, _03925_, _02377_);
  nor (_06367_, _06366_, _06365_);
  and (_06368_, _06367_, _06364_);
  and (_06369_, _06368_, _06361_);
  and (_06370_, _06369_, _06354_);
  not (_06371_, _06370_);
  and (_06372_, _06371_, _06339_);
  and (_06373_, _04515_, _04326_);
  and (_06374_, _04077_, _03946_);
  and (_06375_, _06374_, _06373_);
  and (_06376_, _03934_, _02426_);
  and (_06377_, _03925_, _02413_);
  nor (_06378_, _06377_, _06376_);
  and (_06379_, _03911_, _02409_);
  and (_06380_, _03936_, _02405_);
  nor (_06381_, _06380_, _06379_);
  and (_06382_, _06381_, _06378_);
  and (_06383_, _03898_, _02435_);
  and (_06384_, _03928_, _02407_);
  nor (_06385_, _06384_, _06383_);
  and (_06386_, _03903_, _02447_);
  and (_06387_, _03907_, _02439_);
  nor (_06388_, _06387_, _06386_);
  and (_06389_, _06388_, _06385_);
  and (_06390_, _06389_, _06382_);
  and (_06391_, _03913_, _02423_);
  and (_06392_, _03894_, _02421_);
  nor (_06393_, _06392_, _06391_);
  and (_06394_, _03918_, _02437_);
  and (_06395_, _03923_, _02415_);
  nor (_06396_, _06395_, _06394_);
  and (_06397_, _06396_, _06393_);
  and (_06398_, _03916_, _02429_);
  and (_06399_, _03941_, _02433_);
  nor (_06400_, _06399_, _06398_);
  and (_06401_, _03930_, _02417_);
  and (_06402_, _03939_, _02445_);
  nor (_06403_, _06402_, _06401_);
  and (_06404_, _06403_, _06400_);
  and (_06405_, _06404_, _06397_);
  and (_06406_, _06405_, _06390_);
  nor (_06407_, _06406_, _06070_);
  and (_06408_, _06407_, _06375_);
  and (_06409_, _06408_, _06372_);
  and (_06410_, _06409_, \oc8051_golden_model_1.ACC [7]);
  nor (_06411_, _06370_, _06339_);
  and (_06412_, _06411_, _06408_);
  and (_06413_, _06412_, \oc8051_golden_model_1.B [7]);
  nor (_06414_, _06413_, _06410_);
  not (_06415_, _03946_);
  and (_06416_, _04077_, _06415_);
  and (_06417_, _06416_, _06373_);
  and (_06418_, _06406_, _06307_);
  and (_06419_, _06418_, _06411_);
  and (_06420_, _06419_, _06417_);
  and (_06421_, _06420_, \oc8051_golden_model_1.IP [7]);
  not (_06422_, _06339_);
  and (_06423_, _06370_, _06422_);
  and (_06424_, _06423_, _06408_);
  and (_06425_, _06424_, \oc8051_golden_model_1.PSW [7]);
  nor (_06426_, _06425_, _06421_);
  and (_06427_, _06426_, _06414_);
  not (_06428_, _04326_);
  and (_06429_, _04515_, _06428_);
  and (_06430_, _06370_, _06339_);
  and (_06431_, _06430_, _06418_);
  nor (_06432_, _04077_, _03946_);
  and (_06433_, _06432_, _06431_);
  and (_06434_, _06433_, _06429_);
  and (_06435_, _06434_, \oc8051_golden_model_1.TH1 [7]);
  not (_06436_, _06435_);
  and (_06437_, _06431_, _06374_);
  and (_06438_, _06437_, _06429_);
  and (_06439_, _06438_, \oc8051_golden_model_1.SP [7]);
  not (_06440_, _04515_);
  and (_06441_, _06440_, _04326_);
  and (_06442_, _06431_, _06416_);
  and (_06443_, _06442_, _06441_);
  and (_06444_, _06443_, \oc8051_golden_model_1.TL0 [7]);
  nor (_06445_, _06444_, _06439_);
  and (_06446_, _06445_, _06436_);
  and (_06447_, _06446_, _06427_);
  and (_06448_, _06433_, _06373_);
  and (_06449_, _06448_, \oc8051_golden_model_1.TH0 [7]);
  nor (_06450_, _04515_, _04326_);
  and (_06451_, _06450_, _06431_);
  and (_06452_, _06451_, _06416_);
  and (_06453_, _06452_, \oc8051_golden_model_1.TL1 [7]);
  nor (_06454_, _06453_, _06449_);
  and (_06455_, _06431_, _06417_);
  and (_06456_, _06455_, \oc8051_golden_model_1.TCON [7]);
  not (_06457_, _04077_);
  and (_06458_, _06457_, _03946_);
  and (_06459_, _06458_, _06451_);
  and (_06460_, _06459_, \oc8051_golden_model_1.PCON [7]);
  nor (_06461_, _06460_, _06456_);
  and (_06462_, _06461_, _06454_);
  and (_06463_, _06441_, _06437_);
  and (_06464_, _06463_, \oc8051_golden_model_1.DPL [7]);
  not (_06465_, _06464_);
  and (_06466_, _06431_, _06375_);
  and (_06467_, _06466_, \oc8051_golden_model_1.P0INREG [7]);
  not (_06468_, _06467_);
  and (_06469_, _06423_, _06418_);
  and (_06470_, _06469_, _06375_);
  and (_06471_, _06470_, \oc8051_golden_model_1.P1INREG [7]);
  not (_06472_, _06471_);
  and (_06473_, _06418_, _06372_);
  and (_06474_, _06473_, _06375_);
  and (_06475_, _06474_, \oc8051_golden_model_1.P2INREG [7]);
  and (_06476_, _06419_, _06375_);
  and (_06477_, _06476_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06478_, _06477_, _06475_);
  and (_06479_, _06478_, _06472_);
  and (_06480_, _06479_, _06468_);
  and (_06481_, _06480_, _06465_);
  and (_06482_, _06473_, _06417_);
  and (_06483_, _06482_, \oc8051_golden_model_1.IE [7]);
  and (_06484_, _06429_, _06416_);
  and (_06485_, _06484_, _06469_);
  and (_06486_, _06485_, \oc8051_golden_model_1.SBUF [7]);
  and (_06487_, _06469_, _06417_);
  and (_06488_, _06487_, \oc8051_golden_model_1.SCON [7]);
  or (_06489_, _06488_, _06486_);
  nor (_06490_, _06489_, _06483_);
  and (_06491_, _06451_, _06374_);
  and (_06492_, _06491_, \oc8051_golden_model_1.DPH [7]);
  and (_06493_, _06442_, _06429_);
  and (_06494_, _06493_, \oc8051_golden_model_1.TMOD [7]);
  nor (_06495_, _06494_, _06492_);
  and (_06496_, _06495_, _06490_);
  and (_06497_, _06496_, _06481_);
  and (_06498_, _06497_, _06462_);
  and (_06499_, _06498_, _06447_);
  not (_06500_, _06499_);
  nor (_06501_, _06500_, _06308_);
  nor (_06502_, _06501_, _06296_);
  or (_06503_, _06502_, _06306_);
  or (_06504_, _06503_, _06300_);
  nor (_06505_, _06305_, _03638_);
  nor (_06506_, _06505_, _04695_);
  and (_06507_, _06506_, _06504_);
  and (_06508_, _06307_, _04695_);
  or (_06509_, _06508_, _03483_);
  or (_06510_, _06509_, _06507_);
  and (_06511_, _06273_, _03483_);
  nor (_06512_, _06511_, _04704_);
  and (_06513_, _06512_, _06510_);
  and (_06514_, _06070_, _05500_);
  nor (_06515_, _06514_, _06072_);
  nor (_06516_, _06515_, _04702_);
  nor (_06517_, _06516_, _04705_);
  or (_06518_, _06517_, _06513_);
  not (_06519_, _04709_);
  not (_06520_, _04702_);
  nor (_06521_, _05500_, _06142_);
  and (_06522_, _05500_, _06142_);
  nor (_06523_, _06522_, _06521_);
  or (_06524_, _06523_, _06520_);
  and (_06525_, _06524_, _06519_);
  and (_06526_, _06525_, _06518_);
  or (_06527_, _06526_, _06073_);
  and (_06528_, _06527_, _06030_);
  and (_06529_, _06521_, _04707_);
  or (_06530_, _06529_, _03477_);
  or (_06531_, _06530_, _06528_);
  not (_06532_, _03835_);
  nor (_06533_, _06532_, _03638_);
  and (_06534_, _06273_, _03477_);
  nor (_06535_, _06534_, _06533_);
  and (_06536_, _06535_, _06531_);
  not (_06537_, _03954_);
  nor (_06538_, _06537_, _03638_);
  not (_06539_, _06533_);
  nor (_06540_, _06514_, _06539_);
  or (_06541_, _06540_, _06538_);
  or (_06542_, _06541_, _06536_);
  not (_06543_, _03474_);
  nand (_06544_, _06522_, _06538_);
  and (_06545_, _06544_, _06543_);
  and (_06546_, _06545_, _06542_);
  or (_06547_, _06546_, _06029_);
  not (_06548_, _04891_);
  and (_06549_, _04671_, _03254_);
  not (_06550_, _06549_);
  and (_06551_, _04220_, _03254_);
  not (_06552_, _06551_);
  nand (_06553_, _03867_, _03254_);
  and (_06554_, _06553_, _06552_);
  and (_06555_, _06554_, _06550_);
  and (_06556_, _06555_, _06548_);
  and (_06557_, _06556_, _06547_);
  not (_06558_, _06556_);
  and (_06559_, _06558_, _06138_);
  or (_06560_, _06559_, _04727_);
  or (_06561_, _06560_, _06557_);
  not (_06562_, _04726_);
  or (_06563_, _06182_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_06564_, _06191_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_06565_, _06564_, _06190_);
  and (_06566_, _06565_, _06563_);
  or (_06567_, _06191_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_06568_, _06182_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_06569_, _06568_, _06196_);
  and (_06570_, _06569_, _06567_);
  nor (_06571_, _06570_, _06566_);
  nand (_06572_, _06571_, _06175_);
  or (_06573_, _06182_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_06574_, _06191_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_06575_, _06574_, _06190_);
  and (_06576_, _06575_, _06573_);
  or (_06577_, _06191_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_06578_, _06182_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_06579_, _06578_, _06196_);
  and (_06580_, _06579_, _06577_);
  nor (_06581_, _06580_, _06576_);
  nand (_06582_, _06581_, _06202_);
  nand (_06583_, _06582_, _06572_);
  nand (_06584_, _06583_, _06166_);
  or (_06585_, _06182_, _05951_);
  or (_06586_, _06191_, _05948_);
  and (_06587_, _06586_, _06190_);
  nand (_06588_, _06587_, _06585_);
  or (_06589_, _06191_, _05960_);
  or (_06590_, _06182_, _05957_);
  and (_06591_, _06590_, _06196_);
  nand (_06592_, _06591_, _06589_);
  nand (_06593_, _06592_, _06588_);
  nand (_06594_, _06593_, _06175_);
  or (_06595_, _06191_, _05978_);
  or (_06596_, _06182_, _05981_);
  and (_06597_, _06596_, _06190_);
  nand (_06598_, _06597_, _06595_);
  or (_06599_, _06191_, _05972_);
  or (_06600_, _06182_, _05969_);
  and (_06601_, _06600_, _06196_);
  nand (_06602_, _06601_, _06599_);
  nand (_06603_, _06602_, _06598_);
  nand (_06604_, _06603_, _06202_);
  nand (_06605_, _06604_, _06594_);
  nand (_06606_, _06605_, _06165_);
  nand (_06607_, _06606_, _06584_);
  or (_06608_, _06182_, \oc8051_golden_model_1.IRAM[9] [1]);
  or (_06609_, _06191_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_06610_, _06609_, _06190_);
  and (_06611_, _06610_, _06608_);
  or (_06612_, _06191_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_06613_, _06182_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_06614_, _06613_, _06196_);
  and (_06615_, _06614_, _06612_);
  nor (_06616_, _06615_, _06611_);
  nand (_06617_, _06616_, _06175_);
  or (_06618_, _06182_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_06619_, _06191_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_06620_, _06619_, _06190_);
  and (_06621_, _06620_, _06618_);
  or (_06622_, _06191_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_06623_, _06182_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_06624_, _06623_, _06196_);
  and (_06625_, _06624_, _06622_);
  nor (_06626_, _06625_, _06621_);
  nand (_06627_, _06626_, _06202_);
  nand (_06628_, _06627_, _06617_);
  nand (_06629_, _06628_, _06166_);
  or (_06630_, _06182_, _04763_);
  or (_06631_, _06191_, _04761_);
  and (_06632_, _06631_, _06190_);
  nand (_06633_, _06632_, _06630_);
  or (_06634_, _06191_, _04769_);
  or (_06635_, _06182_, _04767_);
  and (_06636_, _06635_, _06196_);
  nand (_06637_, _06636_, _06634_);
  nand (_06638_, _06637_, _06633_);
  nand (_06639_, _06638_, _06175_);
  or (_06640_, _06191_, _04781_);
  or (_06641_, _06182_, _04783_);
  and (_06642_, _06641_, _06190_);
  nand (_06643_, _06642_, _06640_);
  or (_06644_, _06191_, _04777_);
  or (_06645_, _06182_, _04775_);
  and (_06646_, _06645_, _06196_);
  nand (_06647_, _06646_, _06644_);
  nand (_06648_, _06647_, _06643_);
  nand (_06650_, _06648_, _06202_);
  nand (_06651_, _06650_, _06639_);
  nand (_06652_, _06651_, _06165_);
  nand (_06653_, _06652_, _06629_);
  or (_06654_, _06182_, \oc8051_golden_model_1.IRAM[9] [0]);
  or (_06655_, _06191_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_06656_, _06655_, _06190_);
  and (_06657_, _06656_, _06654_);
  or (_06658_, _06191_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_06659_, _06182_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_06660_, _06659_, _06196_);
  and (_06661_, _06660_, _06658_);
  nor (_06662_, _06661_, _06657_);
  nand (_06663_, _06662_, _06175_);
  or (_06664_, _06182_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_06665_, _06191_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_06666_, _06665_, _06190_);
  and (_06667_, _06666_, _06664_);
  or (_06668_, _06191_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_06669_, _06182_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_06670_, _06669_, _06196_);
  and (_06671_, _06670_, _06668_);
  nor (_06672_, _06671_, _06667_);
  nand (_06673_, _06672_, _06202_);
  nand (_06674_, _06673_, _06663_);
  nand (_06675_, _06674_, _06166_);
  or (_06676_, _06182_, _04554_);
  or (_06677_, _06191_, _04180_);
  and (_06678_, _06677_, _06190_);
  nand (_06679_, _06678_, _06676_);
  or (_06680_, _06191_, _04562_);
  or (_06681_, _06182_, _04559_);
  and (_06682_, _06681_, _06196_);
  nand (_06683_, _06682_, _06680_);
  nand (_06684_, _06683_, _06679_);
  nand (_06685_, _06684_, _06175_);
  or (_06686_, _06191_, _04575_);
  or (_06687_, _06182_, _04577_);
  and (_06688_, _06687_, _06190_);
  nand (_06689_, _06688_, _06686_);
  or (_06690_, _06191_, _04571_);
  or (_06691_, _06182_, _04569_);
  and (_06692_, _06691_, _06196_);
  nand (_06693_, _06692_, _06690_);
  nand (_06694_, _06693_, _06689_);
  nand (_06695_, _06694_, _06202_);
  nand (_06696_, _06695_, _06685_);
  nand (_06697_, _06696_, _06165_);
  nand (_06698_, _06697_, _06675_);
  and (_06699_, _06698_, _06653_);
  or (_06700_, _06182_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_06701_, _06191_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_06702_, _06701_, _06190_);
  and (_06703_, _06702_, _06700_);
  or (_06704_, _06191_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_06705_, _06182_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_06706_, _06705_, _06196_);
  and (_06707_, _06706_, _06704_);
  nor (_06708_, _06707_, _06703_);
  nand (_06709_, _06708_, _06175_);
  or (_06710_, _06182_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_06711_, _06191_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_06712_, _06711_, _06190_);
  and (_06713_, _06712_, _06710_);
  or (_06714_, _06191_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_06715_, _06182_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_06716_, _06715_, _06196_);
  and (_06717_, _06716_, _06714_);
  nor (_06718_, _06717_, _06713_);
  nand (_06719_, _06718_, _06202_);
  nand (_06720_, _06719_, _06709_);
  nand (_06721_, _06720_, _06166_);
  or (_06722_, _06182_, _05000_);
  or (_06723_, _06191_, _04998_);
  and (_06724_, _06723_, _06190_);
  nand (_06725_, _06724_, _06722_);
  or (_06726_, _06191_, _05006_);
  or (_06727_, _06182_, _05004_);
  and (_06728_, _06727_, _06196_);
  nand (_06729_, _06728_, _06726_);
  nand (_06730_, _06729_, _06725_);
  nand (_06731_, _06730_, _06175_);
  or (_06732_, _06191_, _05018_);
  or (_06733_, _06182_, _05020_);
  and (_06734_, _06733_, _06190_);
  nand (_06735_, _06734_, _06732_);
  or (_06736_, _06191_, _05014_);
  or (_06737_, _06182_, _05012_);
  and (_06738_, _06737_, _06196_);
  nand (_06739_, _06738_, _06736_);
  nand (_06740_, _06739_, _06735_);
  nand (_06741_, _06740_, _06202_);
  nand (_06742_, _06741_, _06731_);
  nand (_06743_, _06742_, _06165_);
  nand (_06744_, _06743_, _06721_);
  or (_06745_, _06182_, \oc8051_golden_model_1.IRAM[9] [2]);
  or (_06746_, _06191_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_06747_, _06746_, _06190_);
  and (_06748_, _06747_, _06745_);
  or (_06749_, _06191_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_06750_, _06182_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_06751_, _06750_, _06196_);
  and (_06752_, _06751_, _06749_);
  nor (_06753_, _06752_, _06748_);
  nand (_06754_, _06753_, _06175_);
  or (_06755_, _06182_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_06756_, _06191_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_06757_, _06756_, _06190_);
  and (_06758_, _06757_, _06755_);
  or (_06759_, _06191_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_06760_, _06182_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_06761_, _06760_, _06196_);
  and (_06762_, _06761_, _06759_);
  nor (_06763_, _06762_, _06758_);
  nand (_06764_, _06763_, _06202_);
  nand (_06765_, _06764_, _06754_);
  nand (_06766_, _06765_, _06166_);
  or (_06767_, _06182_, _05186_);
  or (_06768_, _06191_, _05184_);
  and (_06769_, _06768_, _06190_);
  nand (_06770_, _06769_, _06767_);
  or (_06771_, _06191_, _05192_);
  or (_06772_, _06182_, _05190_);
  and (_06773_, _06772_, _06196_);
  nand (_06774_, _06773_, _06771_);
  nand (_06775_, _06774_, _06770_);
  nand (_06776_, _06775_, _06175_);
  or (_06777_, _06191_, _05204_);
  or (_06778_, _06182_, _05206_);
  and (_06779_, _06778_, _06190_);
  nand (_06780_, _06779_, _06777_);
  or (_06781_, _06191_, _05200_);
  or (_06782_, _06182_, _05198_);
  and (_06783_, _06782_, _06196_);
  nand (_06784_, _06783_, _06781_);
  nand (_06785_, _06784_, _06780_);
  nand (_06786_, _06785_, _06202_);
  nand (_06787_, _06786_, _06776_);
  nand (_06788_, _06787_, _06165_);
  nand (_06789_, _06788_, _06766_);
  and (_06790_, _06789_, _06744_);
  and (_06791_, _06790_, _06699_);
  or (_06792_, _06182_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_06793_, _06191_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_06794_, _06793_, _06190_);
  and (_06795_, _06794_, _06792_);
  or (_06796_, _06191_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_06797_, _06182_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_06798_, _06797_, _06196_);
  and (_06799_, _06798_, _06796_);
  nor (_06800_, _06799_, _06795_);
  nand (_06801_, _06800_, _06175_);
  or (_06802_, _06182_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_06803_, _06191_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_06804_, _06803_, _06190_);
  and (_06805_, _06804_, _06802_);
  or (_06806_, _06191_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_06807_, _06182_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_06808_, _06807_, _06196_);
  and (_06809_, _06808_, _06806_);
  nor (_06810_, _06809_, _06805_);
  nand (_06811_, _06810_, _06202_);
  nand (_06812_, _06811_, _06801_);
  nand (_06813_, _06812_, _06166_);
  or (_06814_, _06182_, _05749_);
  or (_06815_, _06191_, _05747_);
  and (_06816_, _06815_, _06190_);
  nand (_06817_, _06816_, _06814_);
  or (_06818_, _06191_, _05755_);
  or (_06819_, _06182_, _05753_);
  and (_06820_, _06819_, _06196_);
  nand (_06821_, _06820_, _06818_);
  nand (_06822_, _06821_, _06817_);
  nand (_06823_, _06822_, _06175_);
  or (_06824_, _06191_, _05767_);
  or (_06825_, _06182_, _05769_);
  and (_06826_, _06825_, _06190_);
  nand (_06827_, _06826_, _06824_);
  or (_06828_, _06191_, _05763_);
  or (_06829_, _06182_, _05761_);
  and (_06830_, _06829_, _06196_);
  nand (_06831_, _06830_, _06828_);
  nand (_06832_, _06831_, _06827_);
  nand (_06833_, _06832_, _06202_);
  nand (_06834_, _06833_, _06823_);
  nand (_06835_, _06834_, _06165_);
  nand (_06836_, _06835_, _06813_);
  or (_06837_, _06182_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_06838_, _06191_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_06839_, _06838_, _06190_);
  and (_06840_, _06839_, _06837_);
  or (_06841_, _06191_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_06842_, _06182_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_06843_, _06842_, _06196_);
  and (_06844_, _06843_, _06841_);
  nor (_06845_, _06844_, _06840_);
  nand (_06846_, _06845_, _06175_);
  or (_06847_, _06182_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_06848_, _06191_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_06849_, _06848_, _06190_);
  and (_06850_, _06849_, _06847_);
  or (_06851_, _06191_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_06852_, _06182_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_06853_, _06852_, _06196_);
  and (_06854_, _06853_, _06851_);
  nor (_06855_, _06854_, _06850_);
  nand (_06856_, _06855_, _06202_);
  nand (_06857_, _06856_, _06846_);
  nand (_06858_, _06857_, _06166_);
  or (_06859_, _06182_, _05848_);
  or (_06860_, _06191_, _05846_);
  and (_06861_, _06860_, _06190_);
  nand (_06862_, _06861_, _06859_);
  or (_06863_, _06191_, _05854_);
  or (_06864_, _06182_, _05852_);
  and (_06865_, _06864_, _06196_);
  nand (_06866_, _06865_, _06863_);
  nand (_06867_, _06866_, _06862_);
  nand (_06868_, _06867_, _06175_);
  or (_06869_, _06191_, _05866_);
  or (_06870_, _06182_, _05868_);
  and (_06871_, _06870_, _06190_);
  nand (_06872_, _06871_, _06869_);
  or (_06873_, _06191_, _05862_);
  or (_06874_, _06182_, _05860_);
  and (_06875_, _06874_, _06196_);
  nand (_06876_, _06875_, _06873_);
  nand (_06877_, _06876_, _06872_);
  nand (_06878_, _06877_, _06202_);
  nand (_06879_, _06878_, _06868_);
  nand (_06880_, _06879_, _06165_);
  nand (_06881_, _06880_, _06858_);
  and (_06882_, _06881_, _06836_);
  and (_06883_, _06882_, _06791_);
  and (_06884_, _06883_, _06607_);
  nor (_06885_, _06884_, _06280_);
  and (_06886_, _06884_, _06280_);
  or (_06887_, _06886_, _06885_);
  or (_06888_, _06887_, _04728_);
  and (_06889_, _06888_, _06562_);
  and (_06890_, _06889_, _06561_);
  and (_06891_, _06250_, _04726_);
  or (_06892_, _06891_, _03833_);
  or (_06893_, _06892_, _06890_);
  and (_06894_, _03134_, \oc8051_golden_model_1.PC [2]);
  and (_06895_, _06894_, \oc8051_golden_model_1.PC [3]);
  and (_06896_, _06895_, _06024_);
  and (_06897_, _06896_, \oc8051_golden_model_1.PC [7]);
  nor (_06898_, _06896_, \oc8051_golden_model_1.PC [7]);
  nor (_06899_, _06898_, _06897_);
  not (_06900_, _06899_);
  nand (_06901_, _06900_, _03833_);
  and (_06902_, _06901_, _06893_);
  or (_06903_, _06902_, _03400_);
  and (_06904_, _06273_, _03400_);
  nor (_06905_, _06904_, _03672_);
  nand (_06906_, _06905_, _06903_);
  nand (_06907_, _06119_, _03672_);
  and (_06908_, _04220_, _03398_);
  nor (_06909_, _04973_, _06908_);
  not (_06910_, _06909_);
  and (_06911_, _04671_, _03398_);
  nor (_06912_, _06911_, _06910_);
  and (_06913_, _06912_, _06907_);
  and (_06914_, _06913_, _06906_);
  and (_06915_, _04813_, _04608_);
  nor (_06916_, _05236_, _05050_);
  and (_06917_, _06916_, _06915_);
  nor (_06918_, _05898_, _05799_);
  and (_06919_, _06918_, _06917_);
  nor (_06920_, _06919_, _06129_);
  and (_06921_, _06013_, _05498_);
  nor (_06922_, _06013_, _05498_);
  nor (_06923_, _06922_, _06921_);
  not (_06924_, _06923_);
  and (_06925_, _06924_, _06919_);
  nor (_06926_, _06925_, _06920_);
  nor (_06927_, _06926_, _06912_);
  or (_06928_, _06927_, _06914_);
  nor (_06929_, _06928_, _04907_);
  and (_06930_, _06926_, _04907_);
  or (_06931_, _06930_, _04743_);
  or (_06932_, _06931_, _06929_);
  and (_06933_, _06606_, _06584_);
  and (_06934_, _06652_, _06629_);
  and (_06935_, _06697_, _06675_);
  and (_06936_, _06935_, _06934_);
  and (_06937_, _06743_, _06721_);
  and (_06938_, _06788_, _06766_);
  and (_06939_, _06938_, _06937_);
  and (_06940_, _06939_, _06936_);
  and (_06941_, _06835_, _06813_);
  and (_06942_, _06880_, _06858_);
  and (_06943_, _06942_, _06941_);
  and (_06944_, _06943_, _06940_);
  and (_06945_, _06944_, _06933_);
  nor (_06946_, _06945_, _06280_);
  and (_06947_, _06945_, _06280_);
  or (_06948_, _06947_, _06946_);
  or (_06949_, _06948_, _04744_);
  and (_06950_, _06949_, _04922_);
  and (_06951_, _06950_, _06932_);
  nor (_06952_, _06951_, _06022_);
  nor (_06953_, _06952_, _04994_);
  or (_06954_, _06953_, _05340_);
  and (_06955_, _06954_, _05339_);
  not (_06956_, _03833_);
  not (_06957_, \oc8051_golden_model_1.PC [15]);
  and (_06958_, _06897_, \oc8051_golden_model_1.PC [8]);
  and (_06959_, _06958_, \oc8051_golden_model_1.PC [9]);
  and (_06960_, _06959_, \oc8051_golden_model_1.PC [10]);
  and (_06961_, _06960_, \oc8051_golden_model_1.PC [11]);
  and (_06962_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and (_06963_, _06962_, _06961_);
  and (_06964_, _06963_, \oc8051_golden_model_1.PC [14]);
  and (_06965_, _06964_, _06957_);
  nor (_06966_, _06964_, _06957_);
  or (_06967_, _06966_, _06965_);
  or (_06968_, _06967_, _06956_);
  and (_06969_, _06026_, \oc8051_golden_model_1.PC [8]);
  and (_06970_, _06969_, \oc8051_golden_model_1.PC [9]);
  and (_06971_, _06970_, \oc8051_golden_model_1.PC [10]);
  and (_06972_, _06971_, \oc8051_golden_model_1.PC [11]);
  and (_06973_, _06972_, _06962_);
  and (_06974_, _06973_, \oc8051_golden_model_1.PC [14]);
  and (_06975_, _06974_, _06957_);
  nor (_06976_, _06974_, _06957_);
  or (_06977_, _06976_, _06975_);
  or (_06978_, _06977_, _03833_);
  and (_06979_, _06978_, _06968_);
  and (_06980_, _06979_, _05334_);
  and (_06981_, _06980_, _05337_);
  or (_40439_, _06981_, _06955_);
  not (_06982_, \oc8051_golden_model_1.B [7]);
  nor (_06983_, _42908_, _06982_);
  nor (_06984_, _05354_, _06982_);
  and (_06985_, _06523_, _05354_);
  or (_06986_, _06985_, _06984_);
  and (_06987_, _06986_, _03959_);
  not (_06988_, _05354_);
  nor (_06989_, _05498_, _06988_);
  or (_06990_, _06989_, _06984_);
  or (_06991_, _03867_, _03799_);
  nor (_06992_, _06991_, _03786_);
  nor (_06993_, _06992_, _03411_);
  nor (_06994_, _06993_, _04287_);
  or (_06995_, _06994_, _06990_);
  nor (_06996_, _06094_, _06982_);
  and (_06997_, _06119_, _06094_);
  or (_06998_, _06997_, _06996_);
  and (_06999_, _06998_, _03691_);
  and (_07000_, _06250_, _05354_);
  or (_07001_, _07000_, _06984_);
  or (_07002_, _07001_, _04630_);
  and (_07003_, _05354_, \oc8051_golden_model_1.ACC [7]);
  or (_07004_, _07003_, _06984_);
  and (_07005_, _07004_, _04615_);
  nor (_07006_, _04615_, _06982_);
  or (_07007_, _07006_, _03757_);
  or (_07008_, _07007_, _07005_);
  and (_07009_, _07008_, _03697_);
  and (_07010_, _07009_, _07002_);
  and (_07011_, _06127_, _06094_);
  or (_07012_, _07011_, _06996_);
  and (_07013_, _07012_, _03696_);
  or (_07014_, _07013_, _03755_);
  or (_07015_, _07014_, _07010_);
  or (_07016_, _06990_, _04537_);
  and (_07017_, _07016_, _07015_);
  or (_07018_, _07017_, _03750_);
  or (_07019_, _07004_, _03751_);
  and (_07020_, _07019_, _03692_);
  and (_07021_, _07020_, _07018_);
  or (_07022_, _07021_, _06999_);
  and (_07023_, _07022_, _03685_);
  and (_07024_, _03846_, _03783_);
  or (_07025_, _06996_, _06268_);
  and (_07026_, _07025_, _03684_);
  and (_07027_, _07026_, _07012_);
  or (_07028_, _07027_, _07024_);
  or (_07029_, _07028_, _07023_);
  not (_07030_, _07024_);
  and (_07031_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_07032_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_07033_, _07032_, _07031_);
  and (_07034_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_07035_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_07036_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_07037_, _07036_, _07035_);
  nor (_07038_, _07037_, _07033_);
  and (_07039_, _07038_, _07034_);
  nor (_07040_, _07039_, _07033_);
  and (_07041_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_07042_, _07041_, _07036_);
  and (_07043_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_07044_, _07043_, _07031_);
  nor (_07045_, _07044_, _07042_);
  not (_07046_, _07045_);
  nor (_07047_, _07046_, _07040_);
  and (_07048_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_07049_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_07050_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_07051_, _07050_, _07049_);
  nor (_07052_, _07050_, _07049_);
  nor (_07053_, _07052_, _07051_);
  and (_07054_, _07053_, _07048_);
  nor (_07055_, _07053_, _07048_);
  nor (_07056_, _07055_, _07054_);
  and (_07057_, _07046_, _07040_);
  nor (_07058_, _07057_, _07047_);
  and (_07059_, _07058_, _07056_);
  nor (_07060_, _07059_, _07047_);
  not (_07061_, _07036_);
  and (_07062_, _07041_, _07061_);
  and (_07063_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_07064_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_07065_, _07064_, _07049_);
  and (_07066_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_07067_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_07068_, _07067_, _07066_);
  nor (_07069_, _07068_, _07065_);
  and (_07070_, _07069_, _07063_);
  nor (_07071_, _07069_, _07063_);
  nor (_07072_, _07071_, _07070_);
  and (_07073_, _07072_, _07062_);
  nor (_07074_, _07072_, _07062_);
  nor (_07075_, _07074_, _07073_);
  not (_07076_, _07075_);
  nor (_07077_, _07076_, _07060_);
  and (_07078_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_07079_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_07080_, _07079_, _07078_);
  nor (_07081_, _07054_, _07051_);
  and (_07082_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_07083_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_07084_, _07083_, _07082_);
  nor (_07085_, _07083_, _07082_);
  nor (_07086_, _07085_, _07084_);
  not (_07087_, _07086_);
  nor (_07088_, _07087_, _07081_);
  and (_07089_, _07087_, _07081_);
  nor (_07090_, _07089_, _07088_);
  and (_07091_, _07090_, _07080_);
  nor (_07092_, _07090_, _07080_);
  nor (_07093_, _07092_, _07091_);
  and (_07094_, _07076_, _07060_);
  nor (_07095_, _07094_, _07077_);
  and (_07096_, _07095_, _07093_);
  nor (_07097_, _07096_, _07077_);
  nor (_07098_, _07070_, _07065_);
  and (_07099_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_07100_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_07101_, _07100_, _07099_);
  nor (_07102_, _07100_, _07099_);
  nor (_07103_, _07102_, _07101_);
  not (_07104_, _07103_);
  nor (_07105_, _07104_, _07098_);
  and (_07106_, _07104_, _07098_);
  nor (_07107_, _07106_, _07105_);
  and (_07108_, _07107_, _07084_);
  nor (_07109_, _07107_, _07084_);
  nor (_07110_, _07109_, _07108_);
  nor (_07111_, _07073_, _07042_);
  and (_07112_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_07113_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_07114_, _07113_, _07064_);
  nor (_07115_, _07113_, _07064_);
  nor (_07116_, _07115_, _07114_);
  and (_07117_, _07116_, _07112_);
  nor (_07118_, _07116_, _07112_);
  nor (_07119_, _07118_, _07117_);
  not (_07120_, _07119_);
  nor (_07121_, _07120_, _07111_);
  and (_07122_, _07120_, _07111_);
  nor (_07123_, _07122_, _07121_);
  and (_07124_, _07123_, _07110_);
  nor (_07125_, _07123_, _07110_);
  nor (_07126_, _07125_, _07124_);
  not (_07127_, _07126_);
  nor (_07128_, _07127_, _07097_);
  nor (_07129_, _07091_, _07088_);
  not (_07130_, _07129_);
  and (_07131_, _07127_, _07097_);
  nor (_07132_, _07131_, _07128_);
  and (_07133_, _07132_, _07130_);
  nor (_07134_, _07133_, _07128_);
  nor (_07135_, _07108_, _07105_);
  not (_07136_, _07135_);
  nor (_07137_, _07124_, _07121_);
  not (_07138_, _07137_);
  and (_07139_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_07140_, _07139_, _07064_);
  and (_07141_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_07142_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_07143_, _07142_, _07141_);
  nor (_07144_, _07143_, _07140_);
  nor (_07145_, _07117_, _07114_);
  and (_07146_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_07147_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_07148_, _07147_, _07146_);
  nor (_07149_, _07147_, _07146_);
  nor (_07150_, _07149_, _07148_);
  not (_07151_, _07150_);
  nor (_07152_, _07151_, _07145_);
  and (_07153_, _07151_, _07145_);
  nor (_07154_, _07153_, _07152_);
  and (_07155_, _07154_, _07101_);
  nor (_07156_, _07154_, _07101_);
  nor (_07157_, _07156_, _07155_);
  and (_07158_, _07157_, _07144_);
  nor (_07159_, _07157_, _07144_);
  nor (_07160_, _07159_, _07158_);
  and (_07161_, _07160_, _07138_);
  nor (_07162_, _07160_, _07138_);
  nor (_07163_, _07162_, _07161_);
  and (_07164_, _07163_, _07136_);
  nor (_07165_, _07163_, _07136_);
  nor (_07166_, _07165_, _07164_);
  not (_07167_, _07166_);
  nor (_07168_, _07167_, _07134_);
  nor (_07169_, _07164_, _07161_);
  nor (_07170_, _07155_, _07152_);
  not (_07171_, _07170_);
  and (_07172_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_07173_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_07174_, _07173_, _07172_);
  nor (_07175_, _07173_, _07172_);
  nor (_07176_, _07175_, _07174_);
  and (_07177_, _07176_, _07140_);
  nor (_07178_, _07176_, _07140_);
  nor (_07179_, _07178_, _07177_);
  and (_07180_, _07179_, _07148_);
  nor (_07181_, _07179_, _07148_);
  nor (_07182_, _07181_, _07180_);
  and (_07183_, _07182_, _07139_);
  nor (_07184_, _07182_, _07139_);
  nor (_07185_, _07184_, _07183_);
  and (_07186_, _07185_, _07158_);
  nor (_07187_, _07185_, _07158_);
  nor (_07188_, _07187_, _07186_);
  and (_07189_, _07188_, _07171_);
  nor (_07190_, _07188_, _07171_);
  nor (_07191_, _07190_, _07189_);
  not (_07192_, _07191_);
  nor (_07193_, _07192_, _07169_);
  and (_07194_, _07192_, _07169_);
  nor (_07195_, _07194_, _07193_);
  and (_07196_, _07195_, _07168_);
  nor (_07197_, _07189_, _07186_);
  nor (_07198_, _07180_, _07177_);
  not (_07199_, _07198_);
  and (_07200_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_07201_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_07202_, _07201_, _07200_);
  nor (_07203_, _07201_, _07200_);
  nor (_07204_, _07203_, _07202_);
  and (_07205_, _07204_, _07174_);
  nor (_07206_, _07204_, _07174_);
  nor (_07207_, _07206_, _07205_);
  and (_07208_, _07207_, _07183_);
  nor (_07209_, _07207_, _07183_);
  nor (_07210_, _07209_, _07208_);
  and (_07211_, _07210_, _07199_);
  nor (_07212_, _07210_, _07199_);
  nor (_07213_, _07212_, _07211_);
  not (_07214_, _07213_);
  nor (_07215_, _07214_, _07197_);
  and (_07216_, _07214_, _07197_);
  nor (_07217_, _07216_, _07215_);
  and (_07218_, _07217_, _07193_);
  nor (_07219_, _07217_, _07193_);
  nor (_07220_, _07219_, _07218_);
  and (_07221_, _07220_, _07196_);
  nor (_07222_, _07220_, _07196_);
  and (_07223_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_07224_, _07223_, _07036_);
  and (_07225_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_07226_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_07227_, _07226_, _07032_);
  nor (_07228_, _07227_, _07224_);
  and (_07229_, _07228_, _07225_);
  nor (_07230_, _07229_, _07224_);
  not (_07231_, _07230_);
  nor (_07232_, _07038_, _07034_);
  nor (_07233_, _07232_, _07039_);
  and (_07234_, _07233_, _07231_);
  and (_07235_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_07236_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_07237_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_07238_, _07237_, _07236_);
  nor (_07239_, _07237_, _07236_);
  nor (_07240_, _07239_, _07238_);
  and (_07241_, _07240_, _07235_);
  nor (_07242_, _07240_, _07235_);
  nor (_07243_, _07242_, _07241_);
  nor (_07244_, _07233_, _07231_);
  nor (_07245_, _07244_, _07234_);
  and (_07246_, _07245_, _07243_);
  nor (_07247_, _07246_, _07234_);
  nor (_07248_, _07058_, _07056_);
  nor (_07249_, _07248_, _07059_);
  not (_07250_, _07249_);
  nor (_07251_, _07250_, _07247_);
  and (_07252_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_07253_, _07252_, _07079_);
  nor (_07254_, _07241_, _07238_);
  nor (_07255_, _07079_, _07078_);
  nor (_07256_, _07255_, _07080_);
  not (_07257_, _07256_);
  nor (_07258_, _07257_, _07254_);
  and (_07259_, _07257_, _07254_);
  nor (_07260_, _07259_, _07258_);
  and (_07261_, _07260_, _07253_);
  nor (_07262_, _07260_, _07253_);
  nor (_07263_, _07262_, _07261_);
  and (_07264_, _07250_, _07247_);
  nor (_07265_, _07264_, _07251_);
  and (_07266_, _07265_, _07263_);
  nor (_07267_, _07266_, _07251_);
  nor (_07268_, _07095_, _07093_);
  nor (_07269_, _07268_, _07096_);
  not (_07270_, _07269_);
  nor (_07271_, _07270_, _07267_);
  nor (_07272_, _07261_, _07258_);
  not (_07273_, _07272_);
  and (_07274_, _07270_, _07267_);
  nor (_07275_, _07274_, _07271_);
  and (_07276_, _07275_, _07273_);
  nor (_07277_, _07276_, _07271_);
  nor (_07278_, _07132_, _07130_);
  nor (_07279_, _07278_, _07133_);
  not (_07280_, _07279_);
  nor (_07281_, _07280_, _07277_);
  and (_07282_, _07167_, _07134_);
  nor (_07283_, _07282_, _07168_);
  and (_07284_, _07283_, _07281_);
  nor (_07285_, _07195_, _07168_);
  nor (_07286_, _07285_, _07196_);
  nand (_07287_, _07286_, _07284_);
  and (_07288_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_07289_, _07288_, _07223_);
  and (_07290_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_07291_, _07288_, _07223_);
  nor (_07292_, _07291_, _07289_);
  and (_07293_, _07292_, _07290_);
  nor (_07294_, _07293_, _07289_);
  not (_07295_, _07294_);
  nor (_07296_, _07228_, _07225_);
  nor (_07297_, _07296_, _07229_);
  and (_07298_, _07297_, _07295_);
  and (_07299_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_07300_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_07301_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_07302_, _07301_, _07300_);
  nor (_07303_, _07301_, _07300_);
  nor (_07304_, _07303_, _07302_);
  and (_07305_, _07304_, _07299_);
  nor (_07306_, _07304_, _07299_);
  nor (_07307_, _07306_, _07305_);
  nor (_07308_, _07297_, _07295_);
  nor (_07309_, _07308_, _07298_);
  and (_07310_, _07309_, _07307_);
  nor (_07311_, _07310_, _07298_);
  not (_07312_, _07311_);
  nor (_07313_, _07245_, _07243_);
  nor (_07314_, _07313_, _07246_);
  and (_07315_, _07314_, _07312_);
  nor (_07316_, _07305_, _07302_);
  and (_07317_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_07318_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_07319_, _07318_, _07317_);
  nor (_07320_, _07319_, _07253_);
  not (_07321_, _07320_);
  nor (_07322_, _07321_, _07316_);
  and (_07323_, _07321_, _07316_);
  nor (_07324_, _07323_, _07322_);
  nor (_07325_, _07314_, _07312_);
  nor (_07326_, _07325_, _07315_);
  and (_07327_, _07326_, _07324_);
  nor (_07328_, _07327_, _07315_);
  nor (_07329_, _07265_, _07263_);
  nor (_07330_, _07329_, _07266_);
  not (_07331_, _07330_);
  nor (_07332_, _07331_, _07328_);
  and (_07333_, _07331_, _07328_);
  nor (_07334_, _07333_, _07332_);
  and (_07335_, _07334_, _07322_);
  nor (_07336_, _07335_, _07332_);
  nor (_07337_, _07275_, _07273_);
  nor (_07338_, _07337_, _07276_);
  not (_07339_, _07338_);
  nor (_07340_, _07339_, _07336_);
  and (_07341_, _07280_, _07277_);
  nor (_07342_, _07341_, _07281_);
  and (_07343_, _07342_, _07340_);
  nor (_07344_, _07283_, _07281_);
  nor (_07345_, _07344_, _07284_);
  and (_07346_, _07345_, _07343_);
  nor (_07347_, _07345_, _07343_);
  nor (_07348_, _07347_, _07346_);
  and (_07349_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_07350_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_07351_, _07350_, _07349_);
  and (_07352_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_07353_, _07350_, _07349_);
  nor (_07354_, _07353_, _07351_);
  and (_07355_, _07354_, _07352_);
  nor (_07356_, _07355_, _07351_);
  not (_07357_, _07356_);
  nor (_07358_, _07292_, _07290_);
  nor (_07359_, _07358_, _07293_);
  and (_07360_, _07359_, _07357_);
  and (_07361_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_07362_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_07363_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_07364_, _07363_, _07362_);
  nor (_07365_, _07363_, _07362_);
  nor (_07366_, _07365_, _07364_);
  and (_07367_, _07366_, _07361_);
  nor (_07368_, _07366_, _07361_);
  nor (_07369_, _07368_, _07367_);
  nor (_07370_, _07359_, _07357_);
  nor (_07371_, _07370_, _07360_);
  and (_07372_, _07371_, _07369_);
  nor (_07373_, _07372_, _07360_);
  not (_07374_, _07373_);
  nor (_07375_, _07309_, _07307_);
  nor (_07376_, _07375_, _07310_);
  and (_07377_, _07376_, _07374_);
  not (_07378_, _07252_);
  nor (_07379_, _07367_, _07364_);
  nor (_07380_, _07379_, _07378_);
  and (_07381_, _07379_, _07378_);
  nor (_07382_, _07381_, _07380_);
  nor (_07383_, _07376_, _07374_);
  nor (_07384_, _07383_, _07377_);
  and (_07385_, _07384_, _07382_);
  nor (_07386_, _07385_, _07377_);
  not (_07387_, _07386_);
  nor (_07388_, _07326_, _07324_);
  nor (_07389_, _07388_, _07327_);
  and (_07390_, _07389_, _07387_);
  nor (_07391_, _07389_, _07387_);
  nor (_07392_, _07391_, _07390_);
  and (_07393_, _07392_, _07380_);
  nor (_07394_, _07393_, _07390_);
  nor (_07395_, _07334_, _07322_);
  nor (_07396_, _07395_, _07335_);
  not (_07397_, _07396_);
  nor (_07398_, _07397_, _07394_);
  and (_07399_, _07339_, _07336_);
  nor (_07400_, _07399_, _07340_);
  and (_07401_, _07400_, _07398_);
  nor (_07402_, _07342_, _07340_);
  nor (_07403_, _07402_, _07343_);
  nand (_07404_, _07403_, _07401_);
  or (_07405_, _07403_, _07401_);
  and (_07406_, _07405_, _07404_);
  and (_07407_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_07408_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_07409_, _07408_, _07407_);
  and (_07410_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07411_, _07408_, _07407_);
  nor (_07412_, _07411_, _07409_);
  and (_07413_, _07412_, _07410_);
  nor (_07414_, _07413_, _07409_);
  not (_07415_, _07414_);
  nor (_07416_, _07354_, _07352_);
  nor (_07417_, _07416_, _07355_);
  and (_07418_, _07417_, _07415_);
  and (_07419_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_07420_, _07419_, _07363_);
  and (_07421_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_07422_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_07423_, _07422_, _07421_);
  nor (_07424_, _07423_, _07420_);
  nor (_07425_, _07417_, _07415_);
  nor (_07426_, _07425_, _07418_);
  and (_07427_, _07426_, _07424_);
  nor (_07428_, _07427_, _07418_);
  not (_07429_, _07428_);
  nor (_07430_, _07371_, _07369_);
  nor (_07431_, _07430_, _07372_);
  and (_07432_, _07431_, _07429_);
  nor (_07433_, _07431_, _07429_);
  nor (_07434_, _07433_, _07432_);
  and (_07435_, _07434_, _07420_);
  nor (_07436_, _07435_, _07432_);
  not (_07437_, _07436_);
  nor (_07438_, _07384_, _07382_);
  nor (_07439_, _07438_, _07385_);
  and (_07440_, _07439_, _07437_);
  nor (_07441_, _07392_, _07380_);
  nor (_07442_, _07441_, _07393_);
  and (_07443_, _07442_, _07440_);
  and (_07444_, _07397_, _07394_);
  nor (_07445_, _07444_, _07398_);
  and (_07446_, _07445_, _07443_);
  nor (_07447_, _07400_, _07398_);
  nor (_07448_, _07447_, _07401_);
  and (_07449_, _07448_, _07446_);
  nor (_07450_, _07448_, _07446_);
  nor (_07451_, _07450_, _07449_);
  and (_07452_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_07453_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_07454_, _07453_, _07452_);
  and (_07455_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_07456_, _07453_, _07452_);
  nor (_07457_, _07456_, _07454_);
  and (_07458_, _07457_, _07455_);
  nor (_07459_, _07458_, _07454_);
  not (_07460_, _07459_);
  nor (_07461_, _07412_, _07410_);
  nor (_07462_, _07461_, _07413_);
  and (_07463_, _07462_, _07460_);
  nor (_07464_, _07462_, _07460_);
  nor (_07465_, _07464_, _07463_);
  and (_07466_, _07465_, _07419_);
  nor (_07467_, _07466_, _07463_);
  not (_07468_, _07467_);
  nor (_07469_, _07426_, _07424_);
  nor (_07470_, _07469_, _07427_);
  and (_07471_, _07470_, _07468_);
  nor (_07472_, _07434_, _07420_);
  nor (_07473_, _07472_, _07435_);
  and (_07474_, _07473_, _07471_);
  nor (_07475_, _07439_, _07437_);
  nor (_07476_, _07475_, _07440_);
  and (_07477_, _07476_, _07474_);
  nor (_07478_, _07442_, _07440_);
  nor (_07479_, _07478_, _07443_);
  and (_07480_, _07479_, _07477_);
  nor (_07481_, _07445_, _07443_);
  nor (_07482_, _07481_, _07446_);
  and (_07483_, _07482_, _07480_);
  and (_07484_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_07485_, _07484_, _07453_);
  nor (_07486_, _07457_, _07455_);
  nor (_07487_, _07486_, _07458_);
  and (_07488_, _07487_, _07485_);
  nor (_07489_, _07465_, _07419_);
  nor (_07490_, _07489_, _07466_);
  and (_07491_, _07490_, _07488_);
  nor (_07492_, _07470_, _07468_);
  nor (_07493_, _07492_, _07471_);
  and (_07494_, _07493_, _07491_);
  nor (_07495_, _07473_, _07471_);
  nor (_07496_, _07495_, _07474_);
  and (_07497_, _07496_, _07494_);
  nor (_07498_, _07476_, _07474_);
  nor (_07499_, _07498_, _07477_);
  and (_07500_, _07499_, _07497_);
  nor (_07501_, _07479_, _07477_);
  nor (_07502_, _07501_, _07480_);
  and (_07503_, _07502_, _07500_);
  nor (_07504_, _07482_, _07480_);
  nor (_07505_, _07504_, _07483_);
  and (_07506_, _07505_, _07503_);
  nor (_07507_, _07506_, _07483_);
  not (_07508_, _07507_);
  and (_07509_, _07508_, _07451_);
  or (_07510_, _07509_, _07449_);
  nand (_07511_, _07510_, _07406_);
  and (_07512_, _07511_, _07404_);
  not (_07513_, _07512_);
  and (_07514_, _07513_, _07348_);
  or (_07515_, _07514_, _07346_);
  or (_07516_, _07286_, _07284_);
  and (_07517_, _07516_, _07287_);
  nand (_07518_, _07517_, _07515_);
  and (_07519_, _07518_, _07287_);
  nor (_07520_, _07519_, _07222_);
  or (_07521_, _07520_, _07221_);
  and (_07522_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_07523_, _07522_);
  nor (_07524_, _07523_, _07173_);
  nor (_07525_, _07524_, _07205_);
  nor (_07526_, _07211_, _07208_);
  nor (_07527_, _07526_, _07525_);
  and (_07528_, _07526_, _07525_);
  nor (_07529_, _07528_, _07527_);
  nor (_07530_, _07218_, _07215_);
  and (_07531_, _07530_, _07529_);
  nor (_07532_, _07530_, _07529_);
  or (_07533_, _07532_, _07531_);
  and (_07534_, _07533_, _07521_);
  and (_07535_, _07529_, _07215_);
  or (_07536_, _07527_, _07202_);
  or (_07537_, _07536_, _07535_);
  and (_07538_, _07529_, _07218_);
  or (_07539_, _07538_, _07537_);
  or (_07540_, _07539_, _07534_);
  or (_07541_, _07540_, _07030_);
  and (_07542_, _07541_, _03680_);
  and (_07543_, _07542_, _07029_);
  not (_07544_, _06994_);
  not (_07545_, _06094_);
  nor (_07546_, _06121_, _07545_);
  or (_07547_, _07546_, _06996_);
  and (_07548_, _07547_, _03679_);
  or (_07549_, _07548_, _07544_);
  or (_07550_, _07549_, _07543_);
  and (_07551_, _07550_, _06995_);
  or (_07552_, _07551_, _04678_);
  and (_07553_, _06237_, _05354_);
  or (_07554_, _06984_, _04679_);
  or (_07555_, _07554_, _07553_);
  and (_07556_, _07555_, _03415_);
  and (_07557_, _07556_, _07552_);
  and (_07558_, _03846_, _03410_);
  not (_07559_, _03415_);
  nor (_07560_, _06501_, _06988_);
  or (_07561_, _07560_, _06984_);
  and (_07562_, _07561_, _07559_);
  or (_07563_, _07562_, _07558_);
  or (_07564_, _07563_, _07557_);
  not (_07565_, _07558_);
  nor (_07566_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_07567_, _07566_, _07035_);
  not (_07568_, \oc8051_golden_model_1.B [1]);
  nor (_07569_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_07570_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and (_07571_, _07570_, _07569_);
  and (_07572_, _07571_, _07568_);
  nor (_07573_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and (_07574_, _07573_, _07572_);
  and (_07575_, \oc8051_golden_model_1.B [0], _06142_);
  not (_07576_, _07575_);
  and (_07577_, _07576_, _07574_);
  and (_07578_, _07577_, _07567_);
  nor (_07579_, _07574_, _06142_);
  not (_07580_, \oc8051_golden_model_1.B [2]);
  not (_07581_, \oc8051_golden_model_1.B [3]);
  nor (_07582_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_07583_, _07582_, _07569_);
  and (_07584_, _07583_, _07581_);
  and (_07585_, _07584_, _07580_);
  not (_07586_, \oc8051_golden_model_1.ACC [6]);
  and (_07587_, \oc8051_golden_model_1.B [0], _07586_);
  nor (_07588_, _07587_, _06142_);
  nor (_07589_, _07588_, _07568_);
  not (_07590_, _07589_);
  and (_07591_, _07590_, _07585_);
  not (_07592_, _07591_);
  and (_07593_, _07592_, _07579_);
  nor (_07594_, _07593_, _07578_);
  and (_07595_, _07591_, \oc8051_golden_model_1.B [0]);
  nor (_07596_, _07595_, _07586_);
  and (_07597_, _07596_, _07568_);
  nor (_07598_, _07596_, _07568_);
  nor (_07599_, _07598_, _07597_);
  nor (_07600_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_07601_, _07600_, _07223_);
  nor (_07602_, _07601_, \oc8051_golden_model_1.ACC [4]);
  nor (_07603_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  not (_07604_, \oc8051_golden_model_1.B [0]);
  and (_07605_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_07606_, _07605_, _07604_);
  nor (_07607_, _07606_, _07603_);
  nor (_07608_, _07607_, _07602_);
  not (_07609_, _07608_);
  and (_07610_, _07609_, _07599_);
  not (_07611_, _07610_);
  nor (_07612_, _07594_, \oc8051_golden_model_1.B [2]);
  nor (_07613_, _07612_, _07597_);
  and (_07614_, _07613_, _07611_);
  and (_07615_, \oc8051_golden_model_1.B [2], _06142_);
  nor (_07616_, _07615_, \oc8051_golden_model_1.B [7]);
  and (_07617_, _07616_, _07571_);
  not (_07618_, _07617_);
  nor (_07619_, _07618_, _07614_);
  nor (_07620_, _07619_, _07594_);
  nor (_07621_, _07620_, _07578_);
  and (_07622_, _07583_, \oc8051_golden_model_1.ACC [7]);
  nor (_07623_, _07622_, _07584_);
  nor (_07624_, _07609_, _07599_);
  nor (_07625_, _07624_, _07610_);
  not (_07626_, _07625_);
  and (_07627_, _07626_, _07619_);
  nor (_07628_, _07619_, _07596_);
  nor (_07629_, _07628_, _07627_);
  and (_07630_, _07629_, _07580_);
  nor (_07631_, _07629_, _07580_);
  nor (_07632_, _07631_, _07630_);
  not (_07633_, _07632_);
  not (_07634_, \oc8051_golden_model_1.ACC [5]);
  nor (_07635_, _07619_, _07634_);
  and (_07636_, _07619_, _07601_);
  or (_07637_, _07636_, _07635_);
  and (_07638_, _07637_, _07568_);
  nor (_07639_, _07637_, _07568_);
  not (_07640_, \oc8051_golden_model_1.ACC [4]);
  and (_07641_, \oc8051_golden_model_1.B [0], _07640_);
  nor (_07642_, _07641_, _07639_);
  nor (_07643_, _07642_, _07638_);
  nor (_07644_, _07643_, _07633_);
  nor (_07645_, _07621_, \oc8051_golden_model_1.B [3]);
  nor (_07646_, _07645_, _07630_);
  not (_07647_, _07646_);
  nor (_07648_, _07647_, _07644_);
  nor (_07649_, _07648_, _07623_);
  nor (_07650_, _07649_, _07621_);
  nor (_07651_, _07650_, _07578_);
  not (_07652_, _07649_);
  and (_07653_, _07643_, _07633_);
  nor (_07654_, _07653_, _07644_);
  nor (_07655_, _07654_, _07652_);
  nor (_07656_, _07649_, _07629_);
  nor (_07657_, _07656_, _07655_);
  and (_07658_, _07657_, _07581_);
  nor (_07659_, _07657_, _07581_);
  nor (_07660_, _07659_, _07658_);
  not (_07661_, _07660_);
  nor (_07662_, _07649_, _07637_);
  nor (_07663_, _07639_, _07638_);
  and (_07664_, _07663_, _07641_);
  nor (_07665_, _07663_, _07641_);
  nor (_07666_, _07665_, _07664_);
  and (_07667_, _07666_, _07649_);
  or (_07668_, _07667_, _07662_);
  nor (_07669_, _07668_, \oc8051_golden_model_1.B [2]);
  and (_07670_, _07668_, \oc8051_golden_model_1.B [2]);
  nor (_07671_, _07649_, _07640_);
  nor (_07672_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_07673_, _07672_, _07349_);
  and (_07674_, _07649_, _07673_);
  or (_07675_, _07674_, _07671_);
  and (_07676_, _07675_, _07568_);
  nor (_07677_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_07678_, _07677_, _07407_);
  nor (_07679_, _07678_, \oc8051_golden_model_1.ACC [2]);
  nor (_07680_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_07681_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_07682_, _07681_, _07604_);
  nor (_07683_, _07682_, _07680_);
  nor (_07684_, _07683_, _07679_);
  not (_07685_, _07684_);
  nor (_07686_, _07675_, _07568_);
  nor (_07687_, _07686_, _07676_);
  and (_07688_, _07687_, _07685_);
  nor (_07689_, _07688_, _07676_);
  nor (_07690_, _07689_, _07670_);
  nor (_07691_, _07690_, _07669_);
  nor (_07692_, _07691_, _07661_);
  nor (_07693_, _07651_, \oc8051_golden_model_1.B [4]);
  nor (_07694_, _07693_, _07658_);
  not (_07695_, _07694_);
  nor (_07696_, _07695_, _07692_);
  not (_07697_, \oc8051_golden_model_1.B [5]);
  and (_07698_, _07582_, _07697_);
  and (_07699_, \oc8051_golden_model_1.B [4], _06142_);
  not (_07700_, _07699_);
  and (_07701_, _07700_, _07698_);
  not (_07702_, _07701_);
  nor (_07703_, _07702_, _07696_);
  nor (_07704_, _07703_, _07651_);
  nor (_07705_, _07704_, _07578_);
  not (_07706_, \oc8051_golden_model_1.B [4]);
  and (_07707_, _07691_, _07661_);
  nor (_07708_, _07707_, _07692_);
  not (_07709_, _07708_);
  and (_07710_, _07709_, _07703_);
  nor (_07711_, _07703_, _07657_);
  nor (_07712_, _07711_, _07710_);
  and (_07713_, _07712_, _07706_);
  nor (_07714_, _07712_, _07706_);
  nor (_07715_, _07714_, _07713_);
  not (_07716_, _07715_);
  nor (_07717_, _07703_, _07668_);
  nor (_07718_, _07670_, _07669_);
  and (_07719_, _07718_, _07689_);
  nor (_07720_, _07718_, _07689_);
  nor (_07721_, _07720_, _07719_);
  not (_07722_, _07721_);
  and (_07723_, _07722_, _07703_);
  nor (_07724_, _07723_, _07717_);
  nor (_07725_, _07724_, \oc8051_golden_model_1.B [3]);
  and (_07726_, _07724_, \oc8051_golden_model_1.B [3]);
  nor (_07727_, _07687_, _07685_);
  nor (_07728_, _07727_, _07688_);
  not (_07729_, _07728_);
  and (_07730_, _07729_, _07703_);
  nor (_07731_, _07703_, _07675_);
  nor (_07732_, _07731_, _07730_);
  and (_07733_, _07732_, _07580_);
  not (_07734_, \oc8051_golden_model_1.ACC [3]);
  nor (_07735_, _07703_, _07734_);
  and (_07736_, _07703_, _07678_);
  or (_07737_, _07736_, _07735_);
  and (_07738_, _07737_, _07568_);
  nor (_07739_, _07737_, _07568_);
  not (_07740_, \oc8051_golden_model_1.ACC [2]);
  and (_07741_, \oc8051_golden_model_1.B [0], _07740_);
  nor (_07742_, _07741_, _07739_);
  nor (_07743_, _07742_, _07738_);
  nor (_07744_, _07732_, _07580_);
  nor (_07745_, _07744_, _07733_);
  not (_07746_, _07745_);
  nor (_07747_, _07746_, _07743_);
  nor (_07748_, _07747_, _07733_);
  nor (_07749_, _07748_, _07726_);
  nor (_07750_, _07749_, _07725_);
  nor (_07751_, _07750_, _07716_);
  nor (_07752_, _07705_, \oc8051_golden_model_1.B [5]);
  nor (_07753_, _07752_, _07713_);
  not (_07754_, _07753_);
  nor (_07755_, _07754_, _07751_);
  not (_07756_, _07755_);
  not (_07757_, _07582_);
  and (_07758_, \oc8051_golden_model_1.B [5], _06142_);
  nor (_07759_, _07758_, _07757_);
  and (_07760_, _07759_, _07756_);
  nor (_07761_, _07760_, _07705_);
  not (_07762_, _07760_);
  and (_07763_, _07750_, _07716_);
  nor (_07764_, _07763_, _07751_);
  nor (_07765_, _07764_, _07762_);
  nor (_07766_, _07760_, _07712_);
  nor (_07767_, _07766_, _07765_);
  and (_07768_, _07767_, _07697_);
  nor (_07769_, _07767_, _07697_);
  nor (_07770_, _07769_, _07768_);
  not (_07771_, _07770_);
  nor (_07772_, _07760_, _07724_);
  nor (_07773_, _07726_, _07725_);
  nor (_07774_, _07773_, _07748_);
  and (_07775_, _07773_, _07748_);
  or (_07776_, _07775_, _07774_);
  and (_07777_, _07776_, _07760_);
  or (_07778_, _07777_, _07772_);
  and (_07779_, _07778_, _07706_);
  nor (_07780_, _07778_, _07706_);
  and (_07781_, _07746_, _07743_);
  nor (_07782_, _07781_, _07747_);
  nor (_07783_, _07782_, _07762_);
  nor (_07784_, _07760_, _07732_);
  nor (_07785_, _07784_, _07783_);
  and (_07786_, _07785_, _07581_);
  nor (_07787_, _07739_, _07738_);
  nor (_07788_, _07787_, _07741_);
  and (_07789_, _07787_, _07741_);
  or (_07790_, _07789_, _07788_);
  nor (_07791_, _07790_, _07762_);
  nor (_07792_, _07760_, _07737_);
  nor (_07793_, _07792_, _07791_);
  and (_07794_, _07793_, _07580_);
  nor (_07795_, _07793_, _07580_);
  nor (_07796_, _07760_, _07740_);
  nor (_07797_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07798_, _07797_, _07452_);
  and (_07799_, _07760_, _07798_);
  or (_07800_, _07799_, _07796_);
  and (_07801_, _07800_, _07568_);
  and (_07802_, \oc8051_golden_model_1.B [0], _03491_);
  not (_07803_, _07802_);
  nor (_07804_, _07800_, _07568_);
  nor (_07805_, _07804_, _07801_);
  and (_07806_, _07805_, _07803_);
  nor (_07807_, _07806_, _07801_);
  nor (_07808_, _07807_, _07795_);
  nor (_07809_, _07808_, _07794_);
  nor (_07810_, _07785_, _07581_);
  nor (_07811_, _07810_, _07786_);
  not (_07812_, _07811_);
  nor (_07813_, _07812_, _07809_);
  nor (_07814_, _07813_, _07786_);
  nor (_07815_, _07814_, _07780_);
  nor (_07816_, _07815_, _07779_);
  nor (_07817_, _07816_, _07771_);
  nor (_07818_, _07817_, _07768_);
  and (_07819_, _06982_, \oc8051_golden_model_1.ACC [7]);
  nor (_07820_, _07819_, _07582_);
  nor (_07821_, _07820_, _07818_);
  nor (_07822_, _07761_, _07578_);
  nor (_07823_, _07822_, _07757_);
  nor (_07824_, _07823_, _07821_);
  and (_07825_, _07824_, _07761_);
  nor (_07826_, _07825_, _07578_);
  and (_07827_, _07826_, \oc8051_golden_model_1.B [7]);
  and (_07828_, _07826_, _06982_);
  nor (_07829_, _07828_, _07522_);
  not (_07830_, _07829_);
  not (_07831_, \oc8051_golden_model_1.B [6]);
  and (_07832_, _07816_, _07771_);
  nor (_07833_, _07832_, _07817_);
  nor (_07834_, _07833_, _07824_);
  not (_07835_, _07824_);
  nor (_07836_, _07835_, _07767_);
  nor (_07837_, _07836_, _07834_);
  nor (_07838_, _07837_, _07831_);
  and (_07839_, _07837_, _07831_);
  nor (_07840_, _07780_, _07779_);
  nor (_07841_, _07840_, _07814_);
  and (_07842_, _07840_, _07814_);
  or (_07843_, _07842_, _07841_);
  nor (_07844_, _07843_, _07824_);
  nor (_07845_, _07835_, _07778_);
  nor (_07846_, _07845_, _07844_);
  nor (_07847_, _07846_, _07697_);
  and (_07848_, _07846_, _07697_);
  not (_07849_, _07848_);
  and (_07850_, _07812_, _07809_);
  nor (_07851_, _07850_, _07813_);
  nor (_07852_, _07851_, _07824_);
  nor (_07853_, _07835_, _07785_);
  nor (_07854_, _07853_, _07852_);
  nor (_07855_, _07854_, _07706_);
  and (_07856_, _07824_, _07793_);
  nor (_07857_, _07795_, _07794_);
  and (_07858_, _07857_, _07807_);
  nor (_07859_, _07857_, _07807_);
  nor (_07860_, _07859_, _07858_);
  nor (_07861_, _07860_, _07824_);
  or (_07862_, _07861_, _07856_);
  and (_07863_, _07862_, _07581_);
  nor (_07864_, _07862_, _07581_);
  nor (_07865_, _07864_, _07863_);
  nor (_07866_, _07805_, _07803_);
  nor (_07867_, _07866_, _07806_);
  nor (_07868_, _07867_, _07824_);
  nor (_07869_, _07835_, _07800_);
  nor (_07870_, _07869_, _07868_);
  nor (_07871_, _07870_, _07580_);
  and (_07872_, _07870_, _07580_);
  nor (_07873_, _07872_, _07871_);
  and (_07874_, _07873_, _07865_);
  and (_07875_, _07824_, _03491_);
  and (_07876_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07877_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07878_, _07877_, _07876_);
  nor (_07879_, _07824_, _07878_);
  nor (_07880_, _07879_, _07875_);
  and (_07881_, _07880_, _07568_);
  nor (_07882_, _07880_, _07568_);
  and (_07883_, _07604_, \oc8051_golden_model_1.ACC [0]);
  not (_07884_, _07883_);
  nor (_07885_, _07884_, _07882_);
  nor (_07886_, _07885_, _07881_);
  and (_07887_, _07886_, _07874_);
  and (_07888_, _07871_, _07865_);
  nor (_07889_, _07888_, _07864_);
  not (_07890_, _07889_);
  nor (_07891_, _07890_, _07887_);
  and (_07892_, _07854_, _07706_);
  nor (_07893_, _07892_, _07891_);
  or (_07894_, _07893_, _07855_);
  and (_07895_, _07894_, _07849_);
  nor (_07896_, _07895_, _07847_);
  nor (_07897_, _07896_, _07839_);
  or (_07898_, _07897_, _07838_);
  and (_07899_, _07898_, _07830_);
  nor (_07900_, _07899_, _07827_);
  nor (_07901_, _07892_, _07855_);
  nor (_07902_, _07848_, _07847_);
  and (_07903_, _07902_, _07901_);
  nor (_07904_, _07839_, _07838_);
  and (_07905_, _07904_, _07830_);
  and (_07906_, _07905_, _07903_);
  nor (_07907_, _07882_, _07881_);
  and (_07908_, \oc8051_golden_model_1.B [0], _03558_);
  not (_07909_, _07908_);
  and (_07910_, _07909_, _07907_);
  and (_07911_, _07910_, _07884_);
  and (_07912_, _07911_, _07874_);
  and (_07913_, _07912_, _07906_);
  nor (_07914_, _07913_, _07900_);
  and (_07915_, _07914_, _07825_);
  or (_07916_, _07915_, _07578_);
  or (_07917_, _07916_, _07565_);
  and (_07918_, _07917_, _04694_);
  and (_07919_, _07918_, _07564_);
  and (_07920_, _06307_, _05354_);
  or (_07921_, _07920_, _06984_);
  and (_07922_, _07921_, _03839_);
  or (_07923_, _07922_, _03838_);
  or (_07924_, _07923_, _07919_);
  and (_07925_, _06515_, _05354_);
  or (_07926_, _07925_, _06984_);
  or (_07927_, _07926_, _04703_);
  and (_07928_, _07927_, _04701_);
  and (_07929_, _07928_, _07924_);
  or (_07930_, _07929_, _06987_);
  and (_07931_, _07930_, _04708_);
  or (_07932_, _06984_, _05501_);
  and (_07933_, _07921_, _03866_);
  and (_07934_, _07933_, _07932_);
  or (_07935_, _07934_, _07931_);
  and (_07936_, _07935_, _04706_);
  and (_07937_, _07004_, _03967_);
  and (_07938_, _07937_, _07932_);
  or (_07939_, _07938_, _03835_);
  or (_07940_, _07939_, _07936_);
  nor (_07941_, _06514_, _06988_);
  or (_07942_, _06984_, _06532_);
  or (_07943_, _07942_, _07941_);
  and (_07944_, _07943_, _06537_);
  and (_07945_, _07944_, _07940_);
  nor (_07946_, _06522_, _06988_);
  or (_07947_, _07946_, _06984_);
  and (_07948_, _07947_, _03954_);
  or (_07949_, _07948_, _03703_);
  or (_07950_, _07949_, _07945_);
  or (_07951_, _07001_, _03704_);
  and (_07952_, _07951_, _03385_);
  and (_07953_, _07952_, _07950_);
  and (_07954_, _06998_, _03384_);
  or (_07955_, _07954_, _03701_);
  or (_07956_, _07955_, _07953_);
  and (_07957_, _06021_, _05354_);
  or (_07958_, _06984_, _03702_);
  or (_07959_, _07958_, _07957_);
  and (_07960_, _07959_, _42908_);
  and (_07961_, _07960_, _07956_);
  or (_07962_, _07961_, _06983_);
  and (_40440_, _07962_, _41654_);
  nor (_07963_, _42908_, _06142_);
  and (_07964_, _03834_, _03393_);
  nand (_07965_, _07964_, _07586_);
  and (_07966_, _03853_, _03393_);
  and (_07967_, _06280_, _06142_);
  and (_07968_, _06237_, \oc8051_golden_model_1.ACC [7]);
  nor (_07969_, _07968_, _07967_);
  and (_07970_, _06933_, \oc8051_golden_model_1.ACC [6]);
  and (_07971_, _06607_, _07586_);
  nor (_07972_, _07971_, _07970_);
  and (_07973_, _06941_, \oc8051_golden_model_1.ACC [5]);
  and (_07974_, _06836_, _07634_);
  nor (_07975_, _07974_, _07973_);
  not (_07976_, _07975_);
  and (_07977_, _06942_, \oc8051_golden_model_1.ACC [4]);
  and (_07978_, _06881_, _07640_);
  nor (_07979_, _07978_, _07977_);
  and (_07980_, _06937_, \oc8051_golden_model_1.ACC [3]);
  and (_07981_, _06744_, _07734_);
  and (_07982_, _06938_, \oc8051_golden_model_1.ACC [2]);
  and (_07983_, _06789_, _07740_);
  nor (_07984_, _07983_, _07982_);
  not (_07985_, _07984_);
  and (_07986_, _06934_, \oc8051_golden_model_1.ACC [1]);
  and (_07987_, _06653_, _03491_);
  nor (_07988_, _07987_, _07986_);
  and (_07989_, _06935_, \oc8051_golden_model_1.ACC [0]);
  and (_07990_, _07989_, _07988_);
  nor (_07991_, _07990_, _07986_);
  nor (_07992_, _07991_, _07985_);
  nor (_07993_, _07992_, _07982_);
  nor (_07994_, _07993_, _07981_);
  or (_07995_, _07994_, _07980_);
  and (_07996_, _07995_, _07979_);
  nor (_07997_, _07996_, _07977_);
  nor (_07998_, _07997_, _07976_);
  or (_07999_, _07998_, _07973_);
  and (_08000_, _07999_, _07972_);
  nor (_08001_, _08000_, _07970_);
  nor (_08002_, _08001_, _07969_);
  and (_08003_, _08001_, _07969_);
  nor (_08004_, _08003_, _08002_);
  nand (_08005_, _08004_, _07966_);
  and (_08006_, _03473_, _03834_);
  not (_08007_, _08006_);
  and (_08008_, _06945_, \oc8051_golden_model_1.PSW [7]);
  nor (_08009_, _08008_, _06280_);
  and (_08010_, _08008_, _06280_);
  nor (_08011_, _08010_, _08009_);
  and (_08012_, _08011_, \oc8051_golden_model_1.ACC [7]);
  nor (_08013_, _08011_, \oc8051_golden_model_1.ACC [7]);
  nor (_08014_, _08013_, _08012_);
  and (_08015_, _06944_, \oc8051_golden_model_1.PSW [7]);
  nor (_08016_, _08015_, _06933_);
  nor (_08017_, _08016_, _08008_);
  and (_08018_, _08017_, \oc8051_golden_model_1.ACC [6]);
  nor (_08019_, _08017_, _07586_);
  and (_08020_, _08017_, _07586_);
  or (_08021_, _08020_, _08019_);
  and (_08022_, _06940_, _06942_);
  and (_08023_, _08022_, \oc8051_golden_model_1.PSW [7]);
  nor (_08024_, _08023_, _06941_);
  nor (_08025_, _08024_, _08015_);
  and (_08026_, _08025_, \oc8051_golden_model_1.ACC [5]);
  nor (_08027_, _08025_, _07634_);
  and (_08028_, _08025_, _07634_);
  nor (_08029_, _08028_, _08027_);
  and (_08030_, _06936_, \oc8051_golden_model_1.PSW [7]);
  and (_08031_, _08030_, _06939_);
  nor (_08032_, _08031_, _06942_);
  nor (_08033_, _08032_, _08023_);
  and (_08034_, _08033_, \oc8051_golden_model_1.ACC [4]);
  nor (_08035_, _08033_, _07640_);
  and (_08036_, _08033_, _07640_);
  or (_08037_, _08036_, _08035_);
  and (_08038_, _06936_, _06938_);
  and (_08039_, _08038_, \oc8051_golden_model_1.PSW [7]);
  nor (_08040_, _08039_, _06937_);
  nor (_08041_, _08040_, _08031_);
  and (_08042_, _08041_, \oc8051_golden_model_1.ACC [3]);
  nor (_08043_, _08041_, _07734_);
  and (_08044_, _08041_, _07734_);
  nor (_08045_, _08044_, _08043_);
  nor (_08046_, _08030_, _06938_);
  nor (_08047_, _08046_, _08039_);
  and (_08048_, _08047_, \oc8051_golden_model_1.ACC [2]);
  nor (_08049_, _08047_, _07740_);
  and (_08050_, _08047_, _07740_);
  nor (_08051_, _08050_, _08049_);
  and (_08052_, _06935_, \oc8051_golden_model_1.PSW [7]);
  nor (_08053_, _08052_, _06934_);
  nor (_08054_, _08053_, _08030_);
  and (_08055_, _08054_, \oc8051_golden_model_1.ACC [1]);
  and (_08056_, _08054_, _03491_);
  nor (_08057_, _08054_, _03491_);
  nor (_08058_, _08057_, _08056_);
  not (_08059_, \oc8051_golden_model_1.PSW [7]);
  and (_08060_, _06698_, _08059_);
  nor (_08061_, _08060_, _08052_);
  and (_08062_, _08061_, \oc8051_golden_model_1.ACC [0]);
  not (_08063_, _08062_);
  nor (_08064_, _08063_, _08058_);
  nor (_08065_, _08064_, _08055_);
  nor (_08066_, _08065_, _08051_);
  nor (_08067_, _08066_, _08048_);
  nor (_08068_, _08067_, _08045_);
  or (_08069_, _08068_, _08042_);
  and (_08070_, _08069_, _08037_);
  nor (_08071_, _08070_, _08034_);
  nor (_08072_, _08071_, _08029_);
  or (_08073_, _08072_, _08026_);
  and (_08074_, _08073_, _08021_);
  nor (_08075_, _08074_, _08018_);
  nor (_08076_, _08075_, _08014_);
  and (_08077_, _08075_, _08014_);
  nor (_08078_, _08077_, _08076_);
  and (_08079_, _03853_, _03473_);
  not (_08080_, _08079_);
  or (_08081_, _08080_, _08078_);
  and (_08082_, _05498_, _06142_);
  and (_08083_, _03480_, _03316_);
  nand (_08084_, _08083_, _08082_);
  and (_08085_, _03789_, _03476_);
  not (_08086_, _08085_);
  nor (_08087_, _03791_, _03786_);
  nor (_08088_, _08087_, _04346_);
  nor (_08089_, _03797_, _03799_);
  nor (_08090_, _08089_, _04346_);
  nor (_08091_, _08090_, _08088_);
  nor (_08092_, _05365_, _06142_);
  and (_08093_, _08092_, _03959_);
  not (_08094_, _05365_);
  nor (_08095_, _05498_, _08094_);
  nor (_08096_, _08095_, _08092_);
  nand (_08097_, _08096_, _07544_);
  and (_08098_, _03846_, _03689_);
  and (_08099_, _08098_, _07734_);
  nand (_08100_, _05498_, _04839_);
  nor (_08101_, _04957_, _04220_);
  nor (_08102_, _03413_, _03382_);
  nor (_08103_, _08102_, _03789_);
  and (_08104_, _08103_, _08101_);
  nor (_08105_, _08104_, _03449_);
  nand (_08106_, _08105_, _05498_);
  and (_08107_, _03846_, _04108_);
  not (_08108_, _08107_);
  nor (_08109_, _04234_, _06142_);
  and (_08110_, _04234_, _06142_);
  or (_08111_, _08110_, _08109_);
  or (_08112_, _08111_, _08105_);
  and (_08113_, _08112_, _08108_);
  and (_08114_, _08113_, _08106_);
  and (_08115_, _08107_, _06237_);
  or (_08116_, _08115_, _08114_);
  not (_08117_, _03450_);
  nor (_08118_, _03757_, _08117_);
  and (_08119_, _08118_, _08116_);
  and (_08120_, _03846_, _03695_);
  not (_08121_, _08092_);
  nand (_08122_, _06250_, _05365_);
  and (_08123_, _08122_, _08121_);
  nor (_08124_, _08123_, _04630_);
  or (_08125_, _08124_, _08120_);
  or (_08126_, _08125_, _08119_);
  nor (_08127_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_08128_, _08127_, _07734_);
  and (_08129_, _08128_, _07605_);
  and (_08130_, _08129_, \oc8051_golden_model_1.ACC [6]);
  and (_08131_, _08130_, \oc8051_golden_model_1.ACC [7]);
  nor (_08132_, _08130_, \oc8051_golden_model_1.ACC [7]);
  nor (_08133_, _08132_, _08131_);
  and (_08134_, _08128_, \oc8051_golden_model_1.ACC [4]);
  nor (_08135_, _08134_, \oc8051_golden_model_1.ACC [5]);
  nor (_08136_, _08135_, _08129_);
  nor (_08137_, _08129_, \oc8051_golden_model_1.ACC [6]);
  nor (_08138_, _08137_, _08130_);
  nor (_08139_, _08138_, _08136_);
  not (_08140_, _08139_);
  and (_08141_, _08140_, _08133_);
  nor (_08142_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_08143_, _08142_, _08139_);
  nor (_08144_, _08143_, _08133_);
  nor (_08145_, _08144_, _08141_);
  not (_08146_, _08145_);
  nand (_08147_, _08146_, _08120_);
  and (_08148_, _08147_, _03761_);
  and (_08149_, _08148_, _08126_);
  nor (_08150_, _06086_, _06142_);
  and (_08151_, _06127_, _06086_);
  nor (_08152_, _08151_, _08150_);
  nor (_08153_, _08152_, _03697_);
  nor (_08154_, _08096_, _04537_);
  or (_08155_, _08154_, _04839_);
  or (_08156_, _08155_, _08153_);
  or (_08157_, _08156_, _08149_);
  and (_08158_, _08157_, _08100_);
  or (_08159_, _08158_, _04645_);
  or (_08160_, _06237_, _04646_);
  and (_08161_, _08160_, _03751_);
  nand (_08162_, _08161_, _08159_);
  nor (_08163_, _05500_, _03751_);
  nor (_08164_, _08163_, _08098_);
  and (_08165_, _08164_, _08162_);
  or (_08166_, _08165_, _08099_);
  and (_08167_, _08166_, _03692_);
  and (_08168_, _06119_, _06086_);
  nor (_08169_, _08168_, _08150_);
  and (_08170_, _08169_, _03691_);
  or (_08171_, _08170_, _03684_);
  or (_08172_, _08171_, _08167_);
  and (_08173_, _08151_, _06268_);
  nor (_08174_, _08173_, _08150_);
  or (_08175_, _08174_, _03685_);
  and (_08176_, _08175_, _07030_);
  and (_08177_, _08176_, _08172_);
  nor (_08178_, _07502_, _07500_);
  nor (_08179_, _08178_, _07503_);
  nor (_08180_, _08179_, _07030_);
  nand (_08181_, _03416_, _03316_);
  not (_08182_, _08181_);
  or (_08183_, _08182_, _08180_);
  nor (_08184_, _08183_, _08177_);
  not (_08185_, _06013_);
  and (_08186_, _06919_, \oc8051_golden_model_1.PSW [7]);
  and (_08187_, _08186_, _08185_);
  nor (_08188_, _08187_, _05498_);
  and (_08189_, _08187_, _05498_);
  nor (_08190_, _08189_, _08188_);
  and (_08191_, _08190_, \oc8051_golden_model_1.ACC [7]);
  nor (_08192_, _08190_, \oc8051_golden_model_1.ACC [7]);
  nor (_08193_, _08192_, _08191_);
  not (_08194_, _08193_);
  nor (_08195_, _08186_, _08185_);
  nor (_08196_, _08195_, _08187_);
  nor (_08197_, _08196_, _07586_);
  not (_08198_, _05799_);
  not (_08199_, _05898_);
  and (_08200_, _06917_, _08199_);
  and (_08201_, _08200_, \oc8051_golden_model_1.PSW [7]);
  nor (_08202_, _08201_, _08198_);
  nor (_08203_, _08202_, _08186_);
  and (_08204_, _08203_, _07634_);
  nor (_08205_, _08203_, _07634_);
  nor (_08206_, _08205_, _08204_);
  not (_08207_, _08206_);
  and (_08208_, _06915_, \oc8051_golden_model_1.PSW [7]);
  and (_08209_, _08208_, _06916_);
  nor (_08210_, _08209_, _08199_);
  nor (_08211_, _08210_, _08201_);
  nor (_08212_, _08211_, _07640_);
  and (_08213_, _08211_, _07640_);
  or (_08214_, _08213_, _08212_);
  or (_08215_, _08214_, _08207_);
  not (_08216_, _05050_);
  not (_08217_, _05236_);
  and (_08218_, _06915_, _08217_);
  and (_08219_, _08218_, \oc8051_golden_model_1.PSW [7]);
  nor (_08220_, _08219_, _08216_);
  nor (_08221_, _08220_, _08209_);
  nor (_08222_, _08221_, _07734_);
  and (_08223_, _08221_, _07734_);
  nor (_08224_, _08223_, _08222_);
  nor (_08225_, _08208_, _08217_);
  nor (_08226_, _08225_, _08219_);
  nor (_08227_, _08226_, _07740_);
  and (_08228_, _08226_, _07740_);
  nor (_08229_, _08228_, _08227_);
  and (_08230_, _08229_, _08224_);
  and (_08231_, _04608_, \oc8051_golden_model_1.PSW [7]);
  nor (_08232_, _08231_, _04813_);
  nor (_08233_, _08232_, _08208_);
  and (_08234_, _08233_, _03491_);
  nor (_08235_, _08233_, _03491_);
  nor (_08236_, _04608_, \oc8051_golden_model_1.PSW [7]);
  nor (_08237_, _08236_, _08231_);
  and (_08238_, _08237_, _03558_);
  not (_08239_, _08238_);
  nor (_08240_, _08239_, _08235_);
  nor (_08241_, _08240_, _08234_);
  nand (_08242_, _08241_, _08230_);
  and (_08243_, _08227_, _08224_);
  nor (_08244_, _08243_, _08222_);
  and (_08245_, _08244_, _08242_);
  nor (_08246_, _08245_, _08215_);
  and (_08247_, _08212_, _08206_);
  nor (_08248_, _08247_, _08205_);
  not (_08249_, _08248_);
  nor (_08250_, _08249_, _08246_);
  and (_08251_, _08196_, _07586_);
  nor (_08252_, _08197_, _08251_);
  not (_08253_, _08252_);
  nor (_08254_, _08253_, _08250_);
  or (_08255_, _08254_, _08197_);
  nor (_08256_, _08255_, _08194_);
  and (_08257_, _08255_, _08194_);
  or (_08258_, _08257_, _08256_);
  nand (_08259_, _08258_, _08182_);
  and (_08260_, _03853_, _03416_);
  not (_08261_, _08260_);
  nand (_08262_, _08261_, _08259_);
  or (_08263_, _08262_, _08184_);
  not (_08264_, _08014_);
  nor (_08265_, _08035_, _08027_);
  or (_08266_, _08265_, _08028_);
  not (_08267_, _08029_);
  or (_08268_, _08037_, _08267_);
  and (_08269_, _08051_, _08045_);
  and (_08270_, _08061_, _03558_);
  nor (_08271_, _08270_, _08056_);
  or (_08272_, _08271_, _08057_);
  and (_08273_, _08272_, _08269_);
  and (_08274_, _08049_, _08045_);
  or (_08275_, _08274_, _08043_);
  nor (_08276_, _08275_, _08273_);
  or (_08277_, _08276_, _08268_);
  and (_08278_, _08277_, _08266_);
  nor (_08279_, _08278_, _08021_);
  or (_08280_, _08279_, _08019_);
  and (_08281_, _08280_, _08264_);
  nor (_08282_, _08280_, _08264_);
  nor (_08283_, _08282_, _08281_);
  nand (_08284_, _08283_, _08260_);
  and (_08285_, _08284_, _08263_);
  or (_08286_, _08285_, _03818_);
  and (_08287_, _03846_, _03416_);
  not (_08288_, _08287_);
  not (_08289_, _06015_);
  and (_08290_, _05902_, \oc8051_golden_model_1.PSW [7]);
  and (_08291_, _08290_, _08289_);
  nor (_08292_, _08291_, _05500_);
  and (_08293_, _08291_, _05500_);
  nor (_08294_, _08293_, _08292_);
  and (_08295_, _08294_, \oc8051_golden_model_1.ACC [7]);
  nor (_08296_, _08294_, \oc8051_golden_model_1.ACC [7]);
  nor (_08297_, _08296_, _08295_);
  not (_08298_, _08297_);
  nor (_08299_, _08290_, _08289_);
  nor (_08300_, _08299_, _08291_);
  nor (_08301_, _08300_, _07586_);
  not (_08302_, _05801_);
  not (_08303_, _05900_);
  and (_08304_, _05652_, \oc8051_golden_model_1.PSW [7]);
  and (_08305_, _08304_, _05603_);
  and (_08306_, _08305_, _05700_);
  and (_08307_, _08306_, _05554_);
  and (_08308_, _08307_, _08303_);
  nor (_08309_, _08308_, _08302_);
  nor (_08310_, _08309_, _08290_);
  and (_08311_, _08310_, _07634_);
  nor (_08312_, _08310_, _07634_);
  nor (_08313_, _08312_, _08311_);
  not (_08314_, _08313_);
  nor (_08315_, _08307_, _08303_);
  nor (_08316_, _08315_, _08308_);
  nor (_08317_, _08316_, _07640_);
  and (_08318_, _08316_, _07640_);
  or (_08319_, _08318_, _08317_);
  or (_08320_, _08319_, _08314_);
  nor (_08321_, _08306_, _05554_);
  nor (_08322_, _08321_, _08307_);
  nor (_08323_, _08322_, _07734_);
  and (_08324_, _08322_, _07734_);
  nor (_08325_, _08324_, _08323_);
  nor (_08326_, _08305_, _05700_);
  nor (_08327_, _08326_, _08306_);
  nor (_08328_, _08327_, _07740_);
  and (_08329_, _08327_, _07740_);
  nor (_08330_, _08329_, _08328_);
  and (_08331_, _08330_, _08325_);
  nor (_08332_, _08304_, _05603_);
  nor (_08333_, _08332_, _08305_);
  and (_08334_, _08333_, _03491_);
  nor (_08335_, _08333_, _03491_);
  nor (_08336_, _05652_, \oc8051_golden_model_1.PSW [7]);
  nor (_08337_, _08336_, _08304_);
  and (_08338_, _08337_, _03558_);
  not (_08339_, _08338_);
  nor (_08340_, _08339_, _08335_);
  nor (_08341_, _08340_, _08334_);
  nand (_08342_, _08341_, _08331_);
  and (_08343_, _08328_, _08325_);
  nor (_08344_, _08343_, _08323_);
  and (_08345_, _08344_, _08342_);
  nor (_08346_, _08345_, _08320_);
  and (_08347_, _08317_, _08313_);
  nor (_08348_, _08347_, _08312_);
  not (_08349_, _08348_);
  nor (_08350_, _08349_, _08346_);
  and (_08351_, _08300_, _07586_);
  nor (_08352_, _08301_, _08351_);
  not (_08353_, _08352_);
  nor (_08354_, _08353_, _08350_);
  or (_08355_, _08354_, _08301_);
  and (_08356_, _08355_, _08298_);
  nor (_08357_, _08355_, _08298_);
  nor (_08358_, _08357_, _08356_);
  nand (_08359_, _08358_, _03818_);
  and (_08360_, _08359_, _08288_);
  and (_08361_, _08360_, _08286_);
  and (_08362_, _05388_, \oc8051_golden_model_1.PSW [7]);
  and (_08363_, _08362_, _05402_);
  and (_08364_, _08363_, _05345_);
  and (_08365_, _08364_, _05165_);
  nor (_08366_, _08365_, _05351_);
  and (_08367_, _08365_, _05351_);
  nor (_08368_, _08367_, _08366_);
  and (_08369_, _08368_, \oc8051_golden_model_1.ACC [7]);
  nor (_08370_, _08368_, \oc8051_golden_model_1.ACC [7]);
  nor (_08371_, _08370_, _08369_);
  nor (_08372_, _08364_, _05165_);
  nor (_08373_, _08372_, _08365_);
  nor (_08374_, _08373_, _07586_);
  and (_08375_, _08363_, _05357_);
  nor (_08376_, _08375_, _05362_);
  nor (_08377_, _08376_, _08364_);
  and (_08378_, _08377_, _07634_);
  nor (_08379_, _08377_, _07634_);
  nor (_08380_, _08379_, _08378_);
  not (_08381_, _08380_);
  nor (_08382_, _08363_, _05357_);
  nor (_08383_, _08382_, _08375_);
  nor (_08384_, _08383_, _07640_);
  and (_08385_, _08383_, _07640_);
  or (_08386_, _08385_, _08384_);
  or (_08387_, _08386_, _08381_);
  nor (_08388_, _06120_, _03742_);
  nor (_08389_, _08388_, _08363_);
  nor (_08390_, _08389_, _07734_);
  and (_08391_, _08389_, _07734_);
  nor (_08392_, _08391_, _08390_);
  nor (_08393_, _08362_, _05174_);
  nor (_08394_, _08393_, _06120_);
  nor (_08395_, _08394_, _07740_);
  and (_08396_, _08394_, _07740_);
  nor (_08397_, _08396_, _08395_);
  and (_08398_, _08397_, _08392_);
  nor (_08399_, _04211_, _08059_);
  nor (_08400_, _08399_, _04750_);
  nor (_08401_, _08400_, _08362_);
  nor (_08402_, _08401_, _03491_);
  and (_08403_, _08401_, _03491_);
  and (_08404_, _04211_, _08059_);
  nor (_08405_, _08404_, _08399_);
  and (_08406_, _08405_, _03558_);
  nor (_08407_, _08406_, _08403_);
  or (_08408_, _08407_, _08402_);
  nand (_08409_, _08408_, _08398_);
  nor (_08410_, _08395_, _08390_);
  or (_08411_, _08410_, _08391_);
  and (_08412_, _08411_, _08409_);
  nor (_08413_, _08412_, _08387_);
  and (_08414_, _08384_, _08380_);
  nor (_08415_, _08414_, _08379_);
  not (_08416_, _08415_);
  nor (_08417_, _08416_, _08413_);
  and (_08418_, _08373_, _07586_);
  nor (_08419_, _08374_, _08418_);
  not (_08420_, _08419_);
  nor (_08421_, _08420_, _08417_);
  or (_08422_, _08421_, _08374_);
  nor (_08423_, _08422_, _08371_);
  and (_08424_, _08422_, _08371_);
  nor (_08425_, _08424_, _08423_);
  and (_08426_, _08425_, _08287_);
  or (_08427_, _08426_, _03547_);
  or (_08428_, _08427_, _08361_);
  or (_08429_, _03638_, _03422_);
  and (_08430_, _08429_, _03680_);
  and (_08431_, _08430_, _08428_);
  not (_08432_, _06086_);
  nor (_08433_, _06121_, _08432_);
  nor (_08434_, _08433_, _08150_);
  nor (_08435_, _08434_, _03680_);
  or (_08436_, _08435_, _07544_);
  or (_08437_, _08436_, _08431_);
  and (_08438_, _08437_, _08097_);
  or (_08439_, _08438_, _04678_);
  and (_08440_, _06237_, _05365_);
  nor (_08441_, _08440_, _08092_);
  nand (_08442_, _08441_, _04678_);
  and (_08443_, _08442_, _03415_);
  and (_08444_, _08443_, _08439_);
  nor (_08445_, _06501_, _08094_);
  nor (_08446_, _08445_, _08092_);
  nor (_08447_, _08446_, _03415_);
  or (_08448_, _08447_, _07558_);
  or (_08449_, _08448_, _08444_);
  or (_08450_, _07577_, _07565_);
  and (_08451_, _08450_, _08449_);
  or (_08452_, _08451_, _03466_);
  or (_08453_, _03638_, _03467_);
  and (_08454_, _08453_, _08452_);
  or (_08455_, _08454_, _03839_);
  and (_08456_, _03846_, _03482_);
  not (_08457_, _08456_);
  and (_08458_, _06307_, _05365_);
  nor (_08459_, _08458_, _08092_);
  nand (_08460_, _08459_, _03839_);
  and (_08461_, _08460_, _08457_);
  and (_08462_, _08461_, _08455_);
  and (_08463_, _08456_, _03638_);
  and (_08464_, _03485_, _03316_);
  or (_08465_, _08464_, _08463_);
  or (_08466_, _08465_, _08462_);
  nor (_08467_, _05498_, _06142_);
  nor (_08468_, _08467_, _08082_);
  not (_08469_, _08464_);
  or (_08470_, _08469_, _08468_);
  and (_08471_, _03853_, _03485_);
  not (_08472_, _08471_);
  and (_08473_, _08472_, _08470_);
  and (_08474_, _08473_, _08466_);
  and (_08475_, _08471_, _07969_);
  or (_08476_, _08475_, _03957_);
  or (_08477_, _08476_, _08474_);
  and (_08478_, _03846_, _03485_);
  not (_08479_, _08478_);
  or (_08480_, _06523_, _03958_);
  and (_08481_, _08480_, _08479_);
  and (_08482_, _08481_, _08477_);
  nor (_08483_, _03638_, \oc8051_golden_model_1.ACC [7]);
  and (_08484_, _03638_, \oc8051_golden_model_1.ACC [7]);
  nor (_08485_, _08484_, _08483_);
  and (_08486_, _08478_, _08485_);
  or (_08487_, _08486_, _03838_);
  or (_08488_, _08487_, _08482_);
  and (_08489_, _06515_, _05365_);
  nor (_08490_, _08489_, _08092_);
  nand (_08491_, _08490_, _03838_);
  and (_08492_, _08491_, _04701_);
  and (_08493_, _08492_, _08488_);
  or (_08494_, _08493_, _08093_);
  and (_08495_, _08494_, _08091_);
  not (_08496_, _08091_);
  and (_08497_, _08467_, _08496_);
  or (_08498_, _08497_, _08495_);
  and (_08499_, _08498_, _08086_);
  and (_08500_, _08467_, _08085_);
  or (_08501_, _08500_, _08499_);
  and (_08502_, _03853_, _03476_);
  not (_08503_, _08502_);
  and (_08504_, _08503_, _08501_);
  and (_08505_, _08502_, _07968_);
  or (_08506_, _08505_, _03965_);
  or (_08507_, _08506_, _08504_);
  and (_08508_, _03846_, _03476_);
  not (_08509_, _08508_);
  or (_08510_, _06521_, _03966_);
  and (_08511_, _08510_, _08509_);
  and (_08512_, _08511_, _08507_);
  and (_08513_, _08508_, _08484_);
  or (_08514_, _08513_, _08512_);
  and (_08515_, _08514_, _04708_);
  or (_08516_, _08459_, _06522_);
  nor (_08517_, _08516_, _04708_);
  or (_08518_, _08517_, _08083_);
  or (_08519_, _08518_, _08515_);
  and (_08520_, _08519_, _08084_);
  and (_08521_, _03853_, _03480_);
  or (_08522_, _08521_, _08520_);
  nand (_08523_, _08521_, _07967_);
  and (_08524_, _08523_, _03953_);
  and (_08525_, _08524_, _08522_);
  and (_08526_, _03846_, _03480_);
  nor (_08527_, _08526_, _03952_);
  not (_08528_, _08527_);
  not (_08529_, _08526_);
  nand (_08530_, _08529_, _06522_);
  and (_08531_, _08530_, _08528_);
  or (_08532_, _08531_, _08525_);
  nand (_08533_, _08526_, _08483_);
  and (_08534_, _08533_, _06532_);
  and (_08535_, _08534_, _08532_);
  nor (_08536_, _06514_, _08094_);
  nor (_08537_, _08536_, _08092_);
  nor (_08538_, _08537_, _06532_);
  not (_08539_, _03473_);
  nor (_08540_, _08089_, _08539_);
  nor (_08541_, _08087_, _08539_);
  nor (_08542_, _08541_, _08540_);
  not (_08543_, _08542_);
  or (_08544_, _08543_, _08538_);
  or (_08545_, _08544_, _08535_);
  not (_08546_, _04374_);
  and (_08547_, _08542_, _08546_);
  and (_08548_, _08196_, \oc8051_golden_model_1.ACC [6]);
  and (_08549_, _08203_, \oc8051_golden_model_1.ACC [5]);
  and (_08550_, _08211_, \oc8051_golden_model_1.ACC [4]);
  and (_08551_, _08221_, \oc8051_golden_model_1.ACC [3]);
  and (_08552_, _08226_, \oc8051_golden_model_1.ACC [2]);
  and (_08553_, _08233_, \oc8051_golden_model_1.ACC [1]);
  nor (_08554_, _08235_, _08234_);
  and (_08555_, _08237_, \oc8051_golden_model_1.ACC [0]);
  not (_08556_, _08555_);
  nor (_08557_, _08556_, _08554_);
  nor (_08558_, _08557_, _08553_);
  nor (_08559_, _08558_, _08229_);
  nor (_08560_, _08559_, _08552_);
  nor (_08561_, _08560_, _08224_);
  or (_08562_, _08561_, _08551_);
  and (_08563_, _08562_, _08214_);
  nor (_08564_, _08563_, _08550_);
  nor (_08565_, _08564_, _08206_);
  or (_08566_, _08565_, _08549_);
  and (_08567_, _08566_, _08253_);
  nor (_08568_, _08567_, _08548_);
  nor (_08569_, _08568_, _08193_);
  and (_08570_, _08568_, _08193_);
  nor (_08571_, _08570_, _08569_);
  and (_08572_, _08571_, _08546_);
  or (_08573_, _08572_, _08547_);
  and (_08574_, _08573_, _08545_);
  and (_08575_, _08571_, _04374_);
  or (_08576_, _08575_, _08079_);
  or (_08577_, _08576_, _08574_);
  and (_08578_, _08577_, _08081_);
  or (_08579_, _08578_, _03963_);
  and (_08580_, _03846_, _03473_);
  not (_08581_, _08580_);
  and (_08582_, _08300_, \oc8051_golden_model_1.ACC [6]);
  and (_08583_, _08310_, \oc8051_golden_model_1.ACC [5]);
  and (_08584_, _08316_, \oc8051_golden_model_1.ACC [4]);
  and (_08585_, _08322_, \oc8051_golden_model_1.ACC [3]);
  and (_08586_, _08327_, \oc8051_golden_model_1.ACC [2]);
  and (_08587_, _08333_, \oc8051_golden_model_1.ACC [1]);
  nor (_08588_, _08335_, _08334_);
  and (_08589_, _08337_, \oc8051_golden_model_1.ACC [0]);
  not (_08590_, _08589_);
  nor (_08591_, _08590_, _08588_);
  nor (_08592_, _08591_, _08587_);
  nor (_08593_, _08592_, _08330_);
  nor (_08594_, _08593_, _08586_);
  nor (_08595_, _08594_, _08325_);
  or (_08596_, _08595_, _08585_);
  and (_08597_, _08596_, _08319_);
  nor (_08598_, _08597_, _08584_);
  nor (_08599_, _08598_, _08313_);
  or (_08600_, _08599_, _08583_);
  and (_08601_, _08600_, _08353_);
  nor (_08602_, _08601_, _08582_);
  nor (_08603_, _08602_, _08297_);
  and (_08604_, _08602_, _08297_);
  nor (_08605_, _08604_, _08603_);
  or (_08606_, _08605_, _03964_);
  and (_08607_, _08606_, _08581_);
  and (_08608_, _08607_, _08579_);
  and (_08609_, _08373_, \oc8051_golden_model_1.ACC [6]);
  and (_08610_, _08377_, \oc8051_golden_model_1.ACC [5]);
  and (_08611_, _08383_, \oc8051_golden_model_1.ACC [4]);
  and (_08612_, _08389_, \oc8051_golden_model_1.ACC [3]);
  and (_08613_, _08394_, \oc8051_golden_model_1.ACC [2]);
  and (_08614_, _08401_, \oc8051_golden_model_1.ACC [1]);
  nor (_08615_, _08403_, _08402_);
  and (_08616_, _08405_, \oc8051_golden_model_1.ACC [0]);
  not (_08617_, _08616_);
  nor (_08618_, _08617_, _08615_);
  nor (_08619_, _08618_, _08614_);
  nor (_08620_, _08619_, _08397_);
  nor (_08621_, _08620_, _08613_);
  nor (_08622_, _08621_, _08392_);
  or (_08623_, _08622_, _08612_);
  and (_08624_, _08623_, _08386_);
  nor (_08625_, _08624_, _08611_);
  nor (_08626_, _08625_, _08380_);
  or (_08627_, _08626_, _08610_);
  and (_08628_, _08627_, _08420_);
  nor (_08629_, _08628_, _08609_);
  nor (_08630_, _08629_, _08371_);
  and (_08631_, _08629_, _08371_);
  nor (_08632_, _08631_, _08630_);
  and (_08633_, _08632_, _08580_);
  or (_08634_, _08633_, _08608_);
  and (_08635_, _08634_, _08007_);
  nand (_08636_, _08006_, \oc8051_golden_model_1.ACC [6]);
  and (_08637_, _03786_, _03393_);
  not (_08638_, _08637_);
  and (_08639_, _04671_, _03393_);
  nor (_08640_, _04220_, _03797_);
  and (_08641_, _08640_, _04291_);
  nor (_08642_, _08641_, _04389_);
  nor (_08643_, _08642_, _08639_);
  and (_08644_, _08643_, _08638_);
  nand (_08645_, _08644_, _08636_);
  or (_08646_, _08645_, _08635_);
  not (_08647_, _04392_);
  nor (_08648_, _06013_, _07586_);
  and (_08649_, _06013_, _07586_);
  nor (_08650_, _08648_, _08649_);
  nor (_08651_, _05799_, _07634_);
  and (_08652_, _05799_, _07634_);
  nor (_08653_, _08652_, _08651_);
  not (_08654_, _08653_);
  nor (_08655_, _05898_, _07640_);
  and (_08656_, _05898_, _07640_);
  nor (_08657_, _08655_, _08656_);
  nor (_08658_, _05050_, _07734_);
  and (_08659_, _05050_, _07734_);
  nor (_08660_, _05236_, _07740_);
  and (_08661_, _05236_, _07740_);
  nor (_08662_, _08660_, _08661_);
  not (_08663_, _08662_);
  and (_08664_, _04813_, \oc8051_golden_model_1.ACC [1]);
  and (_08665_, _04842_, _03491_);
  nor (_08666_, _08664_, _08665_);
  and (_08667_, _04608_, \oc8051_golden_model_1.ACC [0]);
  and (_08668_, _08667_, _08666_);
  nor (_08669_, _08668_, _08664_);
  nor (_08670_, _08669_, _08663_);
  nor (_08671_, _08670_, _08660_);
  nor (_08672_, _08671_, _08659_);
  or (_08673_, _08672_, _08658_);
  and (_08674_, _08673_, _08657_);
  nor (_08675_, _08674_, _08655_);
  nor (_08676_, _08675_, _08654_);
  or (_08677_, _08676_, _08651_);
  and (_08678_, _08677_, _08650_);
  nor (_08679_, _08678_, _08648_);
  nor (_08680_, _08679_, _08468_);
  and (_08681_, _08679_, _08468_);
  or (_08682_, _08681_, _08680_);
  or (_08683_, _08682_, _08644_);
  and (_08684_, _08683_, _08647_);
  and (_08685_, _08684_, _08646_);
  and (_08686_, _08682_, _04392_);
  or (_08687_, _08686_, _07966_);
  or (_08688_, _08687_, _08685_);
  and (_08689_, _08688_, _08005_);
  or (_08690_, _08689_, _03709_);
  and (_08691_, _03846_, _03393_);
  not (_08692_, _08691_);
  nor (_08693_, _06015_, _07586_);
  and (_08694_, _06015_, _07586_);
  nor (_08695_, _08694_, _08693_);
  nor (_08696_, _05801_, _07634_);
  and (_08697_, _05801_, _07634_);
  nor (_08698_, _05900_, _07640_);
  and (_08699_, _05900_, _07640_);
  nor (_08700_, _08699_, _08698_);
  and (_08701_, _05553_, _07734_);
  not (_08702_, _08701_);
  nor (_08703_, _05553_, _07734_);
  not (_08704_, _08703_);
  nor (_08705_, _05699_, _07740_);
  and (_08706_, _05699_, _07740_);
  nor (_08707_, _08706_, _08705_);
  not (_08708_, _08707_);
  nor (_08709_, _05602_, _03491_);
  and (_08710_, _05602_, _03491_);
  nor (_08711_, _08710_, _08709_);
  and (_08712_, _05652_, \oc8051_golden_model_1.ACC [0]);
  and (_08713_, _08712_, _08711_);
  nor (_08714_, _08713_, _08709_);
  nor (_08715_, _08714_, _08708_);
  nor (_08716_, _08715_, _08705_);
  nand (_08717_, _08716_, _08704_);
  and (_08718_, _08717_, _08702_);
  and (_08719_, _08718_, _08700_);
  nor (_08720_, _08719_, _08698_);
  nor (_08721_, _08720_, _08697_);
  or (_08722_, _08721_, _08696_);
  and (_08723_, _08722_, _08695_);
  nor (_08724_, _08723_, _08693_);
  nor (_08725_, _08724_, _06523_);
  and (_08726_, _08724_, _06523_);
  or (_08727_, _08726_, _08725_);
  or (_08728_, _08727_, _04166_);
  and (_08729_, _08728_, _08692_);
  and (_08730_, _08729_, _08690_);
  nor (_08731_, _03740_, _07586_);
  and (_08732_, _03740_, _07586_);
  nor (_08733_, _08731_, _08732_);
  nor (_08734_, _04034_, _07634_);
  and (_08735_, _04034_, _07634_);
  nor (_08736_, _08734_, _08735_);
  not (_08737_, _08736_);
  nor (_08738_, _04446_, _07640_);
  and (_08739_, _04446_, _07640_);
  nor (_08740_, _08738_, _08739_);
  nor (_08741_, _03669_, _07734_);
  and (_08742_, _03669_, _07734_);
  nor (_08743_, _04165_, _07740_);
  and (_08744_, _04165_, _07740_);
  nor (_08745_, _08743_, _08744_);
  not (_08746_, _08745_);
  nor (_08747_, _04482_, _03491_);
  nor (_08748_, _04211_, _03558_);
  not (_08749_, _08748_);
  and (_08750_, _04482_, _03491_);
  or (_08751_, _08750_, _08747_);
  nor (_08752_, _08751_, _08749_);
  nor (_08753_, _08752_, _08747_);
  nor (_08754_, _08753_, _08746_);
  nor (_08755_, _08754_, _08743_);
  nor (_08756_, _08755_, _08742_);
  or (_08757_, _08756_, _08741_);
  and (_08758_, _08757_, _08740_);
  nor (_08759_, _08758_, _08738_);
  nor (_08760_, _08759_, _08737_);
  or (_08761_, _08760_, _08734_);
  and (_08762_, _08761_, _08733_);
  nor (_08763_, _08762_, _08731_);
  nor (_08764_, _08763_, _08485_);
  and (_08765_, _08763_, _08485_);
  or (_08766_, _08765_, _08764_);
  and (_08767_, _08766_, _08691_);
  or (_08768_, _08767_, _07964_);
  or (_08769_, _08768_, _08730_);
  and (_08770_, _08769_, _07965_);
  or (_08771_, _08770_, _03703_);
  and (_08772_, _03846_, _03254_);
  not (_08773_, _08772_);
  nand (_08774_, _08123_, _03703_);
  and (_08775_, _08774_, _08773_);
  and (_08776_, _08775_, _08771_);
  and (_08777_, _03834_, _03254_);
  nor (_08778_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08779_, _08778_, _07680_);
  and (_08780_, _08779_, _07603_);
  and (_08781_, _08780_, _07586_);
  nor (_08782_, _08781_, _06142_);
  and (_08783_, _08781_, _06142_);
  nor (_08784_, _08783_, _08782_);
  nor (_08785_, _08784_, _08773_);
  or (_08786_, _08785_, _08777_);
  or (_08787_, _08786_, _08776_);
  nand (_08788_, _08777_, _08059_);
  and (_08789_, _08788_, _03385_);
  and (_08790_, _08789_, _08787_);
  nor (_08791_, _08169_, _03385_);
  or (_08792_, _08791_, _03701_);
  or (_08793_, _08792_, _08790_);
  and (_08794_, _03846_, _03398_);
  not (_08795_, _08794_);
  and (_08796_, _06021_, _05365_);
  nor (_08797_, _08796_, _08092_);
  nand (_08798_, _08797_, _03701_);
  and (_08799_, _08798_, _08795_);
  and (_08800_, _08799_, _08793_);
  and (_08801_, _03834_, _03398_);
  and (_08802_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08803_, _08802_, _07681_);
  nor (_08804_, _08803_, _07640_);
  and (_08805_, _08804_, \oc8051_golden_model_1.ACC [5]);
  and (_08806_, _08805_, \oc8051_golden_model_1.ACC [6]);
  nor (_08807_, _08806_, \oc8051_golden_model_1.ACC [7]);
  and (_08808_, _08806_, \oc8051_golden_model_1.ACC [7]);
  nor (_08809_, _08808_, _08807_);
  and (_08810_, _08809_, _08794_);
  or (_08811_, _08810_, _08801_);
  or (_08812_, _08811_, _08800_);
  nand (_08813_, _08801_, _03558_);
  and (_08814_, _08813_, _42908_);
  and (_08815_, _08814_, _08812_);
  or (_08816_, _08815_, _07963_);
  and (_40441_, _08816_, _41654_);
  not (_08817_, \oc8051_golden_model_1.SBUF [7]);
  nor (_08818_, _05396_, _08817_);
  and (_08819_, _06021_, _05396_);
  nor (_08820_, _08819_, _08818_);
  nor (_08821_, _08820_, _03702_);
  and (_08822_, _06523_, _05396_);
  nor (_08823_, _08822_, _08818_);
  nor (_08824_, _08823_, _04701_);
  and (_08825_, _06237_, _05396_);
  or (_08826_, _08825_, _08818_);
  and (_08827_, _08826_, _04678_);
  and (_08828_, _05396_, \oc8051_golden_model_1.ACC [7]);
  nor (_08829_, _08828_, _08818_);
  nor (_08830_, _08829_, _04616_);
  nor (_08831_, _04615_, _08817_);
  or (_08832_, _08831_, _08830_);
  and (_08833_, _08832_, _04630_);
  and (_08834_, _06250_, _05396_);
  nor (_08835_, _08834_, _08818_);
  nor (_08836_, _08835_, _04630_);
  or (_08837_, _08836_, _08833_);
  and (_08838_, _08837_, _04537_);
  not (_08839_, _05396_);
  nor (_08840_, _05498_, _08839_);
  nor (_08841_, _08840_, _08818_);
  nor (_08842_, _08841_, _04537_);
  nor (_08843_, _08842_, _08838_);
  nor (_08844_, _08843_, _03750_);
  nor (_08845_, _08829_, _03751_);
  nor (_08846_, _08845_, _07544_);
  not (_08847_, _08846_);
  nor (_08848_, _08847_, _08844_);
  and (_08849_, _08841_, _07544_);
  or (_08850_, _08849_, _04678_);
  nor (_08851_, _08850_, _08848_);
  or (_08852_, _08851_, _08827_);
  and (_08853_, _08852_, _03415_);
  not (_08854_, _03840_);
  nor (_08855_, _06501_, _08839_);
  nor (_08856_, _08855_, _08818_);
  nor (_08857_, _08856_, _03415_);
  or (_08858_, _08857_, _08854_);
  or (_08859_, _08858_, _08853_);
  and (_08860_, _06515_, _05396_);
  or (_08861_, _08818_, _04703_);
  nor (_08862_, _08861_, _08860_);
  and (_08863_, _06307_, _05396_);
  nor (_08864_, _08863_, _08818_);
  and (_08865_, _08864_, _03839_);
  or (_08866_, _08865_, _03959_);
  nor (_08867_, _08866_, _08862_);
  and (_08868_, _08867_, _08859_);
  nor (_08869_, _08868_, _08824_);
  nor (_08870_, _08869_, _03866_);
  nor (_08871_, _08818_, _05501_);
  not (_08872_, _08871_);
  nor (_08873_, _08864_, _04708_);
  and (_08874_, _08873_, _08872_);
  nor (_08875_, _08874_, _08870_);
  nor (_08876_, _08875_, _03967_);
  nor (_08877_, _08829_, _04706_);
  and (_08878_, _08877_, _08872_);
  or (_08879_, _08878_, _08876_);
  and (_08880_, _08879_, _06532_);
  nor (_08881_, _06514_, _08839_);
  nor (_08882_, _08881_, _08818_);
  nor (_08883_, _08882_, _06532_);
  or (_08884_, _08883_, _08880_);
  and (_08885_, _08884_, _06537_);
  nor (_08886_, _06522_, _08839_);
  nor (_08888_, _08886_, _08818_);
  nor (_08889_, _08888_, _06537_);
  or (_08890_, _08889_, _08885_);
  and (_08891_, _08890_, _03704_);
  nor (_08892_, _08835_, _03704_);
  or (_08893_, _08892_, _08891_);
  and (_08894_, _08893_, _03702_);
  nor (_08895_, _08894_, _08821_);
  nand (_08896_, _08895_, _42908_);
  or (_08897_, _42908_, \oc8051_golden_model_1.SBUF [7]);
  and (_08899_, _08897_, _41654_);
  and (_40443_, _08899_, _08896_);
  not (_08900_, \oc8051_golden_model_1.SCON [7]);
  nor (_08901_, _05406_, _08900_);
  and (_08902_, _06237_, _05406_);
  or (_08903_, _08902_, _08901_);
  and (_08904_, _08903_, _04678_);
  and (_08905_, _05406_, \oc8051_golden_model_1.ACC [7]);
  nor (_08906_, _08905_, _08901_);
  nor (_08907_, _08906_, _04616_);
  nor (_08909_, _04615_, _08900_);
  or (_08910_, _08909_, _08907_);
  and (_08911_, _08910_, _04630_);
  and (_08912_, _06250_, _05406_);
  nor (_08913_, _08912_, _08901_);
  nor (_08914_, _08913_, _04630_);
  or (_08915_, _08914_, _08911_);
  and (_08916_, _08915_, _03697_);
  nor (_08917_, _06099_, _08900_);
  and (_08918_, _06127_, _06099_);
  nor (_08920_, _08918_, _08917_);
  nor (_08921_, _08920_, _03697_);
  or (_08922_, _08921_, _03755_);
  or (_08923_, _08922_, _08916_);
  not (_08924_, _05406_);
  nor (_08925_, _05498_, _08924_);
  nor (_08926_, _08925_, _08901_);
  nand (_08927_, _08926_, _03755_);
  and (_08928_, _08927_, _08923_);
  and (_08929_, _08928_, _03751_);
  nor (_08931_, _08906_, _03751_);
  or (_08932_, _08931_, _08929_);
  and (_08933_, _08932_, _03692_);
  and (_08934_, _06119_, _06099_);
  nor (_08935_, _08934_, _08917_);
  nor (_08936_, _08935_, _03692_);
  or (_08937_, _08936_, _03684_);
  or (_08938_, _08937_, _08933_);
  nor (_08939_, _08917_, _06268_);
  nor (_08940_, _08939_, _08920_);
  or (_08942_, _08940_, _03685_);
  and (_08943_, _08942_, _03680_);
  and (_08944_, _08943_, _08938_);
  not (_08945_, _06099_);
  nor (_08946_, _06121_, _08945_);
  nor (_08947_, _08946_, _08917_);
  nor (_08948_, _08947_, _03680_);
  nor (_08949_, _08948_, _07544_);
  not (_08950_, _08949_);
  nor (_08951_, _08950_, _08944_);
  and (_08953_, _08926_, _07544_);
  or (_08954_, _08953_, _04678_);
  nor (_08955_, _08954_, _08951_);
  or (_08956_, _08955_, _08904_);
  and (_08957_, _08956_, _03415_);
  nor (_08958_, _06501_, _08924_);
  nor (_08959_, _08958_, _08901_);
  nor (_08960_, _08959_, _03415_);
  or (_08961_, _08960_, _08854_);
  or (_08962_, _08961_, _08957_);
  and (_08963_, _06515_, _05406_);
  or (_08964_, _08901_, _04703_);
  or (_08965_, _08964_, _08963_);
  and (_08966_, _06307_, _05406_);
  nor (_08967_, _08966_, _08901_);
  and (_08968_, _08967_, _03839_);
  nor (_08969_, _08968_, _03959_);
  and (_08970_, _08969_, _08965_);
  and (_08971_, _08970_, _08962_);
  and (_08972_, _06523_, _05406_);
  nor (_08973_, _08972_, _08901_);
  nor (_08974_, _08973_, _04701_);
  nor (_08975_, _08974_, _08971_);
  nor (_08976_, _08975_, _03866_);
  nor (_08977_, _08901_, _05501_);
  not (_08978_, _08977_);
  nor (_08979_, _08967_, _04708_);
  and (_08980_, _08979_, _08978_);
  nor (_08981_, _08980_, _08976_);
  nor (_08982_, _08981_, _03967_);
  nor (_08983_, _08906_, _04706_);
  and (_08984_, _08983_, _08978_);
  or (_08985_, _08984_, _08982_);
  and (_08986_, _08985_, _06532_);
  nor (_08987_, _06514_, _08924_);
  nor (_08988_, _08987_, _08901_);
  nor (_08989_, _08988_, _06532_);
  or (_08990_, _08989_, _08986_);
  and (_08991_, _08990_, _06537_);
  nor (_08992_, _06522_, _08924_);
  nor (_08993_, _08992_, _08901_);
  nor (_08994_, _08993_, _06537_);
  or (_08995_, _08994_, _08991_);
  and (_08996_, _08995_, _03704_);
  nor (_08997_, _08913_, _03704_);
  or (_08998_, _08997_, _08996_);
  and (_08999_, _08998_, _03385_);
  nor (_09000_, _08935_, _03385_);
  or (_09001_, _09000_, _08999_);
  and (_09002_, _09001_, _03702_);
  and (_09003_, _06021_, _05406_);
  nor (_09004_, _09003_, _08901_);
  nor (_09005_, _09004_, _03702_);
  or (_09006_, _09005_, _09002_);
  or (_09007_, _09006_, _42912_);
  or (_09008_, _42908_, \oc8051_golden_model_1.SCON [7]);
  and (_09009_, _09008_, _41654_);
  and (_40444_, _09009_, _09007_);
  not (_09010_, \oc8051_golden_model_1.PCON [7]);
  nor (_09011_, _05391_, _09010_);
  and (_09012_, _06021_, _05391_);
  nor (_09013_, _09012_, _09011_);
  nor (_09014_, _09013_, _03702_);
  and (_09015_, _06523_, _05391_);
  nor (_09016_, _09015_, _09011_);
  nor (_09017_, _09016_, _04701_);
  and (_09018_, _06237_, _05391_);
  or (_09019_, _09018_, _09011_);
  and (_09020_, _09019_, _04678_);
  and (_09021_, _05391_, \oc8051_golden_model_1.ACC [7]);
  nor (_09022_, _09021_, _09011_);
  nor (_09023_, _09022_, _04616_);
  nor (_09024_, _04615_, _09010_);
  or (_09025_, _09024_, _09023_);
  and (_09026_, _09025_, _04630_);
  and (_09027_, _06250_, _05391_);
  nor (_09028_, _09027_, _09011_);
  nor (_09029_, _09028_, _04630_);
  or (_09030_, _09029_, _09026_);
  and (_09031_, _09030_, _04537_);
  not (_09032_, _05391_);
  nor (_09033_, _05498_, _09032_);
  nor (_09034_, _09033_, _09011_);
  nor (_09035_, _09034_, _04537_);
  nor (_09036_, _09035_, _09031_);
  nor (_09037_, _09036_, _03750_);
  nor (_09038_, _09022_, _03751_);
  nor (_09039_, _09038_, _07544_);
  not (_09040_, _09039_);
  nor (_09041_, _09040_, _09037_);
  and (_09042_, _09034_, _07544_);
  or (_09043_, _09042_, _04678_);
  nor (_09044_, _09043_, _09041_);
  or (_09045_, _09044_, _09020_);
  and (_09046_, _09045_, _03415_);
  nor (_09047_, _06501_, _09032_);
  nor (_09048_, _09047_, _09011_);
  nor (_09049_, _09048_, _03415_);
  or (_09050_, _09049_, _08854_);
  or (_09051_, _09050_, _09046_);
  and (_09052_, _06515_, _05391_);
  or (_09053_, _09011_, _04703_);
  nor (_09054_, _09053_, _09052_);
  and (_09055_, _06307_, _05391_);
  nor (_09056_, _09055_, _09011_);
  and (_09057_, _09056_, _03839_);
  or (_09058_, _09057_, _03959_);
  nor (_09059_, _09058_, _09054_);
  and (_09060_, _09059_, _09051_);
  nor (_09061_, _09060_, _09017_);
  nor (_09062_, _09061_, _03866_);
  nor (_09063_, _09011_, _05501_);
  not (_09064_, _09063_);
  nor (_09065_, _09056_, _04708_);
  and (_09066_, _09065_, _09064_);
  nor (_09067_, _09066_, _09062_);
  nor (_09068_, _09067_, _03967_);
  nor (_09069_, _09022_, _04706_);
  and (_09070_, _09069_, _09064_);
  or (_09071_, _09070_, _09068_);
  and (_09072_, _09071_, _06532_);
  nor (_09073_, _06514_, _09032_);
  nor (_09074_, _09073_, _09011_);
  nor (_09075_, _09074_, _06532_);
  or (_09076_, _09075_, _09072_);
  and (_09077_, _09076_, _06537_);
  nor (_09078_, _06522_, _09032_);
  nor (_09079_, _09078_, _09011_);
  nor (_09080_, _09079_, _06537_);
  or (_09081_, _09080_, _09077_);
  and (_09082_, _09081_, _03704_);
  nor (_09083_, _09028_, _03704_);
  or (_09084_, _09083_, _09082_);
  and (_09085_, _09084_, _03702_);
  nor (_09086_, _09085_, _09014_);
  nand (_09087_, _09086_, _42908_);
  or (_09088_, _42908_, \oc8051_golden_model_1.PCON [7]);
  and (_09089_, _09088_, _41654_);
  and (_40445_, _09089_, _09087_);
  not (_09090_, _05438_);
  and (_09091_, _09090_, \oc8051_golden_model_1.TCON [7]);
  and (_09092_, _06250_, _05438_);
  or (_09093_, _09092_, _09091_);
  or (_09094_, _09093_, _04630_);
  and (_09095_, _05438_, \oc8051_golden_model_1.ACC [7]);
  or (_09096_, _09095_, _09091_);
  and (_09097_, _09096_, _04615_);
  and (_09098_, _04616_, \oc8051_golden_model_1.TCON [7]);
  or (_09099_, _09098_, _03757_);
  or (_09100_, _09099_, _09097_);
  and (_09101_, _09100_, _03697_);
  and (_09102_, _09101_, _09094_);
  not (_09103_, _06081_);
  and (_09104_, _09103_, \oc8051_golden_model_1.TCON [7]);
  and (_09105_, _06127_, _06081_);
  or (_09106_, _09105_, _09104_);
  and (_09107_, _09106_, _03696_);
  or (_09108_, _09107_, _03755_);
  or (_09109_, _09108_, _09102_);
  nor (_09110_, _05498_, _09090_);
  or (_09111_, _09110_, _09091_);
  or (_09112_, _09111_, _04537_);
  and (_09113_, _09112_, _09109_);
  or (_09114_, _09113_, _03750_);
  or (_09115_, _09096_, _03751_);
  and (_09116_, _09115_, _03692_);
  and (_09117_, _09116_, _09114_);
  and (_09118_, _06119_, _06081_);
  or (_09119_, _09118_, _09104_);
  and (_09120_, _09119_, _03691_);
  or (_09121_, _09120_, _03684_);
  or (_09122_, _09121_, _09117_);
  or (_09123_, _09104_, _06268_);
  and (_09124_, _09123_, _09106_);
  or (_09125_, _09124_, _03685_);
  and (_09126_, _09125_, _03680_);
  and (_09127_, _09126_, _09122_);
  nor (_09128_, _06121_, _09103_);
  or (_09129_, _09128_, _09104_);
  and (_09130_, _09129_, _03679_);
  or (_09131_, _09130_, _07544_);
  or (_09132_, _09131_, _09127_);
  or (_09133_, _09111_, _06994_);
  and (_09134_, _09133_, _09132_);
  or (_09135_, _09134_, _04678_);
  and (_09136_, _06237_, _05438_);
  or (_09137_, _09091_, _04679_);
  or (_09138_, _09137_, _09136_);
  and (_09139_, _09138_, _03415_);
  and (_09140_, _09139_, _09135_);
  nor (_09141_, _06501_, _09090_);
  or (_09142_, _09141_, _09091_);
  and (_09143_, _09142_, _07559_);
  or (_09144_, _09143_, _08854_);
  or (_09145_, _09144_, _09140_);
  and (_09146_, _06515_, _05438_);
  or (_09147_, _09091_, _04703_);
  or (_09148_, _09147_, _09146_);
  and (_09149_, _06307_, _05438_);
  or (_09150_, _09149_, _09091_);
  or (_09151_, _09150_, _04694_);
  and (_09152_, _09151_, _04701_);
  and (_09153_, _09152_, _09148_);
  and (_09154_, _09153_, _09145_);
  and (_09155_, _06523_, _05438_);
  or (_09156_, _09155_, _09091_);
  and (_09157_, _09156_, _03959_);
  or (_09158_, _09157_, _09154_);
  and (_09159_, _09158_, _04708_);
  or (_09160_, _09091_, _05501_);
  and (_09161_, _09150_, _03866_);
  and (_09162_, _09161_, _09160_);
  or (_09163_, _09162_, _09159_);
  and (_09164_, _09163_, _04706_);
  and (_09165_, _09096_, _03967_);
  and (_09166_, _09165_, _09160_);
  or (_09167_, _09166_, _03835_);
  or (_09168_, _09167_, _09164_);
  nor (_09169_, _06514_, _09090_);
  or (_09170_, _09091_, _06532_);
  or (_09171_, _09170_, _09169_);
  and (_09172_, _09171_, _06537_);
  and (_09173_, _09172_, _09168_);
  nor (_09174_, _06522_, _09090_);
  or (_09175_, _09174_, _09091_);
  and (_09176_, _09175_, _03954_);
  or (_09177_, _09176_, _03703_);
  or (_09178_, _09177_, _09173_);
  or (_09179_, _09093_, _03704_);
  and (_09180_, _09179_, _03385_);
  and (_09181_, _09180_, _09178_);
  and (_09182_, _09119_, _03384_);
  or (_09183_, _09182_, _03701_);
  or (_09184_, _09183_, _09181_);
  and (_09185_, _06021_, _05438_);
  or (_09186_, _09185_, _09091_);
  or (_09187_, _09186_, _03702_);
  and (_09188_, _09187_, _09184_);
  or (_09189_, _09188_, _42912_);
  or (_09190_, _42908_, \oc8051_golden_model_1.TCON [7]);
  and (_09191_, _09190_, _41654_);
  and (_40446_, _09191_, _09189_);
  not (_09192_, \oc8051_golden_model_1.TL0 [7]);
  nor (_09193_, _05411_, _09192_);
  and (_09194_, _06021_, _05411_);
  nor (_09195_, _09194_, _09193_);
  nor (_09196_, _09195_, _03702_);
  and (_09197_, _06523_, _05411_);
  nor (_09198_, _09197_, _09193_);
  nor (_09199_, _09198_, _04701_);
  and (_09200_, _06237_, _05411_);
  or (_09201_, _09200_, _09193_);
  and (_09202_, _09201_, _04678_);
  and (_09203_, _05411_, \oc8051_golden_model_1.ACC [7]);
  nor (_09204_, _09203_, _09193_);
  nor (_09205_, _09204_, _03751_);
  nor (_09206_, _09204_, _04616_);
  nor (_09207_, _04615_, _09192_);
  or (_09208_, _09207_, _09206_);
  and (_09209_, _09208_, _04630_);
  and (_09210_, _06250_, _05411_);
  nor (_09211_, _09210_, _09193_);
  nor (_09212_, _09211_, _04630_);
  or (_09213_, _09212_, _09209_);
  and (_09214_, _09213_, _04537_);
  not (_09215_, _05411_);
  nor (_09216_, _05498_, _09215_);
  nor (_09217_, _09216_, _09193_);
  nor (_09218_, _09217_, _04537_);
  nor (_09219_, _09218_, _09214_);
  nor (_09220_, _09219_, _03750_);
  or (_09221_, _09220_, _07544_);
  nor (_09222_, _09221_, _09205_);
  and (_09223_, _09217_, _07544_);
  or (_09224_, _09223_, _04678_);
  nor (_09225_, _09224_, _09222_);
  or (_09226_, _09225_, _09202_);
  and (_09227_, _09226_, _03415_);
  nor (_09228_, _06501_, _09215_);
  nor (_09229_, _09228_, _09193_);
  nor (_09230_, _09229_, _03415_);
  or (_09231_, _09230_, _08854_);
  or (_09232_, _09231_, _09227_);
  and (_09233_, _06515_, _05411_);
  or (_09234_, _09193_, _04703_);
  nor (_09235_, _09234_, _09233_);
  and (_09236_, _06307_, _05411_);
  nor (_09237_, _09236_, _09193_);
  and (_09238_, _09237_, _03839_);
  or (_09239_, _09238_, _03959_);
  nor (_09240_, _09239_, _09235_);
  and (_09241_, _09240_, _09232_);
  nor (_09242_, _09241_, _09199_);
  nor (_09243_, _09242_, _03866_);
  nor (_09244_, _09193_, _05501_);
  not (_09245_, _09244_);
  nor (_09246_, _09237_, _04708_);
  and (_09247_, _09246_, _09245_);
  nor (_09248_, _09247_, _09243_);
  nor (_09249_, _09248_, _03967_);
  nor (_09250_, _09204_, _04706_);
  and (_09251_, _09250_, _09245_);
  nor (_09252_, _09251_, _03835_);
  not (_09253_, _09252_);
  nor (_09254_, _09253_, _09249_);
  nor (_09255_, _06514_, _09215_);
  or (_09256_, _09193_, _06532_);
  nor (_09257_, _09256_, _09255_);
  or (_09258_, _09257_, _03954_);
  nor (_09259_, _09258_, _09254_);
  nor (_09260_, _06522_, _09215_);
  nor (_09261_, _09260_, _09193_);
  nor (_09262_, _09261_, _06537_);
  or (_09263_, _09262_, _09259_);
  and (_09264_, _09263_, _03704_);
  nor (_09265_, _09211_, _03704_);
  or (_09266_, _09265_, _09264_);
  and (_09267_, _09266_, _03702_);
  nor (_09268_, _09267_, _09196_);
  nand (_09269_, _09268_, _42908_);
  or (_09270_, _42908_, \oc8051_golden_model_1.TL0 [7]);
  and (_09271_, _09270_, _41654_);
  and (_40447_, _09271_, _09269_);
  not (_09272_, \oc8051_golden_model_1.TL1 [7]);
  nor (_09273_, _05516_, _09272_);
  and (_09274_, _06021_, _05428_);
  nor (_09275_, _09274_, _09273_);
  nor (_09276_, _09275_, _03702_);
  and (_09277_, _06523_, _05428_);
  nor (_09278_, _09277_, _09273_);
  nor (_09279_, _09278_, _04701_);
  and (_09280_, _06237_, _05516_);
  or (_09281_, _09280_, _09273_);
  and (_09282_, _09281_, _04678_);
  and (_09283_, _05516_, \oc8051_golden_model_1.ACC [7]);
  nor (_09284_, _09283_, _09273_);
  nor (_09285_, _09284_, _03751_);
  nor (_09286_, _09284_, _04616_);
  nor (_09287_, _04615_, _09272_);
  or (_09288_, _09287_, _09286_);
  and (_09289_, _09288_, _04630_);
  and (_09290_, _06250_, _05428_);
  nor (_09291_, _09290_, _09273_);
  nor (_09292_, _09291_, _04630_);
  or (_09293_, _09292_, _09289_);
  and (_09294_, _09293_, _04537_);
  not (_09295_, _05428_);
  nor (_09296_, _05498_, _09295_);
  nor (_09297_, _09296_, _09273_);
  nor (_09298_, _09297_, _04537_);
  nor (_09299_, _09298_, _09294_);
  nor (_09300_, _09299_, _03750_);
  or (_09301_, _09300_, _07544_);
  nor (_09302_, _09301_, _09285_);
  and (_09303_, _09297_, _07544_);
  or (_09304_, _09303_, _04678_);
  nor (_09305_, _09304_, _09302_);
  or (_09306_, _09305_, _09282_);
  and (_09307_, _09306_, _03415_);
  nor (_09308_, _06501_, _09295_);
  nor (_09309_, _09308_, _09273_);
  nor (_09310_, _09309_, _03415_);
  or (_09311_, _09310_, _08854_);
  or (_09312_, _09311_, _09307_);
  and (_09313_, _06515_, _05428_);
  or (_09314_, _09273_, _04703_);
  or (_09315_, _09314_, _09313_);
  and (_09316_, _06307_, _05516_);
  nor (_09317_, _09316_, _09273_);
  and (_09318_, _09317_, _03839_);
  nor (_09319_, _09318_, _03959_);
  and (_09320_, _09319_, _09315_);
  and (_09321_, _09320_, _09312_);
  nor (_09322_, _09321_, _09279_);
  nor (_09323_, _09322_, _03866_);
  nor (_09324_, _09273_, _05501_);
  not (_09325_, _09324_);
  nor (_09326_, _09317_, _04708_);
  and (_09327_, _09326_, _09325_);
  nor (_09328_, _09327_, _09323_);
  nor (_09329_, _09328_, _03967_);
  nor (_09330_, _09284_, _04706_);
  and (_09331_, _09330_, _09325_);
  nor (_09332_, _09331_, _03835_);
  not (_09333_, _09332_);
  nor (_09334_, _09333_, _09329_);
  or (_09335_, _06514_, _09295_);
  nor (_09336_, _09273_, _06532_);
  and (_09337_, _09336_, _09335_);
  or (_09338_, _09337_, _03954_);
  nor (_09339_, _09338_, _09334_);
  nor (_09340_, _06522_, _09295_);
  nor (_09341_, _09340_, _09273_);
  nor (_09342_, _09341_, _06537_);
  or (_09343_, _09342_, _09339_);
  and (_09344_, _09343_, _03704_);
  nor (_09345_, _09291_, _03704_);
  or (_09346_, _09345_, _09344_);
  and (_09347_, _09346_, _03702_);
  nor (_09348_, _09347_, _09276_);
  nand (_09349_, _09348_, _42908_);
  or (_09350_, _42908_, \oc8051_golden_model_1.TL1 [7]);
  and (_09351_, _09350_, _41654_);
  and (_40449_, _09351_, _09349_);
  not (_09352_, \oc8051_golden_model_1.TH0 [7]);
  nor (_09353_, _05426_, _09352_);
  and (_09354_, _06021_, _05426_);
  nor (_09355_, _09354_, _09353_);
  nor (_09356_, _09355_, _03702_);
  and (_09357_, _06523_, _05426_);
  nor (_09358_, _09357_, _09353_);
  nor (_09359_, _09358_, _04701_);
  and (_09360_, _06237_, _05426_);
  or (_09361_, _09360_, _09353_);
  and (_09362_, _09361_, _04678_);
  and (_09363_, _05426_, \oc8051_golden_model_1.ACC [7]);
  nor (_09364_, _09363_, _09353_);
  nor (_09365_, _09364_, _03751_);
  nor (_09366_, _09364_, _04616_);
  nor (_09367_, _04615_, _09352_);
  or (_09368_, _09367_, _09366_);
  and (_09369_, _09368_, _04630_);
  and (_09370_, _06250_, _05426_);
  nor (_09371_, _09370_, _09353_);
  nor (_09372_, _09371_, _04630_);
  or (_09373_, _09372_, _09369_);
  and (_09374_, _09373_, _04537_);
  not (_09375_, _05426_);
  nor (_09376_, _05498_, _09375_);
  nor (_09377_, _09376_, _09353_);
  nor (_09378_, _09377_, _04537_);
  nor (_09379_, _09378_, _09374_);
  nor (_09380_, _09379_, _03750_);
  or (_09381_, _09380_, _07544_);
  nor (_09382_, _09381_, _09365_);
  and (_09383_, _09377_, _07544_);
  or (_09384_, _09383_, _04678_);
  nor (_09385_, _09384_, _09382_);
  or (_09386_, _09385_, _09362_);
  and (_09387_, _09386_, _03415_);
  nor (_09388_, _06501_, _09375_);
  nor (_09389_, _09388_, _09353_);
  nor (_09390_, _09389_, _03415_);
  or (_09391_, _09390_, _08854_);
  or (_09392_, _09391_, _09387_);
  and (_09393_, _06515_, _05426_);
  or (_09394_, _09353_, _04703_);
  or (_09395_, _09394_, _09393_);
  and (_09396_, _06307_, _05426_);
  nor (_09397_, _09396_, _09353_);
  and (_09398_, _09397_, _03839_);
  nor (_09399_, _09398_, _03959_);
  and (_09400_, _09399_, _09395_);
  and (_09401_, _09400_, _09392_);
  nor (_09402_, _09401_, _09359_);
  nor (_09403_, _09402_, _03866_);
  nor (_09404_, _09353_, _05501_);
  not (_09405_, _09404_);
  nor (_09406_, _09397_, _04708_);
  and (_09407_, _09406_, _09405_);
  nor (_09408_, _09407_, _09403_);
  nor (_09409_, _09408_, _03967_);
  nor (_09410_, _09364_, _04706_);
  and (_09411_, _09410_, _09405_);
  nor (_09412_, _09411_, _03835_);
  not (_09413_, _09412_);
  nor (_09414_, _09413_, _09409_);
  nor (_09415_, _06514_, _09375_);
  or (_09416_, _09353_, _06532_);
  nor (_09417_, _09416_, _09415_);
  or (_09418_, _09417_, _03954_);
  nor (_09419_, _09418_, _09414_);
  nor (_09420_, _06522_, _09375_);
  nor (_09421_, _09420_, _09353_);
  nor (_09422_, _09421_, _06537_);
  or (_09423_, _09422_, _09419_);
  and (_09424_, _09423_, _03704_);
  nor (_09425_, _09371_, _03704_);
  or (_09426_, _09425_, _09424_);
  and (_09427_, _09426_, _03702_);
  nor (_09428_, _09427_, _09356_);
  nand (_09429_, _09428_, _42908_);
  or (_09430_, _42908_, \oc8051_golden_model_1.TH0 [7]);
  and (_09431_, _09430_, _41654_);
  and (_40450_, _09431_, _09429_);
  not (_09432_, \oc8051_golden_model_1.TH1 [7]);
  nor (_09433_, _05404_, _09432_);
  and (_09434_, _06021_, _05404_);
  nor (_09435_, _09434_, _09433_);
  nor (_09436_, _09435_, _03702_);
  and (_09437_, _06523_, _05404_);
  nor (_09438_, _09437_, _09433_);
  nor (_09439_, _09438_, _04701_);
  and (_09440_, _06237_, _05404_);
  or (_09441_, _09440_, _09433_);
  and (_09442_, _09441_, _04678_);
  and (_09443_, _05404_, \oc8051_golden_model_1.ACC [7]);
  nor (_09444_, _09443_, _09433_);
  nor (_09445_, _09444_, _04616_);
  nor (_09446_, _04615_, _09432_);
  or (_09447_, _09446_, _09445_);
  and (_09448_, _09447_, _04630_);
  and (_09449_, _06250_, _05404_);
  nor (_09450_, _09449_, _09433_);
  nor (_09451_, _09450_, _04630_);
  or (_09452_, _09451_, _09448_);
  and (_09453_, _09452_, _04537_);
  not (_09454_, _05404_);
  nor (_09455_, _05498_, _09454_);
  nor (_09456_, _09455_, _09433_);
  nor (_09457_, _09456_, _04537_);
  nor (_09458_, _09457_, _09453_);
  nor (_09459_, _09458_, _03750_);
  nor (_09460_, _09444_, _03751_);
  nor (_09461_, _09460_, _07544_);
  not (_09462_, _09461_);
  nor (_09463_, _09462_, _09459_);
  and (_09464_, _09456_, _07544_);
  or (_09465_, _09464_, _04678_);
  nor (_09466_, _09465_, _09463_);
  or (_09467_, _09466_, _09442_);
  and (_09468_, _09467_, _03415_);
  nor (_09469_, _06501_, _09454_);
  nor (_09470_, _09469_, _09433_);
  nor (_09471_, _09470_, _03415_);
  or (_09472_, _09471_, _08854_);
  or (_09473_, _09472_, _09468_);
  and (_09474_, _06515_, _05404_);
  or (_09475_, _09433_, _04703_);
  or (_09476_, _09475_, _09474_);
  and (_09477_, _06307_, _05404_);
  nor (_09478_, _09477_, _09433_);
  and (_09479_, _09478_, _03839_);
  nor (_09480_, _09479_, _03959_);
  and (_09481_, _09480_, _09476_);
  and (_09482_, _09481_, _09473_);
  nor (_09483_, _09482_, _09439_);
  nor (_09484_, _09483_, _03866_);
  nor (_09485_, _09433_, _05501_);
  not (_09486_, _09485_);
  nor (_09487_, _09478_, _04708_);
  and (_09488_, _09487_, _09486_);
  nor (_09489_, _09488_, _09484_);
  nor (_09490_, _09489_, _03967_);
  nor (_09491_, _09444_, _04706_);
  and (_09492_, _09491_, _09486_);
  or (_09493_, _09492_, _09490_);
  and (_09494_, _09493_, _06532_);
  nor (_09495_, _06514_, _09454_);
  nor (_09496_, _09495_, _09433_);
  nor (_09498_, _09496_, _06532_);
  or (_09499_, _09498_, _09494_);
  and (_09500_, _09499_, _06537_);
  nor (_09501_, _06522_, _09454_);
  nor (_09502_, _09501_, _09433_);
  nor (_09503_, _09502_, _06537_);
  or (_09504_, _09503_, _09500_);
  and (_09505_, _09504_, _03704_);
  nor (_09506_, _09450_, _03704_);
  or (_09507_, _09506_, _09505_);
  and (_09508_, _09507_, _03702_);
  nor (_09509_, _09508_, _09436_);
  nand (_09510_, _09509_, _42908_);
  or (_09511_, _42908_, \oc8051_golden_model_1.TH1 [7]);
  and (_09512_, _09511_, _41654_);
  and (_40451_, _09512_, _09510_);
  not (_09513_, \oc8051_golden_model_1.TMOD [7]);
  nor (_09514_, _05414_, _09513_);
  and (_09515_, _06021_, _05414_);
  nor (_09516_, _09515_, _09514_);
  nor (_09518_, _09516_, _03702_);
  and (_09519_, _06523_, _05414_);
  nor (_09520_, _09519_, _09514_);
  nor (_09521_, _09520_, _04701_);
  and (_09522_, _06237_, _05414_);
  or (_09523_, _09522_, _09514_);
  and (_09524_, _09523_, _04678_);
  and (_09525_, _05414_, \oc8051_golden_model_1.ACC [7]);
  nor (_09526_, _09525_, _09514_);
  nor (_09527_, _09526_, _04616_);
  nor (_09528_, _04615_, _09513_);
  or (_09529_, _09528_, _09527_);
  and (_09530_, _09529_, _04630_);
  and (_09531_, _06250_, _05414_);
  nor (_09532_, _09531_, _09514_);
  nor (_09533_, _09532_, _04630_);
  or (_09534_, _09533_, _09530_);
  and (_09535_, _09534_, _04537_);
  not (_09536_, _05414_);
  nor (_09537_, _05498_, _09536_);
  nor (_09538_, _09537_, _09514_);
  nor (_09539_, _09538_, _04537_);
  nor (_09540_, _09539_, _09535_);
  nor (_09541_, _09540_, _03750_);
  nor (_09542_, _09526_, _03751_);
  nor (_09543_, _09542_, _07544_);
  not (_09544_, _09543_);
  nor (_09545_, _09544_, _09541_);
  and (_09546_, _09538_, _07544_);
  or (_09547_, _09546_, _04678_);
  nor (_09548_, _09547_, _09545_);
  or (_09549_, _09548_, _09524_);
  and (_09550_, _09549_, _03415_);
  nor (_09551_, _06501_, _09536_);
  nor (_09552_, _09551_, _09514_);
  nor (_09553_, _09552_, _03415_);
  or (_09554_, _09553_, _08854_);
  or (_09555_, _09554_, _09550_);
  and (_09556_, _06515_, _05414_);
  or (_09557_, _09514_, _04703_);
  nor (_09558_, _09557_, _09556_);
  and (_09559_, _06307_, _05414_);
  nor (_09560_, _09559_, _09514_);
  and (_09561_, _09560_, _03839_);
  or (_09562_, _09561_, _03959_);
  nor (_09563_, _09562_, _09558_);
  and (_09564_, _09563_, _09555_);
  nor (_09565_, _09564_, _09521_);
  nor (_09566_, _09565_, _03866_);
  nor (_09567_, _09514_, _05501_);
  not (_09568_, _09567_);
  nor (_09569_, _09560_, _04708_);
  and (_09570_, _09569_, _09568_);
  nor (_09571_, _09570_, _09566_);
  nor (_09572_, _09571_, _03967_);
  nor (_09573_, _09526_, _04706_);
  and (_09574_, _09573_, _09568_);
  or (_09575_, _09574_, _09572_);
  and (_09576_, _09575_, _06532_);
  nor (_09577_, _06514_, _09536_);
  nor (_09578_, _09577_, _09514_);
  nor (_09579_, _09578_, _06532_);
  or (_09580_, _09579_, _09576_);
  and (_09581_, _09580_, _06537_);
  nor (_09582_, _06522_, _09536_);
  nor (_09583_, _09582_, _09514_);
  nor (_09584_, _09583_, _06537_);
  or (_09585_, _09584_, _09581_);
  and (_09586_, _09585_, _03704_);
  nor (_09587_, _09532_, _03704_);
  or (_09588_, _09587_, _09586_);
  and (_09589_, _09588_, _03702_);
  nor (_09590_, _09589_, _09518_);
  nand (_09591_, _09590_, _42908_);
  or (_09592_, _42908_, \oc8051_golden_model_1.TMOD [7]);
  and (_09593_, _09592_, _41654_);
  and (_40452_, _09593_, _09591_);
  not (_09594_, _05398_);
  and (_09595_, _09594_, \oc8051_golden_model_1.IE [7]);
  and (_09596_, _06250_, _05398_);
  or (_09597_, _09596_, _09595_);
  or (_09598_, _09597_, _04630_);
  and (_09599_, _05398_, \oc8051_golden_model_1.ACC [7]);
  or (_09600_, _09599_, _09595_);
  and (_09601_, _09600_, _04615_);
  and (_09602_, _04616_, \oc8051_golden_model_1.IE [7]);
  or (_09603_, _09602_, _03757_);
  or (_09604_, _09603_, _09601_);
  and (_09605_, _09604_, _03697_);
  and (_09606_, _09605_, _09598_);
  not (_09607_, _06101_);
  and (_09608_, _09607_, \oc8051_golden_model_1.IE [7]);
  and (_09609_, _06127_, _06101_);
  or (_09610_, _09609_, _09608_);
  and (_09611_, _09610_, _03696_);
  or (_09612_, _09611_, _03755_);
  or (_09613_, _09612_, _09606_);
  nor (_09614_, _05498_, _09594_);
  or (_09615_, _09614_, _09595_);
  or (_09616_, _09615_, _04537_);
  and (_09617_, _09616_, _09613_);
  or (_09618_, _09617_, _03750_);
  or (_09619_, _09600_, _03751_);
  and (_09620_, _09619_, _03692_);
  and (_09621_, _09620_, _09618_);
  and (_09622_, _06119_, _06101_);
  or (_09623_, _09622_, _09608_);
  and (_09624_, _09623_, _03691_);
  or (_09625_, _09624_, _03684_);
  or (_09626_, _09625_, _09621_);
  or (_09627_, _09608_, _06268_);
  and (_09628_, _09627_, _09610_);
  or (_09629_, _09628_, _03685_);
  and (_09630_, _09629_, _03680_);
  and (_09631_, _09630_, _09626_);
  nor (_09632_, _06121_, _09607_);
  or (_09633_, _09632_, _09608_);
  and (_09634_, _09633_, _03679_);
  or (_09635_, _09634_, _07544_);
  or (_09636_, _09635_, _09631_);
  or (_09637_, _09615_, _06994_);
  and (_09638_, _09637_, _09636_);
  or (_09639_, _09638_, _04678_);
  and (_09640_, _06237_, _05398_);
  or (_09641_, _09595_, _04679_);
  or (_09642_, _09641_, _09640_);
  and (_09643_, _09642_, _03415_);
  and (_09644_, _09643_, _09639_);
  nor (_09645_, _06501_, _09594_);
  or (_09646_, _09645_, _09595_);
  and (_09647_, _09646_, _07559_);
  or (_09648_, _09647_, _08854_);
  or (_09649_, _09648_, _09644_);
  and (_09650_, _06515_, _05398_);
  or (_09651_, _09595_, _04703_);
  or (_09652_, _09651_, _09650_);
  and (_09653_, _06307_, _05398_);
  or (_09654_, _09653_, _09595_);
  or (_09655_, _09654_, _04694_);
  and (_09656_, _09655_, _04701_);
  and (_09657_, _09656_, _09652_);
  and (_09658_, _09657_, _09649_);
  and (_09659_, _06523_, _05398_);
  or (_09660_, _09659_, _09595_);
  and (_09661_, _09660_, _03959_);
  or (_09662_, _09661_, _09658_);
  and (_09663_, _09662_, _04708_);
  or (_09664_, _09595_, _05501_);
  and (_09665_, _09654_, _03866_);
  and (_09666_, _09665_, _09664_);
  or (_09667_, _09666_, _09663_);
  and (_09668_, _09667_, _04706_);
  and (_09669_, _09600_, _03967_);
  and (_09670_, _09669_, _09664_);
  or (_09671_, _09670_, _03835_);
  or (_09672_, _09671_, _09668_);
  nor (_09673_, _06514_, _09594_);
  or (_09674_, _09595_, _06532_);
  or (_09675_, _09674_, _09673_);
  and (_09676_, _09675_, _06537_);
  and (_09677_, _09676_, _09672_);
  nor (_09678_, _06522_, _09594_);
  or (_09679_, _09678_, _09595_);
  and (_09680_, _09679_, _03954_);
  or (_09681_, _09680_, _03703_);
  or (_09682_, _09681_, _09677_);
  or (_09683_, _09597_, _03704_);
  and (_09684_, _09683_, _03385_);
  and (_09685_, _09684_, _09682_);
  and (_09686_, _09623_, _03384_);
  or (_09687_, _09686_, _03701_);
  or (_09688_, _09687_, _09685_);
  and (_09689_, _06021_, _05398_);
  or (_09690_, _09689_, _09595_);
  or (_09691_, _09690_, _03702_);
  and (_09692_, _09691_, _09688_);
  or (_09693_, _09692_, _42912_);
  or (_09694_, _42908_, \oc8051_golden_model_1.IE [7]);
  and (_09695_, _09694_, _41654_);
  and (_40453_, _09695_, _09693_);
  not (_09696_, _05347_);
  and (_09697_, _09696_, \oc8051_golden_model_1.IP [7]);
  and (_09698_, _06250_, _05347_);
  or (_09699_, _09698_, _09697_);
  or (_09700_, _09699_, _04630_);
  and (_09701_, _05347_, \oc8051_golden_model_1.ACC [7]);
  or (_09702_, _09701_, _09697_);
  and (_09703_, _09702_, _04615_);
  and (_09704_, _04616_, \oc8051_golden_model_1.IP [7]);
  or (_09705_, _09704_, _03757_);
  or (_09706_, _09705_, _09703_);
  and (_09707_, _09706_, _03697_);
  and (_09708_, _09707_, _09700_);
  not (_09709_, _06089_);
  and (_09710_, _09709_, \oc8051_golden_model_1.IP [7]);
  and (_09711_, _06127_, _06089_);
  or (_09712_, _09711_, _09710_);
  and (_09713_, _09712_, _03696_);
  or (_09714_, _09713_, _03755_);
  or (_09715_, _09714_, _09708_);
  nor (_09716_, _05498_, _09696_);
  or (_09717_, _09716_, _09697_);
  or (_09718_, _09717_, _04537_);
  and (_09719_, _09718_, _09715_);
  or (_09720_, _09719_, _03750_);
  or (_09721_, _09702_, _03751_);
  and (_09722_, _09721_, _03692_);
  and (_09723_, _09722_, _09720_);
  and (_09724_, _06119_, _06089_);
  or (_09725_, _09724_, _09710_);
  and (_09726_, _09725_, _03691_);
  or (_09727_, _09726_, _03684_);
  or (_09728_, _09727_, _09723_);
  or (_09729_, _09710_, _06268_);
  and (_09730_, _09729_, _09712_);
  or (_09731_, _09730_, _03685_);
  and (_09732_, _09731_, _03680_);
  and (_09733_, _09732_, _09728_);
  nor (_09734_, _06121_, _09709_);
  or (_09735_, _09734_, _09710_);
  and (_09736_, _09735_, _03679_);
  or (_09737_, _09736_, _07544_);
  or (_09738_, _09737_, _09733_);
  or (_09739_, _09717_, _06994_);
  and (_09740_, _09739_, _09738_);
  or (_09741_, _09740_, _04678_);
  and (_09742_, _06237_, _05347_);
  or (_09743_, _09697_, _04679_);
  or (_09744_, _09743_, _09742_);
  and (_09745_, _09744_, _03415_);
  and (_09746_, _09745_, _09741_);
  nor (_09747_, _06501_, _09696_);
  or (_09748_, _09747_, _09697_);
  and (_09749_, _09748_, _07559_);
  or (_09750_, _09749_, _08854_);
  or (_09751_, _09750_, _09746_);
  and (_09752_, _06515_, _05347_);
  or (_09753_, _09697_, _04703_);
  or (_09754_, _09753_, _09752_);
  and (_09755_, _06307_, _05347_);
  or (_09756_, _09755_, _09697_);
  or (_09757_, _09756_, _04694_);
  and (_09758_, _09757_, _04701_);
  and (_09759_, _09758_, _09754_);
  and (_09760_, _09759_, _09751_);
  and (_09761_, _06523_, _05347_);
  or (_09762_, _09761_, _09697_);
  and (_09763_, _09762_, _03959_);
  or (_09764_, _09763_, _09760_);
  and (_09765_, _09764_, _04708_);
  or (_09766_, _09697_, _05501_);
  and (_09767_, _09756_, _03866_);
  and (_09768_, _09767_, _09766_);
  or (_09769_, _09768_, _09765_);
  and (_09770_, _09769_, _04706_);
  and (_09771_, _09702_, _03967_);
  and (_09772_, _09771_, _09766_);
  or (_09773_, _09772_, _03835_);
  or (_09774_, _09773_, _09770_);
  nor (_09775_, _06514_, _09696_);
  or (_09776_, _09697_, _06532_);
  or (_09777_, _09776_, _09775_);
  and (_09778_, _09777_, _06537_);
  and (_09779_, _09778_, _09774_);
  nor (_09780_, _06522_, _09696_);
  or (_09781_, _09780_, _09697_);
  and (_09782_, _09781_, _03954_);
  or (_09783_, _09782_, _03703_);
  or (_09784_, _09783_, _09779_);
  or (_09785_, _09699_, _03704_);
  and (_09786_, _09785_, _03385_);
  and (_09787_, _09786_, _09784_);
  and (_09788_, _09725_, _03384_);
  or (_09789_, _09788_, _03701_);
  or (_09790_, _09789_, _09787_);
  and (_09791_, _06021_, _05347_);
  or (_09792_, _09791_, _09697_);
  or (_09793_, _09792_, _03702_);
  and (_09794_, _09793_, _09790_);
  or (_09795_, _09794_, _42912_);
  or (_09796_, _42908_, \oc8051_golden_model_1.IP [7]);
  and (_09797_, _09796_, _41654_);
  and (_40455_, _09797_, _09795_);
  or (_09798_, _42908_, \oc8051_golden_model_1.DPL [7]);
  and (_09799_, _09798_, _41654_);
  not (_09800_, \oc8051_golden_model_1.DPL [7]);
  nor (_09801_, _05545_, _09800_);
  not (_09802_, _05440_);
  nor (_09803_, _05498_, _09802_);
  or (_09804_, _09803_, _09801_);
  or (_09805_, _09804_, _06994_);
  not (_09806_, _03861_);
  and (_09807_, _06250_, _05440_);
  or (_09808_, _09807_, _09801_);
  or (_09809_, _09808_, _04630_);
  and (_09810_, _05545_, \oc8051_golden_model_1.ACC [7]);
  or (_09811_, _09810_, _09801_);
  and (_09812_, _09811_, _04615_);
  nor (_09813_, _04615_, _09800_);
  or (_09814_, _09813_, _03757_);
  or (_09815_, _09814_, _09812_);
  and (_09816_, _09815_, _04537_);
  and (_09817_, _09816_, _09809_);
  and (_09818_, _09804_, _03755_);
  or (_09819_, _09818_, _03750_);
  or (_09820_, _09819_, _09817_);
  nor (_09821_, _03452_, _03421_);
  not (_09822_, _09821_);
  or (_09823_, _09811_, _03751_);
  and (_09824_, _09823_, _09822_);
  and (_09825_, _09824_, _09820_);
  and (_09826_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_09827_, _09826_, \oc8051_golden_model_1.DPL [2]);
  and (_09828_, _09827_, \oc8051_golden_model_1.DPL [3]);
  and (_09829_, _09828_, \oc8051_golden_model_1.DPL [4]);
  and (_09830_, _09829_, \oc8051_golden_model_1.DPL [5]);
  and (_09831_, _09830_, \oc8051_golden_model_1.DPL [6]);
  nor (_09832_, _09831_, \oc8051_golden_model_1.DPL [7]);
  and (_09833_, _09831_, \oc8051_golden_model_1.DPL [7]);
  nor (_09834_, _09833_, _09832_);
  and (_09835_, _09834_, _09821_);
  or (_09836_, _09835_, _09825_);
  and (_09837_, _09836_, _09806_);
  nor (_09838_, _06070_, _09806_);
  or (_09839_, _09838_, _07544_);
  or (_09840_, _09839_, _09837_);
  and (_09841_, _09840_, _09805_);
  or (_09842_, _09841_, _04678_);
  or (_09843_, _09801_, _04679_);
  and (_09844_, _06237_, _05545_);
  or (_09845_, _09844_, _09843_);
  and (_09846_, _09845_, _03415_);
  and (_09847_, _09846_, _09842_);
  not (_09848_, _05545_);
  nor (_09849_, _06501_, _09848_);
  or (_09850_, _09849_, _09801_);
  and (_09851_, _09850_, _07559_);
  or (_09852_, _09851_, _09847_);
  or (_09853_, _09852_, _08854_);
  and (_09854_, _06515_, _05440_);
  or (_09855_, _09801_, _04703_);
  or (_09856_, _09855_, _09854_);
  and (_09857_, _06307_, _05545_);
  or (_09858_, _09857_, _09801_);
  or (_09859_, _09858_, _04694_);
  and (_09860_, _09859_, _04701_);
  and (_09861_, _09860_, _09856_);
  and (_09862_, _09861_, _09853_);
  and (_09863_, _06523_, _05440_);
  or (_09864_, _09863_, _09801_);
  and (_09865_, _09864_, _03959_);
  or (_09866_, _09865_, _09862_);
  and (_09867_, _09866_, _04708_);
  or (_09868_, _09801_, _05501_);
  and (_09869_, _09858_, _03866_);
  and (_09870_, _09869_, _09868_);
  or (_09871_, _09870_, _09867_);
  and (_09872_, _09871_, _04706_);
  and (_09873_, _09811_, _03967_);
  and (_09874_, _09873_, _09868_);
  or (_09875_, _09874_, _03835_);
  or (_09876_, _09875_, _09872_);
  nor (_09877_, _06514_, _09802_);
  or (_09878_, _09801_, _06532_);
  or (_09879_, _09878_, _09877_);
  and (_09880_, _09879_, _06537_);
  and (_09881_, _09880_, _09876_);
  nor (_09882_, _06522_, _09802_);
  or (_09883_, _09882_, _09801_);
  and (_09884_, _09883_, _03954_);
  or (_09885_, _09884_, _03703_);
  or (_09886_, _09885_, _09881_);
  or (_09887_, _09808_, _03704_);
  and (_09888_, _09887_, _03702_);
  and (_09889_, _09888_, _09886_);
  and (_09890_, _06021_, _05440_);
  or (_09891_, _09890_, _09801_);
  and (_09892_, _09891_, _03701_);
  or (_09893_, _09892_, _42912_);
  or (_09894_, _09893_, _09889_);
  and (_40456_, _09894_, _09799_);
  or (_09895_, _42908_, \oc8051_golden_model_1.DPH [7]);
  and (_09896_, _09895_, _41654_);
  not (_09897_, \oc8051_golden_model_1.DPH [7]);
  nor (_09898_, _05422_, _09897_);
  not (_09899_, _05422_);
  nor (_09900_, _05498_, _09899_);
  or (_09901_, _09900_, _09898_);
  or (_09902_, _09901_, _06994_);
  and (_09903_, _06250_, _05422_);
  or (_09904_, _09903_, _09898_);
  or (_09905_, _09904_, _04630_);
  and (_09906_, _05422_, \oc8051_golden_model_1.ACC [7]);
  or (_09907_, _09906_, _09898_);
  and (_09908_, _09907_, _04615_);
  nor (_09909_, _04615_, _09897_);
  or (_09910_, _09909_, _03757_);
  or (_09911_, _09910_, _09908_);
  and (_09912_, _09911_, _04537_);
  and (_09913_, _09912_, _09905_);
  and (_09914_, _09901_, _03755_);
  or (_09915_, _09914_, _03750_);
  or (_09916_, _09915_, _09913_);
  or (_09917_, _09907_, _03751_);
  and (_09918_, _09917_, _09822_);
  and (_09919_, _09918_, _09916_);
  and (_09920_, _09833_, \oc8051_golden_model_1.DPH [0]);
  and (_09921_, _09920_, \oc8051_golden_model_1.DPH [1]);
  and (_09922_, _09921_, \oc8051_golden_model_1.DPH [2]);
  and (_09923_, _09922_, \oc8051_golden_model_1.DPH [3]);
  and (_09924_, _09923_, \oc8051_golden_model_1.DPH [4]);
  and (_09925_, _09924_, \oc8051_golden_model_1.DPH [5]);
  nand (_09926_, _09925_, \oc8051_golden_model_1.DPH [6]);
  or (_09927_, _09926_, _09897_);
  nand (_09928_, _09926_, _09897_);
  and (_09929_, _09928_, _09821_);
  and (_09930_, _09929_, _09927_);
  or (_09931_, _09930_, _09919_);
  and (_09932_, _09931_, _09806_);
  and (_09933_, _03861_, _03638_);
  or (_09934_, _09933_, _07544_);
  or (_09935_, _09934_, _09932_);
  and (_09936_, _09935_, _09902_);
  or (_09937_, _09936_, _04678_);
  and (_09938_, _06237_, _05422_);
  or (_09939_, _09898_, _04679_);
  or (_09940_, _09939_, _09938_);
  and (_09941_, _09940_, _03415_);
  and (_09942_, _09941_, _09937_);
  nor (_09943_, _06501_, _09899_);
  or (_09944_, _09943_, _09898_);
  and (_09945_, _09944_, _07559_);
  or (_09946_, _09945_, _09942_);
  or (_09947_, _09946_, _08854_);
  and (_09948_, _06515_, _05422_);
  or (_09949_, _09898_, _04703_);
  or (_09950_, _09949_, _09948_);
  and (_09951_, _06307_, _05422_);
  or (_09952_, _09951_, _09898_);
  or (_09953_, _09952_, _04694_);
  and (_09954_, _09953_, _04701_);
  and (_09955_, _09954_, _09950_);
  and (_09956_, _09955_, _09947_);
  and (_09957_, _06523_, _05422_);
  or (_09958_, _09957_, _09898_);
  and (_09959_, _09958_, _03959_);
  or (_09960_, _09959_, _09956_);
  and (_09961_, _09960_, _04708_);
  or (_09962_, _09898_, _05501_);
  and (_09963_, _09952_, _03866_);
  and (_09964_, _09963_, _09962_);
  or (_09965_, _09964_, _09961_);
  and (_09966_, _09965_, _04706_);
  and (_09967_, _09907_, _03967_);
  and (_09968_, _09967_, _09962_);
  or (_09969_, _09968_, _03835_);
  or (_09970_, _09969_, _09966_);
  nor (_09971_, _06514_, _09899_);
  or (_09972_, _09898_, _06532_);
  or (_09973_, _09972_, _09971_);
  and (_09974_, _09973_, _06537_);
  and (_09975_, _09974_, _09970_);
  nor (_09976_, _06522_, _09899_);
  or (_09977_, _09976_, _09898_);
  and (_09978_, _09977_, _03954_);
  or (_09979_, _09978_, _03703_);
  or (_09980_, _09979_, _09975_);
  or (_09981_, _09904_, _03704_);
  and (_09982_, _09981_, _03702_);
  and (_09983_, _09982_, _09980_);
  and (_09984_, _06021_, _05422_);
  or (_09985_, _09984_, _09898_);
  and (_09986_, _09985_, _03701_);
  or (_09987_, _09986_, _42912_);
  or (_09988_, _09987_, _09983_);
  and (_40457_, _09988_, _09896_);
  nor (_09989_, _08691_, _03709_);
  not (_09990_, _09989_);
  not (_09991_, _03115_);
  and (_09992_, _06024_, _09991_);
  and (_09993_, _09992_, \oc8051_golden_model_1.PC [7]);
  and (_09994_, _09993_, \oc8051_golden_model_1.PC [8]);
  and (_09995_, _09994_, \oc8051_golden_model_1.PC [9]);
  and (_09996_, _09995_, \oc8051_golden_model_1.PC [10]);
  and (_09997_, _09996_, \oc8051_golden_model_1.PC [11]);
  and (_09998_, _09997_, \oc8051_golden_model_1.PC [12]);
  and (_09999_, _09998_, \oc8051_golden_model_1.PC [13]);
  and (_10000_, _09999_, \oc8051_golden_model_1.PC [14]);
  or (_10001_, _10000_, \oc8051_golden_model_1.PC [15]);
  nand (_10002_, _10000_, \oc8051_golden_model_1.PC [15]);
  and (_10003_, _10002_, _10001_);
  not (_10004_, _07966_);
  and (_10005_, _03858_, _03393_);
  not (_10006_, _10005_);
  and (_10007_, _10006_, _08643_);
  and (_10008_, _10007_, _10004_);
  or (_10009_, _10008_, _10003_);
  nor (_10010_, _08580_, _03963_);
  not (_10011_, _10010_);
  and (_10012_, _08547_, _08080_);
  or (_10013_, _10012_, _10003_);
  and (_10014_, _03480_, _03383_);
  not (_10015_, _10014_);
  nor (_10016_, _03954_, _03481_);
  or (_10017_, _10016_, _06977_);
  and (_10018_, _10017_, _10015_);
  and (_10019_, _04671_, _03480_);
  not (_10020_, _10019_);
  not (_10021_, _08521_);
  and (_10022_, _03785_, _03480_);
  and (_10023_, _10022_, _03420_);
  nor (_10024_, _08640_, _04353_);
  nor (_10025_, _10024_, _10023_);
  and (_10026_, _10025_, _10021_);
  and (_10027_, _10026_, _10020_);
  or (_10028_, _10027_, _10003_);
  and (_10029_, _03476_, _03383_);
  not (_10030_, _10029_);
  nor (_10031_, _03967_, _03477_);
  or (_10032_, _10031_, _06977_);
  and (_10033_, _10032_, _10030_);
  and (_10034_, _06972_, \oc8051_golden_model_1.PC [12]);
  and (_10035_, _10034_, \oc8051_golden_model_1.PC [13]);
  and (_10036_, _10035_, \oc8051_golden_model_1.PC [14]);
  nor (_10037_, _10035_, \oc8051_golden_model_1.PC [14]);
  nor (_10038_, _10037_, _10036_);
  and (_10039_, _10038_, _03638_);
  nor (_10040_, _10038_, _03638_);
  nor (_10041_, _10040_, _10039_);
  not (_10042_, _10041_);
  nor (_10043_, _10034_, \oc8051_golden_model_1.PC [13]);
  nor (_10044_, _10043_, _10035_);
  and (_10045_, _10044_, _03638_);
  nor (_10046_, _10044_, _03638_);
  nor (_10047_, _06972_, \oc8051_golden_model_1.PC [12]);
  nor (_10048_, _10047_, _10034_);
  and (_10049_, _10048_, _03638_);
  nor (_10050_, _06970_, \oc8051_golden_model_1.PC [10]);
  nor (_10051_, _10050_, _06971_);
  and (_10052_, _10051_, _03638_);
  not (_10053_, _10052_);
  nor (_10054_, _06971_, \oc8051_golden_model_1.PC [11]);
  nor (_10055_, _10054_, _06972_);
  and (_10056_, _10055_, _03638_);
  nor (_10057_, _10055_, _03638_);
  nor (_10058_, _10057_, _10056_);
  nor (_10059_, _10051_, _03638_);
  nor (_10060_, _10059_, _10052_);
  and (_10061_, _10060_, _10058_);
  nor (_10062_, _06969_, \oc8051_golden_model_1.PC [9]);
  nor (_10063_, _10062_, _06970_);
  and (_10064_, _10063_, _03638_);
  nor (_10065_, _10063_, _03638_);
  nor (_10066_, _10065_, _10064_);
  and (_10067_, _06028_, _03638_);
  nor (_10068_, _06028_, _03638_);
  and (_10069_, _06023_, _03514_);
  nor (_10070_, _10069_, \oc8051_golden_model_1.PC [6]);
  nor (_10071_, _10070_, _06025_);
  not (_10072_, _10071_);
  nor (_10073_, _10072_, _03740_);
  and (_10074_, _10072_, _03740_);
  nor (_10075_, _10074_, _10073_);
  not (_10076_, _10075_);
  and (_10077_, _03514_, \oc8051_golden_model_1.PC [4]);
  nor (_10078_, _10077_, \oc8051_golden_model_1.PC [5]);
  nor (_10079_, _10078_, _10069_);
  not (_10080_, _10079_);
  nor (_10081_, _10080_, _04034_);
  and (_10082_, _10080_, _04034_);
  nor (_10083_, _03514_, \oc8051_golden_model_1.PC [4]);
  nor (_10084_, _10083_, _10077_);
  not (_10085_, _10084_);
  nor (_10086_, _10085_, _04446_);
  nor (_10087_, _03669_, _03879_);
  and (_10088_, _03669_, _03879_);
  not (_10089_, _03405_);
  nor (_10090_, _04165_, _10089_);
  nor (_10091_, _04482_, \oc8051_golden_model_1.PC [1]);
  nor (_10092_, _04211_, _03129_);
  and (_10093_, _04482_, \oc8051_golden_model_1.PC [1]);
  nor (_10094_, _10093_, _10091_);
  and (_10095_, _10094_, _10092_);
  nor (_10096_, _10095_, _10091_);
  and (_10097_, _04165_, _10089_);
  nor (_10098_, _10097_, _10090_);
  not (_10099_, _10098_);
  nor (_10100_, _10099_, _10096_);
  nor (_10101_, _10100_, _10090_);
  nor (_10102_, _10101_, _10088_);
  nor (_10103_, _10102_, _10087_);
  and (_10104_, _10085_, _04446_);
  nor (_10105_, _10104_, _10086_);
  not (_10106_, _10105_);
  nor (_10107_, _10106_, _10103_);
  nor (_10108_, _10107_, _10086_);
  nor (_10109_, _10108_, _10082_);
  nor (_10110_, _10109_, _10081_);
  nor (_10111_, _10110_, _10076_);
  nor (_10112_, _10111_, _10073_);
  nor (_10113_, _10112_, _10068_);
  or (_10114_, _10113_, _10067_);
  nor (_10115_, _06026_, \oc8051_golden_model_1.PC [8]);
  nor (_10116_, _10115_, _06969_);
  and (_10117_, _10116_, _03638_);
  nor (_10118_, _10116_, _03638_);
  nor (_10119_, _10118_, _10117_);
  and (_10120_, _10119_, _10114_);
  and (_10121_, _10120_, _10066_);
  and (_10122_, _10121_, _10061_);
  nor (_10123_, _10117_, _10064_);
  not (_10124_, _10123_);
  and (_10125_, _10124_, _10061_);
  or (_10126_, _10125_, _10056_);
  nor (_10127_, _10126_, _10122_);
  and (_10128_, _10127_, _10053_);
  nor (_10129_, _10048_, _03638_);
  nor (_10130_, _10129_, _10049_);
  not (_10131_, _10130_);
  nor (_10132_, _10131_, _10128_);
  nor (_10133_, _10132_, _10049_);
  nor (_10134_, _10133_, _10046_);
  nor (_10135_, _10134_, _10045_);
  nor (_10136_, _10135_, _10042_);
  nor (_10137_, _10136_, _10039_);
  nor (_10138_, _06977_, _03638_);
  and (_10139_, _06977_, _03638_);
  nor (_10140_, _10139_, _10138_);
  and (_10141_, _10140_, _10137_);
  nor (_10142_, _10140_, _10137_);
  or (_10143_, _10142_, _10141_);
  or (_10144_, _10143_, _08783_);
  and (_10145_, _03482_, _03383_);
  not (_10146_, _08783_);
  or (_10147_, _10146_, _06977_);
  and (_10148_, _10147_, _10145_);
  and (_10149_, _10148_, _10144_);
  or (_10150_, _06977_, _06305_);
  and (_10151_, _06967_, _07559_);
  or (_10152_, _06237_, _05351_);
  and (_10153_, _10152_, _06281_);
  or (_10154_, _06933_, _03740_);
  or (_10155_, _06607_, _05165_);
  and (_10156_, _10155_, _10154_);
  and (_10157_, _10156_, _10153_);
  or (_10158_, _06836_, _05362_);
  or (_10159_, _06941_, _04034_);
  and (_10160_, _10159_, _10158_);
  or (_10161_, _06881_, _05357_);
  or (_10162_, _06942_, _04446_);
  and (_10163_, _10162_, _10161_);
  and (_10164_, _10163_, _10160_);
  and (_10165_, _10164_, _10157_);
  or (_10166_, _06937_, _03669_);
  or (_10167_, _06744_, _03742_);
  and (_10168_, _10167_, _10166_);
  or (_10169_, _06938_, _04165_);
  or (_10170_, _06789_, _05174_);
  and (_10171_, _10170_, _10169_);
  and (_10172_, _10171_, _10168_);
  or (_10173_, _06698_, _04344_);
  or (_10174_, _06653_, _04750_);
  or (_10175_, _06934_, _04482_);
  and (_10176_, _10175_, _10174_);
  and (_10177_, _10176_, _10173_);
  or (_10178_, _06935_, _04211_);
  and (_10179_, _10178_, _10177_);
  and (_10180_, _10179_, _10172_);
  and (_10181_, _10180_, _10165_);
  and (_10182_, _10181_, _06967_);
  not (_10183_, _10181_);
  and (_10184_, _06961_, \oc8051_golden_model_1.PC [12]);
  and (_10185_, _10184_, \oc8051_golden_model_1.PC [13]);
  and (_10186_, _10185_, \oc8051_golden_model_1.PC [14]);
  nor (_10187_, _10185_, \oc8051_golden_model_1.PC [14]);
  nor (_10188_, _10187_, _10186_);
  not (_10189_, _10188_);
  nor (_10190_, _10189_, _06070_);
  and (_10191_, _10189_, _06070_);
  nor (_10192_, _10191_, _10190_);
  not (_10193_, _10192_);
  nor (_10194_, _10184_, \oc8051_golden_model_1.PC [13]);
  nor (_10195_, _10194_, _10185_);
  not (_10196_, _10195_);
  nor (_10197_, _10196_, _06070_);
  and (_10198_, _10196_, _06070_);
  nor (_10199_, _06961_, \oc8051_golden_model_1.PC [12]);
  nor (_10200_, _10199_, _10184_);
  not (_10201_, _10200_);
  nor (_10202_, _10201_, _06070_);
  nor (_10203_, _06960_, \oc8051_golden_model_1.PC [11]);
  nor (_10204_, _10203_, _06961_);
  not (_10205_, _10204_);
  nor (_10206_, _10205_, _06070_);
  and (_10207_, _10205_, _06070_);
  nor (_10208_, _10207_, _10206_);
  nor (_10209_, _06959_, \oc8051_golden_model_1.PC [10]);
  nor (_10210_, _10209_, _06960_);
  not (_10211_, _10210_);
  nor (_10212_, _10211_, _06070_);
  and (_10213_, _10211_, _06070_);
  nor (_10214_, _10213_, _10212_);
  and (_10215_, _10214_, _10208_);
  nor (_10216_, _06958_, \oc8051_golden_model_1.PC [9]);
  nor (_10217_, _10216_, _06959_);
  not (_10218_, _10217_);
  nor (_10219_, _10218_, _06070_);
  and (_10220_, _10218_, _06070_);
  nor (_10221_, _10220_, _10219_);
  nor (_10222_, _06900_, _06070_);
  and (_10223_, _06900_, _06070_);
  and (_10224_, _06895_, _06023_);
  nor (_10225_, _10224_, \oc8051_golden_model_1.PC [6]);
  nor (_10226_, _10225_, _06896_);
  not (_10227_, _10226_);
  nor (_10228_, _10227_, _06406_);
  and (_10229_, _10227_, _06406_);
  nor (_10230_, _10229_, _10228_);
  not (_10231_, _10230_);
  and (_10232_, _06895_, \oc8051_golden_model_1.PC [4]);
  nor (_10233_, _10232_, \oc8051_golden_model_1.PC [5]);
  nor (_10234_, _10233_, _10224_);
  not (_10235_, _10234_);
  nor (_10236_, _10235_, _06370_);
  and (_10237_, _10235_, _06370_);
  nor (_10238_, _06895_, \oc8051_golden_model_1.PC [4]);
  nor (_10239_, _10238_, _10232_);
  not (_10240_, _10239_);
  nor (_10241_, _10240_, _06339_);
  nor (_10242_, _06894_, \oc8051_golden_model_1.PC [3]);
  nor (_10243_, _10242_, _06895_);
  not (_10244_, _10243_);
  nor (_10245_, _10244_, _03946_);
  and (_10246_, _10244_, _03946_);
  nor (_10247_, _03134_, \oc8051_golden_model_1.PC [2]);
  nor (_10248_, _10247_, _06894_);
  not (_10249_, _10248_);
  nor (_10250_, _10249_, _04077_);
  not (_10251_, _03492_);
  nor (_10252_, _04515_, _10251_);
  nor (_10253_, _04326_, \oc8051_golden_model_1.PC [0]);
  and (_10254_, _04515_, _10251_);
  nor (_10255_, _10254_, _10252_);
  and (_10256_, _10255_, _10253_);
  nor (_10257_, _10256_, _10252_);
  and (_10258_, _10249_, _04077_);
  nor (_10259_, _10258_, _10250_);
  not (_10260_, _10259_);
  nor (_10261_, _10260_, _10257_);
  nor (_10262_, _10261_, _10250_);
  nor (_10263_, _10262_, _10246_);
  nor (_10264_, _10263_, _10245_);
  and (_10265_, _10240_, _06339_);
  nor (_10266_, _10265_, _10241_);
  not (_10267_, _10266_);
  nor (_10268_, _10267_, _10264_);
  nor (_10269_, _10268_, _10241_);
  nor (_10270_, _10269_, _10237_);
  nor (_10271_, _10270_, _10236_);
  nor (_10272_, _10271_, _10231_);
  nor (_10273_, _10272_, _10228_);
  nor (_10274_, _10273_, _10223_);
  or (_10275_, _10274_, _10222_);
  nor (_10276_, _06897_, \oc8051_golden_model_1.PC [8]);
  nor (_10277_, _10276_, _06958_);
  not (_10278_, _10277_);
  nor (_10279_, _10278_, _06070_);
  and (_10280_, _10278_, _06070_);
  nor (_10281_, _10280_, _10279_);
  and (_10282_, _10281_, _10275_);
  and (_10283_, _10282_, _10221_);
  and (_10284_, _10283_, _10215_);
  nor (_10285_, _10279_, _10219_);
  not (_10286_, _10285_);
  and (_10287_, _10286_, _10215_);
  or (_10288_, _10287_, _10212_);
  or (_10289_, _10288_, _10284_);
  nor (_10290_, _10289_, _10206_);
  and (_10291_, _10201_, _06070_);
  nor (_10292_, _10291_, _10202_);
  not (_10293_, _10292_);
  nor (_10294_, _10293_, _10290_);
  nor (_10295_, _10294_, _10202_);
  nor (_10296_, _10295_, _10198_);
  nor (_10297_, _10296_, _10197_);
  nor (_10298_, _10297_, _10193_);
  nor (_10299_, _10298_, _10190_);
  not (_10300_, _06967_);
  and (_10301_, _10300_, _06070_);
  nor (_10302_, _10300_, _06070_);
  nor (_10303_, _10302_, _10301_);
  and (_10304_, _10303_, _10299_);
  nor (_10305_, _10303_, _10299_);
  or (_10306_, _10305_, _10304_);
  and (_10307_, _10306_, _10183_);
  or (_10308_, _10307_, _03855_);
  or (_10309_, _10308_, _10182_);
  and (_10310_, _06977_, _03750_);
  and (_10311_, _05652_, _05602_);
  and (_10312_, _06243_, _10311_);
  and (_10313_, _06241_, _06016_);
  and (_10314_, _10313_, _10312_);
  and (_10315_, _10314_, _06967_);
  nand (_10316_, _10313_, _10312_);
  and (_10317_, _10316_, _10306_);
  or (_10318_, _10317_, _10315_);
  and (_10319_, _10318_, _03757_);
  not (_10320_, _06140_);
  and (_10321_, _06132_, _06130_);
  and (_10322_, _04842_, _04608_);
  and (_10323_, _06921_, _10322_);
  nand (_10324_, _10323_, _10321_);
  and (_10325_, _10324_, _10143_);
  and (_10326_, _10323_, _10321_);
  and (_10327_, _10326_, _06977_);
  or (_10328_, _10327_, _10325_);
  and (_10329_, _10328_, _10320_);
  and (_10330_, _10003_, _04234_);
  not (_10331_, _04109_);
  and (_10332_, _06977_, _04083_);
  or (_10333_, _10332_, _10331_);
  nand (_10334_, _04944_, _06957_);
  or (_10335_, _10003_, _04944_);
  and (_10336_, _10335_, _10334_);
  or (_10337_, _10336_, _04615_);
  and (_10338_, _10337_, _10333_);
  or (_10339_, _10338_, _10330_);
  and (_10340_, _10339_, _04948_);
  nand (_10341_, _06977_, _04111_);
  not (_10342_, _08105_);
  nor (_10343_, _08107_, _08117_);
  and (_10344_, _10343_, _10342_);
  nand (_10345_, _10344_, _10341_);
  or (_10346_, _10345_, _10340_);
  or (_10347_, _10344_, _10003_);
  and (_10348_, _10347_, _06140_);
  and (_10349_, _10348_, _10346_);
  or (_10350_, _10349_, _04624_);
  or (_10351_, _10350_, _10329_);
  and (_10352_, _10351_, _04630_);
  nor (_10353_, _03444_, _03421_);
  nor (_10354_, _10353_, _08120_);
  not (_10355_, _10354_);
  or (_10356_, _10355_, _10352_);
  or (_10357_, _10356_, _10319_);
  and (_10358_, _04818_, _03318_);
  nor (_10359_, _10358_, _03696_);
  and (_10360_, _10354_, _04625_);
  or (_10361_, _10360_, _10003_);
  and (_10362_, _10361_, _10359_);
  and (_10363_, _10362_, _10357_);
  nor (_10364_, _04839_, _04645_);
  not (_10365_, _10364_);
  not (_10366_, _10359_);
  and (_10367_, _10366_, _06977_);
  or (_10368_, _10367_, _10365_);
  or (_10369_, _10368_, _10363_);
  or (_10370_, _10364_, _10003_);
  and (_10371_, _10370_, _03751_);
  and (_10372_, _10371_, _10369_);
  or (_10373_, _10372_, _10310_);
  nor (_10374_, _03447_, _03421_);
  nor (_10375_, _10374_, _08098_);
  and (_10376_, _10375_, _10373_);
  not (_10377_, _10375_);
  and (_10378_, _10377_, _10003_);
  not (_10379_, _03448_);
  nor (_10380_, _03690_, _10379_);
  and (_10381_, _10380_, _03692_);
  not (_10382_, _10381_);
  or (_10383_, _10382_, _10378_);
  or (_10384_, _10383_, _10376_);
  or (_10385_, _10381_, _06977_);
  and (_10386_, _03789_, _03683_);
  nor (_10387_, _06992_, _03441_);
  nor (_10388_, _10387_, _10386_);
  and (_10389_, _10388_, _10385_);
  and (_10390_, _10389_, _10384_);
  not (_10391_, _05499_);
  and (_10392_, _05498_, _03638_);
  nor (_10393_, _10392_, _10391_);
  nor (_10394_, _06013_, _05165_);
  and (_10395_, _06013_, _05165_);
  nor (_10396_, _10395_, _10394_);
  and (_10397_, _10396_, _10393_);
  or (_10398_, _05799_, _05362_);
  and (_10399_, _05799_, _05362_);
  not (_10400_, _10399_);
  and (_10401_, _10400_, _10398_);
  and (_10402_, _05898_, _05357_);
  nor (_10403_, _05898_, _05357_);
  nor (_10404_, _10403_, _10402_);
  and (_10405_, _10404_, _10401_);
  and (_10406_, _10405_, _10397_);
  and (_10407_, _05050_, _03742_);
  and (_10408_, _05236_, _05174_);
  nor (_10409_, _10408_, _10407_);
  or (_10410_, _05050_, _03742_);
  or (_10411_, _05236_, _05174_);
  and (_10412_, _10411_, _10410_);
  and (_10413_, _10412_, _10409_);
  or (_10414_, _04842_, _04750_);
  and (_10415_, _04842_, _04750_);
  not (_10416_, _10415_);
  and (_10417_, _10416_, _10414_);
  nand (_10418_, _04608_, _04211_);
  or (_10419_, _04608_, _04211_);
  and (_10420_, _10419_, _10418_);
  and (_10421_, _10420_, _10417_);
  and (_10422_, _10421_, _10413_);
  and (_10423_, _10422_, _10406_);
  nand (_10424_, _10423_, _10300_);
  not (_10425_, _10388_);
  or (_10426_, _10423_, _10306_);
  and (_10427_, _10426_, _10425_);
  and (_10428_, _10427_, _10424_);
  or (_10429_, _10428_, _03854_);
  or (_10430_, _10429_, _10390_);
  nor (_10431_, _03441_, _03421_);
  not (_10432_, _10431_);
  and (_10433_, _10432_, _03848_);
  and (_10434_, _10433_, _10430_);
  and (_10435_, _10434_, _10309_);
  nor (_10436_, _08736_, _08740_);
  nor (_10437_, _08733_, _08485_);
  and (_10438_, _10437_, _10436_);
  nor (_10439_, _08741_, _08742_);
  nor (_10440_, _10439_, _08745_);
  and (_10441_, _04211_, _03558_);
  nor (_10442_, _10441_, _08748_);
  not (_10443_, _10442_);
  and (_10444_, _08751_, _10443_);
  and (_10445_, _10444_, _10440_);
  and (_10446_, _10445_, _10438_);
  or (_10447_, _10446_, _10306_);
  nand (_10448_, _10446_, _10300_);
  and (_10449_, _10448_, _03847_);
  and (_10450_, _10449_, _10447_);
  nor (_10451_, _08697_, _08696_);
  nor (_10452_, _10451_, _08700_);
  nor (_10453_, _08695_, _06523_);
  and (_10454_, _10453_, _10452_);
  nor (_10455_, _08703_, _08701_);
  nor (_10456_, _10455_, _08707_);
  not (_10457_, _08711_);
  nor (_10458_, _05652_, \oc8051_golden_model_1.ACC [0]);
  or (_10459_, _10458_, _08712_);
  and (_10460_, _10459_, _10457_);
  and (_10461_, _10460_, _10456_);
  and (_10462_, _10461_, _10454_);
  nand (_10463_, _10462_, _10300_);
  or (_10464_, _10462_, _10306_);
  and (_10465_, _10464_, _03773_);
  and (_10466_, _10465_, _10463_);
  or (_10467_, _10466_, _10450_);
  nand (_10468_, _10431_, _10003_);
  and (_10469_, _05106_, _03778_);
  and (_10470_, _10469_, _03807_);
  nand (_10471_, _10470_, _10468_);
  or (_10472_, _10471_, _10467_);
  or (_10473_, _10472_, _10435_);
  nor (_10474_, _03452_, _03414_);
  not (_10475_, _10474_);
  nor (_10476_, _09821_, _07024_);
  and (_10477_, _10476_, _10475_);
  or (_10478_, _10470_, _06977_);
  and (_10479_, _10478_, _10477_);
  and (_10480_, _10479_, _10473_);
  not (_10481_, _10477_);
  and (_10482_, _10481_, _10003_);
  and (_10483_, _04856_, _03318_);
  nor (_10484_, _10483_, _03811_);
  not (_10485_, _10484_);
  or (_10486_, _10485_, _10482_);
  or (_10487_, _10486_, _10480_);
  nor (_10488_, _08260_, _08182_);
  or (_10489_, _10484_, _06977_);
  and (_10490_, _10489_, _10488_);
  and (_10491_, _10490_, _10487_);
  nor (_10492_, _08287_, _03818_);
  not (_10493_, _10492_);
  not (_10494_, _10488_);
  and (_10495_, _10494_, _10003_);
  or (_10496_, _10495_, _10493_);
  or (_10497_, _10496_, _10491_);
  or (_10498_, _10492_, _06977_);
  and (_10499_, _10498_, _03422_);
  and (_10500_, _10499_, _10497_);
  and (_10501_, _10003_, _03547_);
  nor (_10502_, _03679_, _03676_);
  not (_10503_, _10502_);
  or (_10504_, _10503_, _10501_);
  or (_10505_, _10504_, _10500_);
  or (_10506_, _10502_, _06977_);
  and (_10507_, _10506_, _09806_);
  and (_10508_, _10507_, _10505_);
  nand (_10509_, _06967_, _03861_);
  and (_10510_, _06994_, _04679_);
  nand (_10511_, _10510_, _10509_);
  or (_10512_, _10511_, _10508_);
  or (_10513_, _10510_, _06977_);
  and (_10514_, _10513_, _03415_);
  and (_10515_, _10514_, _10512_);
  or (_10516_, _10515_, _10151_);
  nor (_10517_, _07558_, _03466_);
  and (_10518_, _10517_, _10516_);
  nor (_10519_, _03746_, _03487_);
  not (_10520_, _10519_);
  not (_10521_, _10517_);
  and (_10522_, _10521_, _10003_);
  or (_10523_, _10522_, _10520_);
  or (_10524_, _10523_, _10518_);
  and (_10525_, _03410_, _03383_);
  not (_10526_, _10525_);
  or (_10527_, _10519_, _06977_);
  and (_10528_, _10527_, _10526_);
  and (_10529_, _10528_, _10524_);
  and (_10530_, _10525_, _10143_);
  or (_10531_, _10530_, _06306_);
  or (_10532_, _10531_, _10529_);
  and (_10533_, _10532_, _10150_);
  or (_10534_, _10533_, _03839_);
  or (_10535_, _06967_, _04694_);
  and (_10536_, _10535_, _08457_);
  and (_10537_, _10536_, _10534_);
  and (_10538_, _08456_, _06977_);
  or (_10539_, _10538_, _10537_);
  and (_10540_, _03482_, _03834_);
  not (_10541_, _10540_);
  and (_10542_, _10541_, _10539_);
  nor (_10543_, _03745_, _03483_);
  not (_10544_, _10543_);
  not (_10545_, \oc8051_golden_model_1.DPH [0]);
  and (_10546_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_10547_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_10548_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_10549_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_10550_, _10549_, _10548_);
  not (_10551_, _10550_);
  and (_10552_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_10553_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  and (_10554_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_10555_, _03524_, _03520_);
  nor (_10556_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_10557_, _10556_, _10554_);
  not (_10558_, _10557_);
  nor (_10559_, _10558_, _10555_);
  nor (_10560_, _10559_, _10554_);
  nor (_10561_, _10560_, _10553_);
  nor (_10562_, _10561_, _10552_);
  nor (_10563_, _10562_, _10551_);
  nor (_10564_, _10563_, _10548_);
  nor (_10565_, _10564_, _10547_);
  nor (_10566_, _10565_, _10546_);
  nor (_10567_, _10566_, _10545_);
  and (_10568_, _10567_, \oc8051_golden_model_1.DPH [1]);
  and (_10569_, _10568_, \oc8051_golden_model_1.DPH [2]);
  and (_10570_, _10569_, \oc8051_golden_model_1.DPH [3]);
  and (_10571_, _10570_, \oc8051_golden_model_1.DPH [4]);
  and (_10572_, _10571_, \oc8051_golden_model_1.DPH [5]);
  and (_10573_, _10572_, \oc8051_golden_model_1.DPH [6]);
  nand (_10574_, _10573_, \oc8051_golden_model_1.DPH [7]);
  or (_10575_, _10573_, \oc8051_golden_model_1.DPH [7]);
  and (_10576_, _10575_, _10540_);
  and (_10577_, _10576_, _10574_);
  or (_10578_, _10577_, _10544_);
  or (_10579_, _10578_, _10542_);
  not (_10580_, _10145_);
  or (_10581_, _10543_, _06977_);
  and (_10582_, _10581_, _10580_);
  and (_10583_, _10582_, _10579_);
  or (_10584_, _10583_, _10149_);
  nor (_10585_, _08471_, _08464_);
  and (_10586_, _10585_, _10584_);
  not (_10587_, _10585_);
  and (_10588_, _10587_, _10003_);
  nor (_10589_, _08478_, _03957_);
  not (_10590_, _10589_);
  or (_10591_, _10590_, _10588_);
  or (_10592_, _10591_, _10586_);
  or (_10593_, _10589_, _06977_);
  and (_10594_, _10593_, _04703_);
  and (_10595_, _10594_, _10592_);
  and (_10596_, _06967_, _03838_);
  nor (_10597_, _03959_, _03486_);
  not (_10598_, _10597_);
  or (_10599_, _10598_, _10596_);
  or (_10600_, _10599_, _10595_);
  and (_10601_, _03485_, _03383_);
  not (_10602_, _10601_);
  or (_10603_, _10597_, _06977_);
  and (_10604_, _10603_, _10602_);
  and (_10605_, _10604_, _10600_);
  or (_10606_, _10143_, _10146_);
  or (_10607_, _08783_, _06977_);
  and (_10608_, _10607_, _10601_);
  and (_10609_, _10608_, _10606_);
  or (_10610_, _10609_, _10605_);
  and (_10611_, _03476_, _03316_);
  nor (_10612_, _08502_, _10611_);
  and (_10613_, _10612_, _10610_);
  nor (_10614_, _08508_, _03965_);
  not (_10615_, _10614_);
  not (_10616_, _10612_);
  and (_10617_, _10616_, _10003_);
  or (_10618_, _10617_, _10615_);
  or (_10619_, _10618_, _10613_);
  or (_10620_, _10614_, _06977_);
  and (_10621_, _10620_, _04708_);
  and (_10622_, _10621_, _10619_);
  not (_10623_, _10031_);
  and (_10624_, _06967_, _03866_);
  or (_10625_, _10624_, _10623_);
  or (_10626_, _10625_, _10622_);
  and (_10627_, _10626_, _10033_);
  not (_10628_, _10027_);
  or (_10629_, _10143_, \oc8051_golden_model_1.PSW [7]);
  or (_10630_, _06977_, _08059_);
  and (_10631_, _10630_, _10029_);
  and (_10632_, _10631_, _10629_);
  or (_10633_, _10632_, _10628_);
  or (_10634_, _10633_, _10627_);
  and (_10635_, _10634_, _10028_);
  or (_10636_, _10635_, _08528_);
  or (_10637_, _08527_, _06977_);
  and (_10638_, _10637_, _06532_);
  and (_10639_, _10638_, _10636_);
  not (_10640_, _10016_);
  and (_10641_, _06967_, _03835_);
  or (_10642_, _10641_, _10640_);
  or (_10644_, _10642_, _10639_);
  and (_10645_, _10644_, _10018_);
  not (_10646_, _10012_);
  or (_10647_, _10143_, _08059_);
  or (_10648_, _06977_, \oc8051_golden_model_1.PSW [7]);
  and (_10649_, _10648_, _10014_);
  and (_10650_, _10649_, _10647_);
  or (_10651_, _10650_, _10646_);
  or (_10652_, _10651_, _10645_);
  and (_10653_, _10652_, _10013_);
  or (_10655_, _10653_, _10011_);
  or (_10656_, _10010_, _06977_);
  and (_10657_, _10656_, _08007_);
  and (_10658_, _10657_, _10655_);
  and (_10659_, _10003_, _08006_);
  or (_10660_, _10659_, _03974_);
  or (_10661_, _10660_, _10658_);
  nand (_10662_, _05498_, _03974_);
  and (_10663_, _10662_, _10661_);
  or (_10664_, _10663_, _03474_);
  or (_10666_, _06977_, _06543_);
  and (_10667_, _10666_, _04386_);
  and (_10668_, _10667_, _10664_);
  not (_10669_, _10008_);
  and (_10670_, _06110_, \oc8051_golden_model_1.P0INREG [2]);
  and (_10671_, _06112_, \oc8051_golden_model_1.P1INREG [2]);
  nor (_10672_, _10671_, _10670_);
  and (_10673_, _06099_, \oc8051_golden_model_1.SCON [2]);
  and (_10674_, _06101_, \oc8051_golden_model_1.IE [2]);
  nor (_10675_, _10674_, _10673_);
  and (_10677_, _06089_, \oc8051_golden_model_1.IP [2]);
  and (_10678_, _06086_, \oc8051_golden_model_1.ACC [2]);
  nor (_10679_, _10678_, _10677_);
  and (_10680_, _06092_, \oc8051_golden_model_1.PSW [2]);
  and (_10681_, _06094_, \oc8051_golden_model_1.B [2]);
  nor (_10682_, _10681_, _10680_);
  and (_10683_, _10682_, _10679_);
  and (_10684_, _06081_, \oc8051_golden_model_1.TCON [2]);
  and (_10685_, _06106_, \oc8051_golden_model_1.P3INREG [2]);
  and (_10686_, _06104_, \oc8051_golden_model_1.P2INREG [2]);
  or (_10688_, _10686_, _10685_);
  nor (_10689_, _10688_, _10684_);
  and (_10690_, _10689_, _10683_);
  and (_10691_, _10690_, _10675_);
  and (_10692_, _10691_, _10672_);
  and (_10693_, _10692_, _05698_);
  and (_10694_, _05409_, _04165_);
  not (_10695_, _10694_);
  nor (_10696_, _10695_, _10693_);
  and (_10697_, _05394_, _04165_);
  not (_10699_, _10697_);
  and (_10700_, _06081_, \oc8051_golden_model_1.TCON [1]);
  and (_10701_, _06086_, \oc8051_golden_model_1.ACC [1]);
  nor (_10702_, _10701_, _10700_);
  and (_10703_, _06092_, \oc8051_golden_model_1.PSW [1]);
  not (_10704_, _10703_);
  and (_10705_, _06089_, \oc8051_golden_model_1.IP [1]);
  and (_10706_, _06094_, \oc8051_golden_model_1.B [1]);
  nor (_10707_, _10706_, _10705_);
  and (_10708_, _10707_, _10704_);
  and (_10710_, _10708_, _10702_);
  and (_10711_, _06099_, \oc8051_golden_model_1.SCON [1]);
  and (_10712_, _06101_, \oc8051_golden_model_1.IE [1]);
  nor (_10713_, _10712_, _10711_);
  and (_10714_, _06104_, \oc8051_golden_model_1.P2INREG [1]);
  and (_10715_, _06106_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_10716_, _10715_, _10714_);
  and (_10717_, _06110_, \oc8051_golden_model_1.P0INREG [1]);
  and (_10718_, _06112_, \oc8051_golden_model_1.P1INREG [1]);
  nor (_10719_, _10718_, _10717_);
  and (_10720_, _10719_, _10716_);
  and (_10721_, _10720_, _10713_);
  and (_10722_, _10721_, _10710_);
  and (_10723_, _10722_, _05601_);
  nor (_10724_, _10723_, _10699_);
  nor (_10725_, _10724_, _10696_);
  and (_10726_, _06089_, \oc8051_golden_model_1.IP [4]);
  and (_10727_, _06094_, \oc8051_golden_model_1.B [4]);
  nor (_10728_, _10727_, _10726_);
  and (_10729_, _06092_, \oc8051_golden_model_1.PSW [4]);
  and (_10730_, _06086_, \oc8051_golden_model_1.ACC [4]);
  nor (_10731_, _10730_, _10729_);
  and (_10732_, _10731_, _10728_);
  and (_10733_, _06081_, \oc8051_golden_model_1.TCON [4]);
  and (_10734_, _06106_, \oc8051_golden_model_1.P3INREG [4]);
  and (_10735_, _06104_, \oc8051_golden_model_1.P2INREG [4]);
  or (_10736_, _10735_, _10734_);
  nor (_10737_, _10736_, _10733_);
  and (_10738_, _06099_, \oc8051_golden_model_1.SCON [4]);
  and (_10739_, _06101_, \oc8051_golden_model_1.IE [4]);
  nor (_10740_, _10739_, _10738_);
  and (_10741_, _06110_, \oc8051_golden_model_1.P0INREG [4]);
  and (_10742_, _06112_, \oc8051_golden_model_1.P1INREG [4]);
  nor (_10743_, _10742_, _10741_);
  and (_10744_, _10743_, _10740_);
  and (_10745_, _10744_, _10737_);
  and (_10746_, _10745_, _10732_);
  and (_10747_, _10746_, _05899_);
  and (_10748_, _05341_, _05174_);
  not (_10749_, _10748_);
  nor (_10750_, _10749_, _10747_);
  nor (_10751_, _10750_, _06267_);
  and (_10752_, _10751_, _10725_);
  and (_10753_, _05341_, _04165_);
  not (_10754_, _10753_);
  not (_10755_, _05651_);
  and (_10756_, _06081_, \oc8051_golden_model_1.TCON [0]);
  and (_10757_, _06094_, \oc8051_golden_model_1.B [0]);
  nor (_10758_, _10757_, _10756_);
  and (_10759_, _06089_, \oc8051_golden_model_1.IP [0]);
  not (_10760_, _10759_);
  and (_10761_, _06092_, \oc8051_golden_model_1.PSW [0]);
  and (_10762_, _06086_, \oc8051_golden_model_1.ACC [0]);
  nor (_10763_, _10762_, _10761_);
  and (_10764_, _10763_, _10760_);
  and (_10765_, _10764_, _10758_);
  and (_10766_, _06099_, \oc8051_golden_model_1.SCON [0]);
  and (_10767_, _06101_, \oc8051_golden_model_1.IE [0]);
  nor (_10768_, _10767_, _10766_);
  and (_10769_, _06104_, \oc8051_golden_model_1.P2INREG [0]);
  and (_10770_, _06106_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_10771_, _10770_, _10769_);
  and (_10772_, _06110_, \oc8051_golden_model_1.P0INREG [0]);
  and (_10773_, _06112_, \oc8051_golden_model_1.P1INREG [0]);
  nor (_10774_, _10773_, _10772_);
  and (_10775_, _10774_, _10771_);
  and (_10776_, _10775_, _10768_);
  and (_10777_, _10776_, _10765_);
  and (_10778_, _10777_, _10755_);
  nor (_10779_, _10778_, _10754_);
  and (_10780_, _06081_, \oc8051_golden_model_1.TCON [6]);
  and (_10781_, _06094_, \oc8051_golden_model_1.B [6]);
  nor (_10782_, _10781_, _10780_);
  and (_10783_, _06089_, \oc8051_golden_model_1.IP [6]);
  not (_10784_, _10783_);
  and (_10785_, _06092_, \oc8051_golden_model_1.PSW [6]);
  and (_10786_, _06086_, \oc8051_golden_model_1.ACC [6]);
  nor (_10787_, _10786_, _10785_);
  and (_10788_, _10787_, _10784_);
  and (_10789_, _10788_, _10782_);
  and (_10790_, _06099_, \oc8051_golden_model_1.SCON [6]);
  and (_10791_, _06101_, \oc8051_golden_model_1.IE [6]);
  nor (_10792_, _10791_, _10790_);
  and (_10793_, _06104_, \oc8051_golden_model_1.P2INREG [6]);
  and (_10794_, _06106_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_10795_, _10794_, _10793_);
  and (_10796_, _06110_, \oc8051_golden_model_1.P0INREG [6]);
  and (_10797_, _06112_, \oc8051_golden_model_1.P1INREG [6]);
  nor (_10798_, _10797_, _10796_);
  and (_10799_, _10798_, _10795_);
  and (_10800_, _10799_, _10792_);
  and (_10801_, _10800_, _10789_);
  and (_10802_, _10801_, _06014_);
  and (_10803_, _05409_, _05174_);
  not (_10804_, _10803_);
  nor (_10805_, _10804_, _10802_);
  nor (_10806_, _10805_, _10779_);
  and (_10807_, _06081_, \oc8051_golden_model_1.TCON [3]);
  and (_10808_, _06086_, \oc8051_golden_model_1.ACC [3]);
  nor (_10809_, _10808_, _10807_);
  and (_10810_, _06092_, \oc8051_golden_model_1.PSW [3]);
  not (_10811_, _10810_);
  and (_10812_, _06089_, \oc8051_golden_model_1.IP [3]);
  and (_10813_, _06094_, \oc8051_golden_model_1.B [3]);
  nor (_10814_, _10813_, _10812_);
  and (_10815_, _10814_, _10811_);
  and (_10816_, _10815_, _10809_);
  and (_10817_, _06099_, \oc8051_golden_model_1.SCON [3]);
  and (_10818_, _06101_, \oc8051_golden_model_1.IE [3]);
  nor (_10819_, _10818_, _10817_);
  and (_10820_, _06104_, \oc8051_golden_model_1.P2INREG [3]);
  and (_10821_, _06106_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_10822_, _10821_, _10820_);
  and (_10823_, _06110_, \oc8051_golden_model_1.P0INREG [3]);
  and (_10824_, _06112_, \oc8051_golden_model_1.P1INREG [3]);
  nor (_10825_, _10824_, _10823_);
  and (_10826_, _10825_, _10822_);
  and (_10827_, _10826_, _10819_);
  and (_10828_, _10827_, _10816_);
  and (_10829_, _10828_, _05552_);
  and (_10830_, _05388_, _04165_);
  not (_10831_, _10830_);
  nor (_10832_, _10831_, _10829_);
  and (_10833_, _06110_, \oc8051_golden_model_1.P0INREG [5]);
  and (_10834_, _06112_, \oc8051_golden_model_1.P1INREG [5]);
  nor (_10835_, _10834_, _10833_);
  and (_10836_, _06099_, \oc8051_golden_model_1.SCON [5]);
  and (_10837_, _06101_, \oc8051_golden_model_1.IE [5]);
  nor (_10838_, _10837_, _10836_);
  and (_10839_, _06089_, \oc8051_golden_model_1.IP [5]);
  and (_10840_, _06086_, \oc8051_golden_model_1.ACC [5]);
  nor (_10841_, _10840_, _10839_);
  and (_10842_, _06092_, \oc8051_golden_model_1.PSW [5]);
  and (_10843_, _06094_, \oc8051_golden_model_1.B [5]);
  nor (_10844_, _10843_, _10842_);
  and (_10845_, _10844_, _10841_);
  and (_10846_, _06081_, \oc8051_golden_model_1.TCON [5]);
  and (_10847_, _06106_, \oc8051_golden_model_1.P3INREG [5]);
  and (_10848_, _06104_, \oc8051_golden_model_1.P2INREG [5]);
  or (_10849_, _10848_, _10847_);
  nor (_10850_, _10849_, _10846_);
  and (_10851_, _10850_, _10845_);
  and (_10852_, _10851_, _10838_);
  and (_10853_, _10852_, _10835_);
  and (_10854_, _10853_, _05800_);
  and (_10855_, _05394_, _05174_);
  not (_10856_, _10855_);
  nor (_10857_, _10856_, _10854_);
  nor (_10858_, _10857_, _10832_);
  and (_10859_, _10858_, _10806_);
  and (_10860_, _10859_, _10752_);
  not (_10861_, _10860_);
  or (_10862_, _10306_, _10861_);
  or (_10863_, _06967_, _10860_);
  and (_10864_, _10863_, _03831_);
  and (_10865_, _10864_, _10862_);
  or (_10866_, _10865_, _10669_);
  or (_10867_, _10866_, _10668_);
  and (_10868_, _10867_, _10009_);
  or (_10869_, _10868_, _09990_);
  not (_10870_, _07964_);
  or (_10871_, _09989_, _06977_);
  and (_10872_, _10871_, _10870_);
  and (_10873_, _10872_, _10869_);
  and (_10874_, _10003_, _07964_);
  or (_10875_, _10874_, _03707_);
  or (_10876_, _10875_, _10873_);
  nand (_10877_, _05498_, _03707_);
  and (_10878_, _10877_, _10876_);
  or (_10879_, _10878_, _03394_);
  or (_10880_, _06977_, _03395_);
  and (_10881_, _10880_, _03706_);
  and (_10882_, _10881_, _10879_);
  or (_10883_, _10306_, _10860_);
  nand (_10884_, _10300_, _10860_);
  and (_10885_, _10884_, _10883_);
  and (_10886_, _10885_, _03705_);
  and (_10887_, _06556_, _04728_);
  not (_10888_, _10887_);
  or (_10889_, _10888_, _10886_);
  or (_10890_, _10889_, _10882_);
  or (_10891_, _10887_, _10003_);
  and (_10892_, _10891_, _03704_);
  and (_10893_, _10892_, _10890_);
  nor (_10894_, _08777_, _08772_);
  nand (_10895_, _06977_, _03703_);
  nand (_10896_, _10895_, _10894_);
  or (_10897_, _10896_, _10893_);
  or (_10898_, _10003_, _10894_);
  and (_10899_, _10898_, _06956_);
  and (_10900_, _10899_, _10897_);
  and (_10901_, _03833_, _03638_);
  or (_10902_, _10901_, _03400_);
  or (_10903_, _10902_, _10900_);
  not (_10904_, _03400_);
  or (_10905_, _06977_, _10904_);
  and (_10906_, _10905_, _03385_);
  and (_10907_, _10906_, _10903_);
  and (_10908_, _10885_, _03384_);
  nand (_10909_, _03398_, _03316_);
  and (_10910_, _10909_, _04744_);
  not (_10911_, _10910_);
  or (_10912_, _10911_, _10908_);
  or (_10913_, _10912_, _10907_);
  or (_10914_, _10910_, _10003_);
  and (_10915_, _10914_, _03702_);
  and (_10916_, _10915_, _10913_);
  nor (_10917_, _08801_, _08794_);
  nand (_10918_, _06977_, _03701_);
  nand (_10919_, _10918_, _10917_);
  or (_10920_, _10919_, _10916_);
  not (_10921_, _03841_);
  or (_10922_, _10003_, _10917_);
  and (_10923_, _10922_, _10921_);
  and (_10924_, _10923_, _10920_);
  and (_10925_, _03841_, _03638_);
  or (_10926_, _10925_, _03399_);
  or (_10927_, _10926_, _10924_);
  and (_10928_, _03398_, _03383_);
  not (_10929_, _10928_);
  not (_10930_, _03399_);
  or (_10931_, _06977_, _10930_);
  and (_10932_, _10931_, _10929_);
  and (_10933_, _10932_, _10927_);
  and (_10934_, _10928_, _10003_);
  or (_10935_, _10934_, _10933_);
  or (_10936_, _10935_, _42912_);
  or (_10937_, _42908_, \oc8051_golden_model_1.PC [15]);
  and (_10938_, _10937_, _41654_);
  and (_40458_, _10938_, _10936_);
  not (_10939_, \oc8051_golden_model_1.P2 [7]);
  nor (_10940_, _42908_, _10939_);
  or (_10941_, _10940_, rst);
  nor (_10942_, _05380_, _10939_);
  not (_10943_, _05380_);
  nor (_10944_, _05498_, _10943_);
  or (_10945_, _10944_, _10942_);
  or (_10946_, _10945_, _06994_);
  nor (_10947_, _06104_, _10939_);
  and (_10948_, _06112_, \oc8051_golden_model_1.P1 [7]);
  and (_10949_, _06106_, \oc8051_golden_model_1.P3 [7]);
  nor (_10950_, _10949_, _10948_);
  and (_10951_, _06110_, \oc8051_golden_model_1.P0 [7]);
  and (_10952_, _06104_, \oc8051_golden_model_1.P2 [7]);
  nor (_10953_, _10952_, _10951_);
  and (_10954_, _10953_, _10950_);
  and (_10955_, _10954_, _06103_);
  and (_10956_, _10955_, _06098_);
  and (_10957_, _10956_, _05499_);
  nor (_10958_, _10957_, _05389_);
  and (_10959_, _10958_, _06104_);
  or (_10960_, _10959_, _10947_);
  and (_10961_, _10960_, _03691_);
  and (_10962_, _05380_, \oc8051_golden_model_1.P2 [7]);
  and (_10963_, _05382_, \oc8051_golden_model_1.P3 [7]);
  nor (_10964_, _10963_, _10962_);
  and (_10965_, _05372_, \oc8051_golden_model_1.P0 [7]);
  and (_10966_, _05376_, \oc8051_golden_model_1.P1 [7]);
  nor (_10967_, _10966_, _10965_);
  and (_10968_, _10967_, _10964_);
  and (_10969_, _10968_, _05368_);
  and (_10970_, _10969_, _05418_);
  and (_10971_, _10970_, _05444_);
  and (_10972_, _10971_, _05499_);
  not (_10973_, _10972_);
  and (_10974_, _05380_, \oc8051_golden_model_1.P2 [6]);
  and (_10975_, _05382_, \oc8051_golden_model_1.P3 [6]);
  nor (_10976_, _10975_, _10974_);
  and (_10977_, _05376_, \oc8051_golden_model_1.P1 [6]);
  and (_10978_, _05372_, \oc8051_golden_model_1.P0 [6]);
  nor (_10979_, _10978_, _10977_);
  and (_10980_, _10979_, _10976_);
  and (_10981_, _10980_, _05944_);
  and (_10982_, _10981_, _05924_);
  and (_10983_, _10982_, _05921_);
  and (_10984_, _10983_, _06014_);
  and (_10985_, _05380_, \oc8051_golden_model_1.P2 [5]);
  and (_10986_, _05382_, \oc8051_golden_model_1.P3 [5]);
  nor (_10987_, _10986_, _10985_);
  and (_10988_, _05372_, \oc8051_golden_model_1.P0 [5]);
  and (_10989_, _05376_, \oc8051_golden_model_1.P1 [5]);
  nor (_10990_, _10989_, _10988_);
  and (_10991_, _10990_, _10987_);
  and (_10992_, _10991_, _05709_);
  and (_10993_, _05722_, _05731_);
  nor (_10994_, _05714_, _05711_);
  nand (_10995_, _10994_, _05719_);
  nor (_10996_, _10995_, _05710_);
  and (_10997_, _10996_, _05743_);
  and (_10998_, _10997_, _10993_);
  and (_10999_, _10998_, _10992_);
  and (_11000_, _10999_, _05800_);
  and (_11001_, _05380_, \oc8051_golden_model_1.P2 [4]);
  and (_11002_, _05382_, \oc8051_golden_model_1.P3 [4]);
  nor (_11003_, _11002_, _11001_);
  and (_11004_, _05376_, \oc8051_golden_model_1.P1 [4]);
  and (_11005_, _05372_, \oc8051_golden_model_1.P0 [4]);
  nor (_11006_, _11005_, _11004_);
  and (_11007_, _11006_, _11003_);
  and (_11008_, _11007_, _05842_);
  and (_11009_, _11008_, _05822_);
  and (_11010_, _11009_, _05819_);
  and (_11011_, _11010_, _05899_);
  and (_11012_, _05548_, _05510_);
  and (_11013_, _05537_, _05530_);
  and (_11014_, _11013_, _05522_);
  not (_11015_, _05511_);
  and (_11016_, _05525_, _11015_);
  nor (_11017_, _05517_, _05512_);
  and (_11018_, _11017_, _11016_);
  and (_11019_, _05372_, \oc8051_golden_model_1.P0 [3]);
  and (_11020_, _05376_, \oc8051_golden_model_1.P1 [3]);
  nor (_11021_, _11020_, _11019_);
  and (_11022_, _05380_, \oc8051_golden_model_1.P2 [3]);
  and (_11023_, _05382_, \oc8051_golden_model_1.P3 [3]);
  nor (_11024_, _11023_, _11022_);
  and (_11025_, _11024_, _11021_);
  and (_11026_, _11025_, _11018_);
  and (_11027_, _11026_, _11014_);
  and (_11028_, _11027_, _11012_);
  and (_11029_, _11028_, _05552_);
  and (_11030_, _05694_, _05660_);
  and (_11031_, _05673_, _05682_);
  and (_11032_, _05380_, \oc8051_golden_model_1.P2 [2]);
  and (_11033_, _05382_, \oc8051_golden_model_1.P3 [2]);
  nor (_11034_, _11033_, _11032_);
  and (_11035_, _05372_, \oc8051_golden_model_1.P0 [2]);
  and (_11036_, _05376_, \oc8051_golden_model_1.P1 [2]);
  nor (_11037_, _11036_, _11035_);
  and (_11038_, _11037_, _11034_);
  not (_11039_, _05662_);
  and (_11040_, _11039_, _05670_);
  nor (_11041_, _05665_, _05661_);
  and (_11042_, _11041_, _11040_);
  and (_11043_, _11042_, _11038_);
  and (_11044_, _11043_, _11031_);
  and (_11045_, _11044_, _11030_);
  and (_11046_, _11045_, _05698_);
  and (_11047_, _05380_, \oc8051_golden_model_1.P2 [1]);
  and (_11048_, _05382_, \oc8051_golden_model_1.P3 [1]);
  nor (_11049_, _11048_, _11047_);
  and (_11050_, _05372_, \oc8051_golden_model_1.P0 [1]);
  and (_11051_, _05376_, \oc8051_golden_model_1.P1 [1]);
  nor (_11052_, _11051_, _11050_);
  and (_11053_, _11052_, _11049_);
  and (_11054_, _11053_, _05561_);
  and (_11055_, _11054_, _05585_);
  and (_11056_, _11055_, _05599_);
  and (_11057_, _11056_, _05601_);
  nor (_11058_, _05617_, _05613_);
  nand (_11059_, _11058_, _05625_);
  nor (_11060_, _11059_, _05614_);
  and (_11061_, _05622_, _05630_);
  and (_11062_, _11061_, _05637_);
  and (_11063_, _05372_, \oc8051_golden_model_1.P0 [0]);
  and (_11064_, _05376_, \oc8051_golden_model_1.P1 [0]);
  nor (_11065_, _11064_, _11063_);
  and (_11066_, _05380_, \oc8051_golden_model_1.P2 [0]);
  and (_11067_, _05382_, \oc8051_golden_model_1.P3 [0]);
  nor (_11068_, _11067_, _11066_);
  and (_11069_, _11068_, _11065_);
  and (_11070_, _11069_, _05612_);
  and (_11071_, _11070_, _11062_);
  and (_11072_, _11071_, _05646_);
  and (_11073_, _11072_, _11060_);
  and (_11074_, _11073_, _10755_);
  and (_11075_, _11074_, _11057_);
  and (_11076_, _11075_, _11046_);
  and (_11077_, _11076_, _11029_);
  and (_11078_, _11077_, _11011_);
  and (_11079_, _11078_, _11000_);
  and (_11080_, _11079_, _10984_);
  or (_11081_, _11080_, _10973_);
  nand (_11082_, _11080_, _10973_);
  and (_11083_, _11082_, _11081_);
  and (_11084_, _11083_, _05380_);
  or (_11085_, _11084_, _10942_);
  or (_11086_, _11085_, _04630_);
  and (_11087_, _05380_, \oc8051_golden_model_1.ACC [7]);
  or (_11088_, _11087_, _10942_);
  and (_11089_, _11088_, _04615_);
  nor (_11090_, _04615_, _10939_);
  or (_11091_, _11090_, _03757_);
  or (_11092_, _11091_, _11089_);
  and (_11093_, _11092_, _03697_);
  and (_11094_, _11093_, _11086_);
  nand (_11095_, _10957_, _06126_);
  and (_11096_, _11095_, _06104_);
  or (_11097_, _11096_, _10947_);
  and (_11098_, _11097_, _03696_);
  or (_11099_, _11098_, _03755_);
  or (_11100_, _11099_, _11094_);
  or (_11101_, _10945_, _04537_);
  and (_11102_, _11101_, _11100_);
  or (_11103_, _11102_, _03750_);
  or (_11104_, _11088_, _03751_);
  and (_11105_, _11104_, _03692_);
  and (_11106_, _11105_, _11103_);
  or (_11107_, _11106_, _10961_);
  and (_11108_, _11107_, _03685_);
  or (_11109_, _10957_, _06126_);
  or (_11110_, _11109_, _10947_);
  and (_11111_, _11097_, _03684_);
  and (_11112_, _11111_, _11110_);
  or (_11113_, _11112_, _11108_);
  and (_11114_, _11113_, _03680_);
  or (_11115_, _10958_, _06120_);
  and (_11116_, _11115_, _06104_);
  or (_11117_, _11116_, _10947_);
  and (_11118_, _11117_, _03679_);
  or (_11119_, _11118_, _07544_);
  or (_11120_, _11119_, _11114_);
  and (_11121_, _11120_, _10946_);
  or (_11122_, _11121_, _04678_);
  and (_11123_, _06237_, _05380_);
  or (_11124_, _10942_, _04679_);
  or (_11125_, _11124_, _11123_);
  and (_11126_, _11125_, _03415_);
  and (_11127_, _11126_, _11122_);
  and (_11128_, _06470_, \oc8051_golden_model_1.P1 [7]);
  and (_11129_, _06466_, \oc8051_golden_model_1.P0 [7]);
  and (_11130_, _06474_, \oc8051_golden_model_1.P2 [7]);
  and (_11131_, _06476_, \oc8051_golden_model_1.P3 [7]);
  or (_11132_, _11131_, _11130_);
  or (_11133_, _11132_, _11129_);
  or (_11134_, _11133_, _11128_);
  nor (_11135_, _11134_, _06464_);
  and (_11136_, _11135_, _06496_);
  and (_11137_, _11136_, _06462_);
  nand (_11138_, _11137_, _06447_);
  or (_11139_, _11138_, _06308_);
  and (_11140_, _11139_, _05380_);
  or (_11141_, _11140_, _10942_);
  and (_11142_, _11141_, _07559_);
  or (_11143_, _11142_, _08854_);
  or (_11144_, _11143_, _11127_);
  nand (_11145_, _10972_, _06070_);
  or (_11146_, _10972_, _06070_);
  and (_11147_, _11146_, _11145_);
  and (_11148_, _11147_, _05380_);
  or (_11149_, _10942_, _04703_);
  or (_11150_, _11149_, _11148_);
  and (_11151_, _06307_, _05380_);
  or (_11152_, _11151_, _10942_);
  or (_11153_, _11152_, _04694_);
  and (_11154_, _11153_, _04701_);
  and (_11155_, _11154_, _11150_);
  and (_11156_, _11155_, _11144_);
  nand (_11157_, _10972_, _06142_);
  or (_11158_, _10972_, _06142_);
  and (_11159_, _11158_, _11157_);
  and (_11160_, _11159_, _05380_);
  or (_11161_, _11160_, _10942_);
  and (_11162_, _11161_, _03959_);
  or (_11163_, _11162_, _11156_);
  and (_11164_, _11163_, _04708_);
  or (_11165_, _10973_, _10942_);
  and (_11166_, _11152_, _03866_);
  and (_11167_, _11166_, _11165_);
  or (_11168_, _11167_, _11164_);
  and (_11169_, _11168_, _04706_);
  and (_11170_, _11088_, _03967_);
  and (_11171_, _11170_, _11165_);
  or (_11172_, _11171_, _03835_);
  or (_11173_, _11172_, _11169_);
  and (_11174_, _11145_, _05380_);
  or (_11175_, _10942_, _06532_);
  or (_11176_, _11175_, _11174_);
  and (_11177_, _11176_, _06537_);
  and (_11178_, _11177_, _11173_);
  and (_11179_, _11157_, _05380_);
  or (_11180_, _11179_, _10942_);
  and (_11181_, _11180_, _03954_);
  or (_11182_, _11181_, _03703_);
  or (_11183_, _11182_, _11178_);
  or (_11184_, _11085_, _03704_);
  and (_11185_, _11184_, _03385_);
  and (_11186_, _11185_, _11183_);
  and (_11187_, _10960_, _03384_);
  or (_11188_, _11187_, _03701_);
  or (_11189_, _11188_, _11186_);
  not (_11190_, _10984_);
  not (_11191_, _11000_);
  not (_11192_, _11011_);
  not (_11193_, _11029_);
  not (_11194_, _11046_);
  nor (_11195_, _11074_, _11057_);
  and (_11196_, _11195_, _11194_);
  and (_11197_, _11196_, _11193_);
  and (_11198_, _11197_, _11192_);
  and (_11199_, _11198_, _11191_);
  nand (_11200_, _11199_, _11190_);
  nand (_11201_, _11200_, _10972_);
  or (_11202_, _11200_, _10972_);
  and (_11203_, _11202_, _11201_);
  and (_11204_, _11203_, _05380_);
  or (_11205_, _10942_, _03702_);
  or (_11206_, _11205_, _11204_);
  and (_11207_, _11206_, _42908_);
  and (_11208_, _11207_, _11189_);
  or (_40459_, _11208_, _10941_);
  not (_11209_, _05382_);
  and (_11210_, _11209_, \oc8051_golden_model_1.P3 [7]);
  nor (_11211_, _05498_, _11209_);
  or (_11212_, _11211_, _11210_);
  or (_11213_, _11212_, _06994_);
  not (_11214_, _06106_);
  and (_11215_, _11214_, \oc8051_golden_model_1.P3 [7]);
  and (_11216_, _10958_, _06106_);
  or (_11217_, _11216_, _11215_);
  and (_11218_, _11217_, _03691_);
  and (_11219_, _11083_, _05382_);
  or (_11220_, _11219_, _11210_);
  or (_11221_, _11220_, _04630_);
  and (_11222_, _05382_, \oc8051_golden_model_1.ACC [7]);
  or (_11223_, _11222_, _11210_);
  and (_11224_, _11223_, _04615_);
  and (_11225_, _04616_, \oc8051_golden_model_1.P3 [7]);
  or (_11226_, _11225_, _03757_);
  or (_11227_, _11226_, _11224_);
  and (_11228_, _11227_, _03697_);
  and (_11229_, _11228_, _11221_);
  and (_11230_, _11095_, _06106_);
  or (_11231_, _11230_, _11215_);
  and (_11232_, _11231_, _03696_);
  or (_11233_, _11232_, _03755_);
  or (_11234_, _11233_, _11229_);
  or (_11235_, _11212_, _04537_);
  and (_11236_, _11235_, _11234_);
  or (_11237_, _11236_, _03750_);
  or (_11238_, _11223_, _03751_);
  and (_11239_, _11238_, _03692_);
  and (_11240_, _11239_, _11237_);
  or (_11241_, _11240_, _11218_);
  and (_11242_, _11241_, _03685_);
  or (_11243_, _11215_, _11109_);
  and (_11244_, _11243_, _03684_);
  and (_11245_, _11244_, _11231_);
  or (_11246_, _11245_, _11242_);
  and (_11247_, _11246_, _03680_);
  and (_11248_, _11115_, _06106_);
  or (_11249_, _11248_, _11215_);
  and (_11250_, _11249_, _03679_);
  or (_11251_, _11250_, _07544_);
  or (_11252_, _11251_, _11247_);
  and (_11253_, _11252_, _11213_);
  or (_11254_, _11253_, _04678_);
  and (_11255_, _06237_, _05382_);
  or (_11256_, _11210_, _04679_);
  or (_11257_, _11256_, _11255_);
  and (_11258_, _11257_, _03415_);
  and (_11259_, _11258_, _11254_);
  and (_11260_, _11139_, _05382_);
  or (_11261_, _11260_, _11210_);
  and (_11262_, _11261_, _07559_);
  or (_11263_, _11262_, _08854_);
  or (_11264_, _11263_, _11259_);
  and (_11265_, _11147_, _05382_);
  or (_11266_, _11210_, _04703_);
  or (_11267_, _11266_, _11265_);
  and (_11268_, _06307_, _05382_);
  or (_11269_, _11268_, _11210_);
  or (_11270_, _11269_, _04694_);
  and (_11271_, _11270_, _04701_);
  and (_11272_, _11271_, _11267_);
  and (_11273_, _11272_, _11264_);
  and (_11274_, _11159_, _05382_);
  or (_11275_, _11274_, _11210_);
  and (_11276_, _11275_, _03959_);
  or (_11277_, _11276_, _11273_);
  and (_11278_, _11277_, _04708_);
  or (_11279_, _11210_, _10973_);
  and (_11280_, _11269_, _03866_);
  and (_11281_, _11280_, _11279_);
  or (_11282_, _11281_, _11278_);
  and (_11283_, _11282_, _04706_);
  and (_11284_, _11223_, _03967_);
  and (_11285_, _11284_, _11279_);
  or (_11286_, _11285_, _03835_);
  or (_11287_, _11286_, _11283_);
  and (_11288_, _11145_, _05382_);
  or (_11289_, _11210_, _06532_);
  or (_11290_, _11289_, _11288_);
  and (_11291_, _11290_, _06537_);
  and (_11292_, _11291_, _11287_);
  and (_11293_, _11157_, _05382_);
  or (_11294_, _11293_, _11210_);
  and (_11295_, _11294_, _03954_);
  or (_11296_, _11295_, _03703_);
  or (_11297_, _11296_, _11292_);
  or (_11298_, _11220_, _03704_);
  and (_11299_, _11298_, _03385_);
  and (_11300_, _11299_, _11297_);
  and (_11301_, _11217_, _03384_);
  or (_11302_, _11301_, _03701_);
  or (_11303_, _11302_, _11300_);
  and (_11304_, _11203_, _05382_);
  or (_11305_, _11210_, _03702_);
  or (_11306_, _11305_, _11304_);
  and (_11307_, _11306_, _42908_);
  and (_11308_, _11307_, _11303_);
  nor (_11309_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_11310_, _11309_, _05330_);
  or (_40461_, _11310_, _11308_);
  not (_11311_, _05372_);
  and (_11312_, _11311_, \oc8051_golden_model_1.P0 [7]);
  nor (_11313_, _05498_, _11311_);
  or (_11314_, _11313_, _11312_);
  or (_11315_, _11314_, _06994_);
  not (_11316_, _06110_);
  and (_11317_, _11316_, \oc8051_golden_model_1.P0 [7]);
  and (_11318_, _10958_, _06110_);
  or (_11319_, _11318_, _11317_);
  and (_11320_, _11319_, _03691_);
  and (_11321_, _11083_, _05372_);
  or (_11322_, _11321_, _11312_);
  or (_11323_, _11322_, _04630_);
  and (_11324_, _05372_, \oc8051_golden_model_1.ACC [7]);
  or (_11325_, _11324_, _11312_);
  and (_11326_, _11325_, _04615_);
  and (_11327_, _04616_, \oc8051_golden_model_1.P0 [7]);
  or (_11328_, _11327_, _03757_);
  or (_11329_, _11328_, _11326_);
  and (_11330_, _11329_, _03697_);
  and (_11331_, _11330_, _11323_);
  and (_11332_, _11095_, _06110_);
  or (_11333_, _11332_, _11317_);
  and (_11334_, _11333_, _03696_);
  or (_11335_, _11334_, _03755_);
  or (_11336_, _11335_, _11331_);
  or (_11337_, _11314_, _04537_);
  and (_11338_, _11337_, _11336_);
  or (_11339_, _11338_, _03750_);
  or (_11340_, _11325_, _03751_);
  and (_11341_, _11340_, _03692_);
  and (_11342_, _11341_, _11339_);
  or (_11343_, _11342_, _11320_);
  and (_11344_, _11343_, _03685_);
  or (_11345_, _11317_, _11109_);
  and (_11346_, _11345_, _03684_);
  and (_11347_, _11346_, _11333_);
  or (_11348_, _11347_, _11344_);
  and (_11349_, _11348_, _03680_);
  and (_11350_, _11115_, _06110_);
  or (_11351_, _11350_, _11317_);
  and (_11352_, _11351_, _03679_);
  or (_11353_, _11352_, _07544_);
  or (_11354_, _11353_, _11349_);
  and (_11355_, _11354_, _11315_);
  or (_11356_, _11355_, _04678_);
  and (_11357_, _06237_, _05372_);
  or (_11358_, _11312_, _04679_);
  or (_11359_, _11358_, _11357_);
  and (_11360_, _11359_, _03415_);
  and (_11361_, _11360_, _11356_);
  and (_11362_, _11139_, _05372_);
  or (_11363_, _11362_, _11312_);
  and (_11364_, _11363_, _07559_);
  or (_11365_, _11364_, _08854_);
  or (_11366_, _11365_, _11361_);
  and (_11367_, _11147_, _05372_);
  or (_11368_, _11312_, _04703_);
  or (_11369_, _11368_, _11367_);
  and (_11370_, _06307_, _05372_);
  or (_11371_, _11370_, _11312_);
  or (_11372_, _11371_, _04694_);
  and (_11373_, _11372_, _04701_);
  and (_11374_, _11373_, _11369_);
  and (_11375_, _11374_, _11366_);
  and (_11376_, _11159_, _05372_);
  or (_11377_, _11376_, _11312_);
  and (_11378_, _11377_, _03959_);
  or (_11379_, _11378_, _11375_);
  and (_11380_, _11379_, _04708_);
  or (_11381_, _11312_, _10973_);
  and (_11382_, _11371_, _03866_);
  and (_11383_, _11382_, _11381_);
  or (_11384_, _11383_, _11380_);
  and (_11385_, _11384_, _04706_);
  and (_11386_, _11325_, _03967_);
  and (_11387_, _11386_, _11381_);
  or (_11388_, _11387_, _03835_);
  or (_11389_, _11388_, _11385_);
  and (_11390_, _11145_, _05372_);
  or (_11391_, _11312_, _06532_);
  or (_11392_, _11391_, _11390_);
  and (_11393_, _11392_, _06537_);
  and (_11394_, _11393_, _11389_);
  and (_11395_, _11157_, _05372_);
  or (_11396_, _11395_, _11312_);
  and (_11397_, _11396_, _03954_);
  or (_11398_, _11397_, _03703_);
  or (_11399_, _11398_, _11394_);
  or (_11400_, _11322_, _03704_);
  and (_11401_, _11400_, _03385_);
  and (_11402_, _11401_, _11399_);
  and (_11403_, _11319_, _03384_);
  or (_11404_, _11403_, _03701_);
  or (_11405_, _11404_, _11402_);
  and (_11406_, _11203_, _05372_);
  or (_11407_, _11312_, _03702_);
  or (_11408_, _11407_, _11406_);
  and (_11409_, _11408_, _42908_);
  and (_11410_, _11409_, _11405_);
  nor (_11411_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_11412_, _11411_, _05330_);
  or (_40462_, _11412_, _11410_);
  not (_11413_, _05376_);
  and (_11414_, _11413_, \oc8051_golden_model_1.P1 [7]);
  nor (_11415_, _05498_, _11413_);
  or (_11416_, _11415_, _11414_);
  or (_11417_, _11416_, _06994_);
  not (_11418_, _06112_);
  and (_11419_, _11418_, \oc8051_golden_model_1.P1 [7]);
  and (_11420_, _10958_, _06112_);
  or (_11421_, _11420_, _11419_);
  and (_11422_, _11421_, _03691_);
  and (_11423_, _11083_, _05376_);
  or (_11424_, _11423_, _11414_);
  or (_11425_, _11424_, _04630_);
  and (_11426_, _05376_, \oc8051_golden_model_1.ACC [7]);
  or (_11427_, _11426_, _11414_);
  and (_11428_, _11427_, _04615_);
  and (_11429_, _04616_, \oc8051_golden_model_1.P1 [7]);
  or (_11430_, _11429_, _03757_);
  or (_11431_, _11430_, _11428_);
  and (_11432_, _11431_, _03697_);
  and (_11433_, _11432_, _11425_);
  and (_11434_, _11095_, _06112_);
  or (_11435_, _11434_, _11419_);
  and (_11436_, _11435_, _03696_);
  or (_11437_, _11436_, _03755_);
  or (_11438_, _11437_, _11433_);
  or (_11439_, _11416_, _04537_);
  and (_11440_, _11439_, _11438_);
  or (_11441_, _11440_, _03750_);
  or (_11442_, _11427_, _03751_);
  and (_11443_, _11442_, _03692_);
  and (_11444_, _11443_, _11441_);
  or (_11445_, _11444_, _11422_);
  and (_11446_, _11445_, _03685_);
  or (_11447_, _11419_, _11109_);
  and (_11448_, _11435_, _03684_);
  and (_11449_, _11448_, _11447_);
  or (_11450_, _11449_, _11446_);
  and (_11451_, _11450_, _03680_);
  and (_11452_, _11115_, _06112_);
  or (_11453_, _11452_, _11419_);
  and (_11454_, _11453_, _03679_);
  or (_11455_, _11454_, _07544_);
  or (_11456_, _11455_, _11451_);
  and (_11457_, _11456_, _11417_);
  or (_11458_, _11457_, _04678_);
  and (_11459_, _06237_, _05376_);
  or (_11460_, _11414_, _04679_);
  or (_11461_, _11460_, _11459_);
  and (_11462_, _11461_, _03415_);
  and (_11463_, _11462_, _11458_);
  and (_11464_, _11139_, _05376_);
  or (_11465_, _11464_, _11414_);
  and (_11466_, _11465_, _07559_);
  or (_11467_, _11466_, _08854_);
  or (_11468_, _11467_, _11463_);
  and (_11469_, _11147_, _05376_);
  or (_11470_, _11414_, _04703_);
  or (_11471_, _11470_, _11469_);
  and (_11472_, _06307_, _05376_);
  or (_11473_, _11472_, _11414_);
  or (_11474_, _11473_, _04694_);
  and (_11475_, _11474_, _04701_);
  and (_11476_, _11475_, _11471_);
  and (_11477_, _11476_, _11468_);
  and (_11478_, _11159_, _05376_);
  or (_11479_, _11478_, _11414_);
  and (_11480_, _11479_, _03959_);
  or (_11481_, _11480_, _11477_);
  and (_11482_, _11481_, _04708_);
  or (_11483_, _11414_, _10973_);
  and (_11484_, _11473_, _03866_);
  and (_11485_, _11484_, _11483_);
  or (_11486_, _11485_, _11482_);
  and (_11487_, _11486_, _04706_);
  and (_11488_, _11427_, _03967_);
  and (_11489_, _11488_, _11483_);
  or (_11490_, _11489_, _03835_);
  or (_11491_, _11490_, _11487_);
  and (_11492_, _11145_, _05376_);
  or (_11493_, _11414_, _06532_);
  or (_11494_, _11493_, _11492_);
  and (_11495_, _11494_, _06537_);
  and (_11496_, _11495_, _11491_);
  and (_11497_, _11157_, _05376_);
  or (_11498_, _11497_, _11414_);
  and (_11499_, _11498_, _03954_);
  or (_11500_, _11499_, _03703_);
  or (_11501_, _11500_, _11496_);
  or (_11502_, _11424_, _03704_);
  and (_11503_, _11502_, _03385_);
  and (_11504_, _11503_, _11501_);
  and (_11505_, _11421_, _03384_);
  or (_11506_, _11505_, _03701_);
  or (_11507_, _11506_, _11504_);
  and (_11508_, _11203_, _05376_);
  or (_11509_, _11414_, _03702_);
  or (_11510_, _11509_, _11508_);
  and (_11511_, _11510_, _42908_);
  and (_11512_, _11511_, _11507_);
  nor (_11513_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_11514_, _11513_, _05330_);
  or (_40463_, _11514_, _11512_);
  not (_11515_, \oc8051_golden_model_1.SP [7]);
  nor (_11516_, _42908_, _11515_);
  and (_11517_, _05059_, \oc8051_golden_model_1.SP [4]);
  and (_11518_, _11517_, \oc8051_golden_model_1.SP [5]);
  and (_11519_, _11518_, \oc8051_golden_model_1.SP [6]);
  or (_11520_, _11519_, \oc8051_golden_model_1.SP [7]);
  nand (_11521_, _11519_, \oc8051_golden_model_1.SP [7]);
  and (_11522_, _11521_, _11520_);
  or (_11523_, _11522_, _04735_);
  nor (_11524_, _05434_, _11515_);
  and (_11525_, _06523_, _05434_);
  or (_11526_, _11525_, _11524_);
  and (_11527_, _11526_, _03959_);
  not (_11528_, _10510_);
  not (_11529_, _05434_);
  nor (_11530_, _05498_, _11529_);
  or (_11531_, _11524_, _04678_);
  or (_11532_, _11531_, _11530_);
  and (_11533_, _11532_, _11528_);
  not (_11534_, \oc8051_golden_model_1.SP [6]);
  not (_11535_, \oc8051_golden_model_1.SP [5]);
  not (_11536_, \oc8051_golden_model_1.SP [4]);
  and (_11537_, _06155_, _11536_);
  and (_11538_, _11537_, _11535_);
  and (_11539_, _11538_, _11534_);
  and (_11540_, _11539_, _03674_);
  or (_11541_, _11540_, \oc8051_golden_model_1.SP [7]);
  nand (_11542_, _11540_, \oc8051_golden_model_1.SP [7]);
  nand (_11543_, _11542_, _11541_);
  nand (_11544_, _11543_, _03755_);
  and (_11545_, _06250_, _05434_);
  or (_11546_, _11545_, _11524_);
  or (_11547_, _11546_, _04630_);
  and (_11548_, _05434_, \oc8051_golden_model_1.ACC [7]);
  or (_11549_, _11548_, _11524_);
  or (_11550_, _11549_, _04616_);
  or (_11551_, _04615_, \oc8051_golden_model_1.SP [7]);
  and (_11552_, _11551_, _04948_);
  and (_11553_, _11552_, _11550_);
  and (_11554_, _11522_, _04111_);
  or (_11555_, _11554_, _03757_);
  or (_11556_, _11555_, _11553_);
  and (_11557_, _11556_, _03445_);
  and (_11558_, _11557_, _11547_);
  and (_11559_, _11522_, _04933_);
  or (_11560_, _11559_, _03755_);
  or (_11561_, _11560_, _11558_);
  and (_11562_, _11561_, _11544_);
  or (_11563_, _11562_, _03750_);
  or (_11564_, _11549_, _03751_);
  and (_11565_, _11564_, _04759_);
  and (_11566_, _11565_, _11563_);
  and (_11567_, _11518_, \oc8051_golden_model_1.SP [0]);
  and (_11568_, _11567_, \oc8051_golden_model_1.SP [6]);
  or (_11569_, _11568_, \oc8051_golden_model_1.SP [7]);
  nand (_11570_, _11568_, \oc8051_golden_model_1.SP [7]);
  and (_11571_, _11570_, _11569_);
  nand (_11572_, _11571_, _03690_);
  nand (_11573_, _11572_, _04968_);
  or (_11574_, _11573_, _11566_);
  or (_11575_, _11522_, _04968_);
  and (_11576_, _11575_, _06994_);
  and (_11577_, _11576_, _11574_);
  or (_11578_, _11577_, _11533_);
  and (_11579_, _06237_, _05434_);
  or (_11580_, _11524_, _04679_);
  or (_11581_, _11580_, _11579_);
  and (_11582_, _11581_, _03415_);
  and (_11583_, _11582_, _11578_);
  nor (_11584_, _06501_, _11529_);
  or (_11585_, _11584_, _11524_);
  and (_11586_, _11585_, _07559_);
  or (_11587_, _11586_, _03839_);
  or (_11588_, _11587_, _11583_);
  and (_11589_, _06307_, _05434_);
  or (_11590_, _11589_, _11524_);
  or (_11591_, _11590_, _04694_);
  and (_11592_, _11591_, _11588_);
  or (_11593_, _11592_, _03483_);
  not (_11594_, _03483_);
  or (_11595_, _11522_, _11594_);
  and (_11596_, _11595_, _11593_);
  or (_11597_, _11596_, _03838_);
  and (_11598_, _06515_, _05434_);
  or (_11599_, _11524_, _04703_);
  or (_11600_, _11599_, _11598_);
  and (_11601_, _11600_, _04701_);
  and (_11602_, _11601_, _11597_);
  or (_11603_, _11602_, _11527_);
  and (_11604_, _11603_, _04708_);
  or (_11605_, _11524_, _05501_);
  and (_11606_, _11590_, _03866_);
  and (_11607_, _11606_, _11605_);
  or (_11608_, _11607_, _11604_);
  and (_11609_, _11608_, _10031_);
  and (_11610_, _11549_, _03967_);
  and (_11611_, _11610_, _11605_);
  and (_11612_, _11522_, _03477_);
  or (_11613_, _11612_, _03835_);
  or (_11614_, _11613_, _11611_);
  or (_11615_, _11614_, _11609_);
  nor (_11616_, _06514_, _11529_);
  or (_11617_, _11616_, _11524_);
  or (_11618_, _11617_, _06532_);
  and (_11619_, _11618_, _11615_);
  or (_11620_, _11619_, _03954_);
  not (_11621_, _03974_);
  nor (_11622_, _06522_, _11529_);
  or (_11623_, _11524_, _06537_);
  or (_11624_, _11623_, _11622_);
  and (_11625_, _11624_, _11621_);
  and (_11626_, _11625_, _11620_);
  or (_11627_, _11539_, \oc8051_golden_model_1.SP [7]);
  nand (_11628_, _11539_, \oc8051_golden_model_1.SP [7]);
  and (_11629_, _11628_, _11627_);
  and (_11630_, _11629_, _03974_);
  or (_11631_, _11630_, _03474_);
  or (_11632_, _11631_, _11626_);
  or (_11633_, _11522_, _06543_);
  and (_11634_, _11633_, _11632_);
  or (_11635_, _11634_, _03707_);
  or (_11636_, _11629_, _03708_);
  and (_11637_, _11636_, _03704_);
  and (_11638_, _11637_, _11635_);
  and (_11639_, _11546_, _03703_);
  or (_11640_, _11639_, _05156_);
  or (_11641_, _11640_, _11638_);
  and (_11642_, _11641_, _11523_);
  or (_11643_, _11642_, _03701_);
  and (_11644_, _06021_, _05434_);
  or (_11645_, _11524_, _03702_);
  or (_11646_, _11645_, _11644_);
  and (_11647_, _11646_, _42908_);
  and (_11648_, _11647_, _11643_);
  or (_11649_, _11648_, _11516_);
  and (_40464_, _11649_, _41654_);
  nor (_11650_, _42908_, _08059_);
  nor (_11651_, _06092_, _08059_);
  and (_11652_, _06119_, _06092_);
  or (_11653_, _11652_, _11651_);
  or (_11654_, _11653_, _03385_);
  nor (_11655_, _05360_, _08059_);
  and (_11656_, _06523_, _05360_);
  or (_11657_, _11656_, _11655_);
  and (_11658_, _11657_, _03959_);
  not (_11659_, _05360_);
  nor (_11660_, _06501_, _11659_);
  or (_11661_, _11660_, _11655_);
  and (_11662_, _11661_, _07559_);
  nor (_11663_, _05498_, _11659_);
  or (_11664_, _11663_, _11655_);
  or (_11665_, _11664_, _06994_);
  not (_11666_, _03810_);
  not (_11667_, _03811_);
  nor (_11668_, _10860_, _11667_);
  and (_11669_, _10431_, _08059_);
  nand (_11670_, _05553_, \oc8051_golden_model_1.ACC [3]);
  nor (_11671_, _05553_, \oc8051_golden_model_1.ACC [3]);
  nor (_11672_, _05699_, \oc8051_golden_model_1.ACC [2]);
  or (_11673_, _11672_, _11671_);
  and (_11674_, _11673_, _11670_);
  nor (_11675_, _05602_, \oc8051_golden_model_1.ACC [1]);
  nor (_11676_, _05652_, _03558_);
  nor (_11677_, _11676_, _08711_);
  or (_11678_, _11677_, _11675_);
  and (_11679_, _11678_, _10456_);
  or (_11680_, _11679_, _11674_);
  and (_11681_, _11680_, _10454_);
  nand (_11682_, _05801_, \oc8051_golden_model_1.ACC [5]);
  nor (_11683_, _05801_, \oc8051_golden_model_1.ACC [5]);
  nor (_11684_, _05900_, \oc8051_golden_model_1.ACC [4]);
  or (_11685_, _11684_, _11683_);
  and (_11686_, _11685_, _11682_);
  and (_11687_, _11686_, _10453_);
  nor (_11688_, _05500_, \oc8051_golden_model_1.ACC [7]);
  or (_11689_, _06015_, \oc8051_golden_model_1.ACC [6]);
  nor (_11690_, _11689_, _06523_);
  or (_11691_, _11690_, _11688_);
  or (_11692_, _11691_, _11687_);
  or (_11693_, _11692_, _11681_);
  nor (_11694_, _10462_, _04216_);
  and (_11695_, _11694_, _11693_);
  nor (_11696_, _04482_, \oc8051_golden_model_1.ACC [1]);
  and (_11697_, _04482_, \oc8051_golden_model_1.ACC [1]);
  and (_11698_, _04211_, \oc8051_golden_model_1.ACC [0]);
  nor (_11699_, _11698_, _11697_);
  or (_11700_, _11699_, _11696_);
  and (_11701_, _11700_, _10440_);
  nand (_11702_, _03669_, \oc8051_golden_model_1.ACC [3]);
  nor (_11703_, _03669_, \oc8051_golden_model_1.ACC [3]);
  nor (_11704_, _04165_, \oc8051_golden_model_1.ACC [2]);
  or (_11705_, _11704_, _11703_);
  and (_11706_, _11705_, _11702_);
  or (_11707_, _11706_, _11701_);
  and (_11708_, _11707_, _10438_);
  and (_11709_, _03638_, _06142_);
  or (_11710_, _03740_, \oc8051_golden_model_1.ACC [6]);
  nor (_11711_, _11710_, _08485_);
  or (_11712_, _11711_, _11709_);
  nand (_11713_, _04034_, \oc8051_golden_model_1.ACC [5]);
  nor (_11714_, _04034_, \oc8051_golden_model_1.ACC [5]);
  nor (_11715_, _04446_, \oc8051_golden_model_1.ACC [4]);
  or (_11716_, _11715_, _11714_);
  and (_11717_, _11716_, _11713_);
  and (_11718_, _11717_, _10437_);
  or (_11719_, _11718_, _11712_);
  or (_11720_, _11719_, _11708_);
  not (_11721_, _03847_);
  nor (_11722_, _10446_, _11721_);
  and (_11723_, _11722_, _11720_);
  or (_11724_, _11723_, _11695_);
  or (_11725_, _11724_, _11669_);
  and (_11726_, _10418_, _10414_);
  or (_11727_, _10415_, _11726_);
  and (_11728_, _11727_, _10413_);
  and (_11729_, _10410_, _10408_);
  or (_11730_, _11729_, _10407_);
  or (_11731_, _11730_, _11728_);
  and (_11732_, _11731_, _10406_);
  or (_11733_, _10402_, _10399_);
  and (_11734_, _10397_, _11733_);
  and (_11735_, _11734_, _10398_);
  and (_11736_, _10395_, _05499_);
  or (_11737_, _11736_, _10392_);
  or (_11738_, _11737_, _11735_);
  or (_11739_, _11738_, _11732_);
  nor (_11740_, _10423_, _10388_);
  and (_11741_, _11740_, _11739_);
  and (_11742_, _11653_, _03691_);
  and (_11743_, _06250_, _05360_);
  or (_11744_, _11743_, _11655_);
  or (_11745_, _11744_, _04630_);
  not (_11746_, _08120_);
  and (_11747_, _05360_, \oc8051_golden_model_1.ACC [7]);
  or (_11748_, _11747_, _11655_);
  and (_11749_, _11748_, _04615_);
  nor (_11750_, _04615_, _08059_);
  or (_11751_, _11750_, _03757_);
  or (_11752_, _11751_, _11749_);
  and (_11753_, _11752_, _11746_);
  and (_11754_, _11753_, _11745_);
  nor (_11755_, _08131_, \oc8051_golden_model_1.PSW [7]);
  not (_11756_, _11755_);
  nor (_11757_, _11756_, _08141_);
  nor (_11758_, _11757_, _11746_);
  not (_11759_, _10353_);
  nand (_11760_, _11759_, _03761_);
  or (_11761_, _11760_, _11758_);
  or (_11762_, _11761_, _11754_);
  and (_11763_, _06127_, _06092_);
  or (_11764_, _11763_, _11651_);
  or (_11765_, _11764_, _03697_);
  or (_11766_, _11664_, _04537_);
  and (_11767_, _11766_, _11765_);
  and (_11768_, _11767_, _11762_);
  or (_11769_, _11768_, _03750_);
  or (_11770_, _11748_, _03751_);
  nor (_11771_, _10374_, _03691_);
  and (_11772_, _11771_, _11770_);
  and (_11773_, _11772_, _11769_);
  or (_11774_, _11773_, _11742_);
  and (_11775_, _11774_, _10388_);
  or (_11776_, _11775_, _11741_);
  and (_11777_, _11776_, _03855_);
  not (_11778_, _10175_);
  or (_11779_, _10177_, _11778_);
  and (_11780_, _11779_, _10172_);
  not (_11781_, _10169_);
  nand (_11782_, _10167_, _11781_);
  nand (_11783_, _11782_, _10166_);
  or (_11784_, _11783_, _11780_);
  and (_11785_, _11784_, _10165_);
  nand (_11786_, _10162_, _10159_);
  and (_11787_, _10157_, _11786_);
  and (_11788_, _11787_, _10158_);
  nand (_11789_, _10152_, _10154_);
  and (_11790_, _11789_, _06281_);
  or (_11791_, _11790_, _11788_);
  or (_11792_, _11791_, _11785_);
  nor (_11793_, _10181_, _03855_);
  and (_11794_, _11793_, _11792_);
  or (_11795_, _11794_, _11777_);
  and (_11796_, _11795_, _10433_);
  or (_11797_, _11796_, _11725_);
  and (_11798_, _11797_, _03778_);
  and (_11799_, _10860_, \oc8051_golden_model_1.PSW [7]);
  and (_11800_, _11799_, _03777_);
  or (_11801_, _11651_, _06268_);
  and (_11802_, _11801_, _03684_);
  and (_11803_, _11802_, _11764_);
  or (_11804_, _11803_, _11800_);
  or (_11805_, _11804_, _11798_);
  nor (_11806_, _07024_, _03811_);
  and (_11807_, _11806_, _11805_);
  or (_11808_, _11807_, _11668_);
  and (_11809_, _11808_, _11666_);
  nor (_11810_, _06992_, _03417_);
  or (_11811_, _10860_, \oc8051_golden_model_1.PSW [7]);
  and (_11812_, _11811_, _03810_);
  or (_11813_, _11812_, _11810_);
  or (_11814_, _11813_, _11809_);
  not (_11815_, _04276_);
  and (_11816_, _08186_, _06922_);
  and (_11817_, _08197_, _08193_);
  nor (_11818_, _11817_, _08191_);
  nand (_11819_, _08252_, _08193_);
  or (_11820_, _11819_, _08250_);
  and (_11821_, _11820_, _11818_);
  or (_11822_, _11821_, _11816_);
  and (_11823_, _11822_, _11815_);
  or (_11824_, _11823_, _08181_);
  and (_11825_, _11824_, _11814_);
  and (_11826_, _11822_, _04276_);
  or (_11827_, _11826_, _08260_);
  or (_11828_, _11827_, _11825_);
  and (_11829_, _08019_, _08014_);
  nor (_11830_, _11829_, _08012_);
  or (_11831_, _08021_, _08264_);
  or (_11832_, _11831_, _08278_);
  and (_11833_, _11832_, _11830_);
  and (_11834_, _08015_, _06933_);
  and (_11835_, _11834_, _06237_);
  or (_11836_, _08261_, _11835_);
  or (_11837_, _11836_, _11833_);
  and (_11838_, _11837_, _11828_);
  or (_11839_, _11838_, _03818_);
  and (_11840_, _08308_, _08302_);
  and (_11841_, _11840_, _06017_);
  and (_11842_, _08301_, _08297_);
  nor (_11843_, _11842_, _08295_);
  nand (_11844_, _08352_, _08297_);
  or (_11845_, _11844_, _08350_);
  and (_11846_, _11845_, _11843_);
  or (_11847_, _11846_, _11841_);
  or (_11848_, _11847_, _03823_);
  and (_11849_, _11848_, _08288_);
  and (_11850_, _11849_, _11839_);
  and (_11851_, _08363_, _05353_);
  and (_11852_, _08374_, _08371_);
  nor (_11853_, _11852_, _08369_);
  nand (_11854_, _08419_, _08371_);
  or (_11855_, _11854_, _08417_);
  and (_11856_, _11855_, _11853_);
  or (_11857_, _11856_, _11851_);
  and (_11858_, _11857_, _08287_);
  or (_11859_, _11858_, _07544_);
  or (_11860_, _11859_, _11850_);
  and (_11861_, _11860_, _11665_);
  or (_11862_, _11861_, _04678_);
  and (_11863_, _06237_, _05360_);
  or (_11864_, _11655_, _04679_);
  or (_11865_, _11864_, _11863_);
  and (_11866_, _11865_, _03415_);
  and (_11867_, _11866_, _11862_);
  or (_11868_, _11867_, _11662_);
  nor (_11869_, _07558_, _03746_);
  and (_11870_, _11869_, _11868_);
  nor (_11871_, _10860_, _08059_);
  and (_11872_, _11871_, _03746_);
  or (_11873_, _11872_, _03839_);
  or (_11874_, _11873_, _11870_);
  and (_11875_, _06307_, _05360_);
  or (_11876_, _11875_, _11655_);
  or (_11877_, _11876_, _04694_);
  and (_11878_, _11877_, _11874_);
  and (_11879_, _11878_, _04336_);
  nand (_11880_, _10860_, _08059_);
  and (_11881_, _11880_, _03745_);
  or (_11882_, _11881_, _11879_);
  or (_11883_, _11882_, _03838_);
  and (_11884_, _06515_, _05360_);
  or (_11885_, _11884_, _11655_);
  or (_11886_, _11885_, _04703_);
  and (_11887_, _11886_, _04701_);
  and (_11888_, _11887_, _11883_);
  or (_11889_, _11888_, _11658_);
  and (_11890_, _11889_, _04708_);
  or (_11891_, _11655_, _05501_);
  and (_11892_, _11876_, _03866_);
  and (_11893_, _11892_, _11891_);
  or (_11894_, _11893_, _11890_);
  and (_11895_, _11894_, _04706_);
  and (_11896_, _11748_, _03967_);
  and (_11897_, _11896_, _11891_);
  or (_11898_, _11897_, _03835_);
  or (_11899_, _11898_, _11895_);
  nor (_11900_, _06514_, _11659_);
  or (_11901_, _11655_, _06532_);
  or (_11902_, _11901_, _11900_);
  and (_11903_, _11902_, _06537_);
  and (_11904_, _11903_, _11899_);
  nor (_11905_, _06522_, _11659_);
  or (_11906_, _11905_, _11655_);
  and (_11907_, _11906_, _03954_);
  or (_11908_, _11907_, _08540_);
  or (_11909_, _11908_, _11904_);
  nor (_11910_, _08541_, _04374_);
  not (_11911_, _08540_);
  nor (_11912_, _08190_, _06142_);
  or (_11913_, _11912_, _08569_);
  or (_11914_, _11913_, _11816_);
  or (_11915_, _11914_, _11911_);
  and (_11916_, _11915_, _11910_);
  and (_11917_, _11916_, _11909_);
  not (_11918_, _11910_);
  and (_11919_, _11914_, _11918_);
  or (_11920_, _11919_, _08079_);
  or (_11921_, _11920_, _11917_);
  or (_11922_, _08080_, _11835_);
  nor (_11923_, _08011_, _06142_);
  or (_11924_, _11923_, _08076_);
  or (_11925_, _11924_, _11922_);
  and (_11926_, _11925_, _03964_);
  and (_11927_, _11926_, _11921_);
  nor (_11928_, _08294_, _06142_);
  or (_11929_, _11928_, _08603_);
  or (_11930_, _11929_, _11841_);
  and (_11931_, _11930_, _03963_);
  or (_11932_, _11931_, _08580_);
  or (_11933_, _11932_, _11927_);
  nor (_11934_, _08368_, _06142_);
  or (_11935_, _11934_, _08630_);
  or (_11936_, _11851_, _08581_);
  or (_11937_, _11936_, _11935_);
  and (_11938_, _11937_, _08007_);
  and (_11939_, _11938_, _11933_);
  nand (_11940_, _08006_, \oc8051_golden_model_1.ACC [7]);
  nand (_11941_, _11940_, _10007_);
  or (_11942_, _11941_, _11939_);
  and (_11943_, _08678_, _08468_);
  not (_11944_, _08082_);
  and (_11945_, _08648_, _11944_);
  or (_11946_, _10007_, _08467_);
  or (_11947_, _11946_, _11945_);
  or (_11948_, _11947_, _11943_);
  and (_11949_, _11948_, _11942_);
  or (_11950_, _11949_, _07966_);
  and (_11951_, _08000_, _07969_);
  not (_11952_, _07967_);
  or (_11953_, _07970_, _07968_);
  and (_11954_, _11953_, _11952_);
  or (_11955_, _11954_, _10004_);
  or (_11956_, _11955_, _11951_);
  and (_11957_, _11956_, _04166_);
  and (_11958_, _11957_, _11950_);
  not (_11959_, _06522_);
  not (_11960_, _06521_);
  nand (_11961_, _08724_, _11960_);
  and (_11962_, _11961_, _03709_);
  and (_11963_, _11962_, _11959_);
  or (_11964_, _11963_, _08691_);
  or (_11965_, _11964_, _11958_);
  not (_11966_, _08484_);
  or (_11967_, _08763_, _08483_);
  and (_11968_, _11967_, _08691_);
  nand (_11969_, _11968_, _11966_);
  and (_11970_, _11969_, _11965_);
  or (_11971_, _11970_, _03703_);
  not (_11972_, _08777_);
  or (_11973_, _11744_, _03704_);
  and (_11974_, _11973_, _11972_);
  and (_11975_, _11974_, _11971_);
  and (_11976_, _08777_, \oc8051_golden_model_1.ACC [0]);
  or (_11977_, _11976_, _03384_);
  or (_11978_, _11977_, _11975_);
  and (_11979_, _11978_, _11654_);
  or (_11980_, _11979_, _03701_);
  and (_11981_, _06021_, _05360_);
  or (_11982_, _11655_, _03702_);
  or (_11983_, _11982_, _11981_);
  and (_11984_, _11983_, _42908_);
  and (_11985_, _11984_, _11980_);
  or (_11986_, _11985_, _11650_);
  and (_40465_, _11986_, _41654_);
  and (_11987_, _42912_, \oc8051_golden_model_1.P0INREG [7]);
  or (_11988_, _11987_, _01289_);
  and (_40467_, _11988_, _41654_);
  and (_11989_, _42912_, \oc8051_golden_model_1.P1INREG [7]);
  or (_11990_, _11989_, _01381_);
  and (_40468_, _11990_, _41654_);
  and (_11991_, _42912_, \oc8051_golden_model_1.P2INREG [7]);
  or (_11992_, _11991_, _01125_);
  and (_40469_, _11992_, _41654_);
  and (_11993_, _42912_, \oc8051_golden_model_1.P3INREG [7]);
  or (_11994_, _11993_, _01055_);
  and (_40470_, _11994_, _41654_);
  nor (_11995_, _04994_, _04749_);
  nor (_11996_, _11995_, _04995_);
  nor (_11997_, _05173_, _04994_);
  nor (_11998_, _11997_, _05319_);
  and (_11999_, _11998_, _11996_);
  and (_12000_, _11999_, _04993_);
  or (_12001_, _12000_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_12002_, _05333_, _04915_);
  and (_12003_, _12002_, _05326_);
  and (_12004_, _12002_, _05329_);
  nor (_12005_, _12004_, _12003_);
  and (_12006_, _12005_, _04753_);
  and (_12007_, _12006_, _12002_);
  not (_12008_, _12007_);
  and (_12009_, _12008_, _12001_);
  not (_12010_, _12000_);
  nand (_12011_, _03400_, _03129_);
  nand (_12012_, _10458_, _06538_);
  and (_12013_, _05652_, _06428_);
  and (_12014_, _12013_, _04709_);
  or (_12015_, _04677_, _04608_);
  and (_12016_, _06935_, _05351_);
  or (_12017_, _12016_, _05650_);
  and (_12018_, _12017_, _04269_);
  or (_12019_, _05652_, _04759_);
  nor (_12020_, _10778_, _10753_);
  or (_12021_, _12020_, _06123_);
  nand (_12022_, _10320_, _04608_);
  nand (_12023_, _04111_, _03129_);
  or (_12024_, _04111_, \oc8051_golden_model_1.ACC [0]);
  and (_12025_, _12024_, _12023_);
  nor (_12026_, _12025_, _10320_);
  nor (_12027_, _12026_, _04631_);
  and (_12028_, _12027_, _12022_);
  nor (_12029_, _05652_, _04816_);
  or (_12030_, _12029_, _12028_);
  and (_12031_, _12030_, _06125_);
  nand (_12032_, _10778_, _10754_);
  and (_12033_, _12032_, _04629_);
  or (_12034_, _12033_, _04933_);
  or (_12035_, _12034_, _12031_);
  nor (_12036_, _03445_, \oc8051_golden_model_1.PC [0]);
  nor (_12037_, _12036_, _04640_);
  and (_12038_, _12037_, _12035_);
  and (_12039_, _04640_, _04608_);
  or (_12040_, _12039_, _03694_);
  or (_12041_, _12040_, _12038_);
  and (_12042_, _12041_, _12021_);
  or (_12043_, _12042_, _03690_);
  and (_12044_, _12043_, _12019_);
  or (_12045_, _12044_, _03687_);
  not (_12046_, _10779_);
  and (_12047_, _12032_, _12046_);
  or (_12048_, _12047_, _03688_);
  and (_12049_, _12048_, _03442_);
  and (_12050_, _12049_, _12045_);
  or (_12051_, _03442_, _03129_);
  nand (_12052_, _03807_, _12051_);
  or (_12053_, _12052_, _12050_);
  or (_12054_, _05652_, _03807_);
  and (_12055_, _12054_, _04663_);
  and (_12056_, _12055_, _12053_);
  or (_12057_, _12056_, _12018_);
  and (_12058_, _12057_, _05114_);
  and (_12059_, _10753_, \oc8051_golden_model_1.PSW [7]);
  nor (_12060_, _12059_, _12020_);
  nor (_12061_, _12060_, _05114_);
  or (_12062_, _12061_, _12058_);
  and (_12063_, _12062_, _03418_);
  or (_12064_, _03418_, _03129_);
  nand (_12065_, _04677_, _12064_);
  or (_12066_, _12065_, _12063_);
  and (_12067_, _12066_, _12015_);
  or (_12068_, _12067_, _04680_);
  not (_12069_, _04681_);
  not (_12070_, _04680_);
  or (_12071_, _06935_, _12070_);
  and (_12072_, _12071_, _12069_);
  and (_12073_, _12072_, _12068_);
  and (_12074_, _06070_, _04608_);
  and (_12075_, _06463_, \oc8051_golden_model_1.DPL [0]);
  and (_12076_, _06443_, \oc8051_golden_model_1.TL0 [0]);
  nor (_12077_, _12076_, _12075_);
  and (_12078_, _06491_, \oc8051_golden_model_1.DPH [0]);
  and (_12079_, _06434_, \oc8051_golden_model_1.TH1 [0]);
  nor (_12080_, _12079_, _12078_);
  and (_12081_, _12080_, _12077_);
  and (_12082_, _06412_, \oc8051_golden_model_1.B [0]);
  and (_12083_, _06409_, \oc8051_golden_model_1.ACC [0]);
  nor (_12084_, _12083_, _12082_);
  and (_12085_, _06420_, \oc8051_golden_model_1.IP [0]);
  and (_12086_, _06424_, \oc8051_golden_model_1.PSW [0]);
  nor (_12087_, _12086_, _12085_);
  and (_12088_, _12087_, _12084_);
  and (_12089_, _06482_, \oc8051_golden_model_1.IE [0]);
  and (_12090_, _06485_, \oc8051_golden_model_1.SBUF [0]);
  and (_12091_, _06487_, \oc8051_golden_model_1.SCON [0]);
  or (_12092_, _12091_, _12090_);
  nor (_12093_, _12092_, _12089_);
  and (_12094_, _12093_, _12088_);
  and (_12095_, _12094_, _12081_);
  and (_12096_, _06448_, \oc8051_golden_model_1.TH0 [0]);
  and (_12097_, _06452_, \oc8051_golden_model_1.TL1 [0]);
  nor (_12098_, _12097_, _12096_);
  and (_12099_, _06455_, \oc8051_golden_model_1.TCON [0]);
  and (_12100_, _06459_, \oc8051_golden_model_1.PCON [0]);
  nor (_12101_, _12100_, _12099_);
  and (_12102_, _12101_, _12098_);
  and (_12103_, _06470_, \oc8051_golden_model_1.P1INREG [0]);
  not (_12104_, _12103_);
  and (_12105_, _06466_, \oc8051_golden_model_1.P0INREG [0]);
  not (_12106_, _12105_);
  and (_12107_, _06474_, \oc8051_golden_model_1.P2INREG [0]);
  and (_12108_, _06476_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_12109_, _12108_, _12107_);
  and (_12110_, _12109_, _12106_);
  and (_12111_, _12110_, _12104_);
  and (_12112_, _06438_, \oc8051_golden_model_1.SP [0]);
  and (_12113_, _06493_, \oc8051_golden_model_1.TMOD [0]);
  nor (_12114_, _12113_, _12112_);
  and (_12115_, _12114_, _12111_);
  and (_12116_, _12115_, _12102_);
  and (_12117_, _12116_, _12095_);
  not (_12118_, _12117_);
  nor (_12119_, _12118_, _12074_);
  nor (_12120_, _12119_, _06296_);
  or (_12121_, _12120_, _06306_);
  or (_12122_, _12121_, _12073_);
  and (_12123_, _06306_, _04211_);
  nor (_12124_, _12123_, _04695_);
  and (_12125_, _12124_, _12122_);
  and (_12126_, _04695_, _06428_);
  or (_12127_, _12126_, _03483_);
  or (_12128_, _12127_, _12125_);
  and (_12129_, _03483_, _03129_);
  nor (_12130_, _12129_, _04704_);
  and (_12131_, _12130_, _12128_);
  nor (_12132_, _05652_, _06428_);
  nor (_12133_, _12132_, _12013_);
  nor (_12134_, _12133_, _04702_);
  nor (_12135_, _12134_, _04705_);
  or (_12136_, _12135_, _12131_);
  nand (_12137_, _10459_, _04702_);
  and (_12138_, _12137_, _06519_);
  and (_12139_, _12138_, _12136_);
  or (_12140_, _12139_, _12014_);
  and (_12141_, _12140_, _06030_);
  and (_12142_, _08712_, _04707_);
  or (_12143_, _12142_, _03477_);
  or (_12144_, _12143_, _12141_);
  and (_12145_, _03477_, _03129_);
  nor (_12146_, _12145_, _06533_);
  and (_12147_, _12146_, _12144_);
  nor (_12148_, _12132_, _06539_);
  or (_12149_, _12148_, _06538_);
  or (_12150_, _12149_, _12147_);
  and (_12151_, _12150_, _12012_);
  or (_12152_, _12151_, _03474_);
  nand (_12153_, _03474_, _03129_);
  and (_12154_, _12153_, _06556_);
  and (_12155_, _12154_, _12152_);
  nor (_12156_, _06556_, _04608_);
  or (_12157_, _12156_, _12155_);
  and (_12158_, _12157_, _04728_);
  and (_12159_, _06698_, _04727_);
  or (_12160_, _12159_, _04726_);
  or (_12161_, _12160_, _12158_);
  nand (_12162_, _05652_, _04726_);
  and (_12163_, _12162_, _06956_);
  and (_12164_, _12163_, _12161_);
  and (_12165_, _03833_, _03129_);
  or (_12166_, _12165_, _03400_);
  or (_12167_, _12166_, _12164_);
  and (_12168_, _12167_, _12011_);
  or (_12169_, _12168_, _03672_);
  or (_12170_, _12020_, _03673_);
  and (_12171_, _12170_, _10909_);
  and (_12172_, _12171_, _12169_);
  nor (_12173_, _10909_, _04608_);
  or (_12174_, _12173_, _12172_);
  and (_12175_, _12174_, _04744_);
  and (_12176_, _06698_, _04743_);
  or (_12177_, _12176_, _04742_);
  or (_12178_, _12177_, _12175_);
  nand (_12179_, _05652_, _04742_);
  and (_12180_, _12179_, _04993_);
  and (_12181_, _12180_, _12178_);
  or (_12182_, _12181_, _12010_);
  and (_12183_, _12182_, _12009_);
  and (_12184_, _05334_, _05326_);
  nor (_12185_, _12184_, _05335_);
  and (_12186_, _05334_, _04753_);
  and (_12187_, _12186_, _12185_);
  nand (_12188_, _10278_, _03833_);
  or (_12189_, _10116_, _03833_);
  and (_12190_, _12189_, _12188_);
  and (_12191_, _12190_, _05334_);
  and (_12192_, _12191_, _12187_);
  or (_40486_, _12192_, _12183_);
  or (_12193_, _12000_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_12194_, _12193_, _12008_);
  and (_12195_, _04223_, _03398_);
  not (_12196_, _12195_);
  nor (_12197_, _06936_, _06699_);
  or (_12198_, _12197_, _12196_);
  and (_12199_, _03803_, _03398_);
  nor (_12200_, _10723_, _10697_);
  or (_12201_, _12200_, _03673_);
  and (_12202_, _04223_, _03254_);
  not (_12203_, _12202_);
  and (_12204_, _03474_, _03100_);
  and (_12205_, _05602_, _04515_);
  nor (_12206_, _05602_, _04515_);
  nor (_12207_, _12206_, _12205_);
  and (_12208_, _12207_, _04704_);
  or (_12209_, _04813_, _04677_);
  nand (_12210_, _05602_, _03808_);
  not (_12211_, _10724_);
  nand (_12212_, _10723_, _10699_);
  and (_12213_, _12212_, _03687_);
  and (_12214_, _12213_, _12211_);
  or (_12215_, _12200_, _06123_);
  nor (_12216_, _06915_, _06131_);
  nand (_12217_, _12216_, _10320_);
  and (_12218_, _04111_, _03100_);
  or (_12219_, _04111_, _03491_);
  nand (_12220_, _12219_, _06140_);
  or (_12221_, _12220_, _12218_);
  and (_12222_, _12221_, _12217_);
  and (_12223_, _12222_, _04816_);
  not (_12224_, _05653_);
  and (_12225_, _06242_, _12224_);
  nor (_12226_, _12225_, _04816_);
  or (_12227_, _12226_, _12223_);
  or (_12228_, _12227_, _04629_);
  or (_12229_, _12212_, _06125_);
  and (_12230_, _12229_, _12228_);
  or (_12231_, _12230_, _04933_);
  nor (_12232_, _03445_, _03100_);
  nor (_12233_, _12232_, _04640_);
  and (_12234_, _12233_, _12231_);
  and (_12235_, _04813_, _04640_);
  or (_12236_, _12235_, _03694_);
  or (_12237_, _12236_, _12234_);
  and (_12238_, _12237_, _12215_);
  or (_12239_, _12238_, _03690_);
  nand (_12240_, _05602_, _03690_);
  and (_12241_, _12240_, _03688_);
  and (_12242_, _12241_, _12239_);
  or (_12243_, _12242_, _12214_);
  and (_12244_, _12243_, _03442_);
  or (_12245_, _03442_, \oc8051_golden_model_1.PC [1]);
  nand (_12246_, _03807_, _12245_);
  or (_12247_, _12246_, _12244_);
  and (_12248_, _12247_, _12210_);
  or (_12249_, _12248_, _04269_);
  and (_12250_, _06934_, _05351_);
  nand (_12251_, _05600_, _04269_);
  or (_12252_, _12251_, _12250_);
  and (_12253_, _12252_, _12249_);
  or (_12254_, _12253_, _04662_);
  and (_12255_, _10697_, \oc8051_golden_model_1.PSW [7]);
  nor (_12256_, _12255_, _12200_);
  nand (_12257_, _12256_, _04662_);
  and (_12258_, _12257_, _03418_);
  and (_12259_, _12258_, _12254_);
  or (_12260_, _03418_, \oc8051_golden_model_1.PC [1]);
  nand (_12261_, _04677_, _12260_);
  or (_12262_, _12261_, _12259_);
  and (_12263_, _12262_, _12209_);
  or (_12264_, _12263_, _04680_);
  or (_12265_, _06934_, _06297_);
  and (_12266_, _12265_, _06296_);
  and (_12267_, _12266_, _12264_);
  and (_12268_, _06070_, _04813_);
  and (_12269_, _06470_, \oc8051_golden_model_1.P1INREG [1]);
  not (_12270_, _12269_);
  and (_12271_, _06466_, \oc8051_golden_model_1.P0INREG [1]);
  not (_12272_, _12271_);
  and (_12273_, _06474_, \oc8051_golden_model_1.P2INREG [1]);
  and (_12274_, _06476_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_12275_, _12274_, _12273_);
  and (_12276_, _12275_, _12272_);
  and (_12277_, _12276_, _12270_);
  and (_12278_, _06438_, \oc8051_golden_model_1.SP [1]);
  and (_12279_, _06443_, \oc8051_golden_model_1.TL0 [1]);
  nor (_12280_, _12279_, _12278_);
  and (_12281_, _12280_, _12277_);
  and (_12282_, _06420_, \oc8051_golden_model_1.IP [1]);
  and (_12283_, _06412_, \oc8051_golden_model_1.B [1]);
  nor (_12284_, _12283_, _12282_);
  and (_12285_, _06424_, \oc8051_golden_model_1.PSW [1]);
  and (_12286_, _06409_, \oc8051_golden_model_1.ACC [1]);
  nor (_12287_, _12286_, _12285_);
  and (_12288_, _12287_, _12284_);
  and (_12289_, _06482_, \oc8051_golden_model_1.IE [1]);
  and (_12290_, _06485_, \oc8051_golden_model_1.SBUF [1]);
  and (_12291_, _06487_, \oc8051_golden_model_1.SCON [1]);
  or (_12292_, _12291_, _12290_);
  nor (_12293_, _12292_, _12289_);
  and (_12294_, _12293_, _12288_);
  and (_12295_, _12294_, _12281_);
  and (_12296_, _06448_, \oc8051_golden_model_1.TH0 [1]);
  and (_12297_, _06452_, \oc8051_golden_model_1.TL1 [1]);
  nor (_12298_, _12297_, _12296_);
  and (_12299_, _06455_, \oc8051_golden_model_1.TCON [1]);
  and (_12300_, _06459_, \oc8051_golden_model_1.PCON [1]);
  nor (_12301_, _12300_, _12299_);
  and (_12302_, _12301_, _12298_);
  and (_12303_, _06491_, \oc8051_golden_model_1.DPH [1]);
  and (_12304_, _06493_, \oc8051_golden_model_1.TMOD [1]);
  nor (_12305_, _12304_, _12303_);
  and (_12306_, _06463_, \oc8051_golden_model_1.DPL [1]);
  and (_12307_, _06434_, \oc8051_golden_model_1.TH1 [1]);
  nor (_12308_, _12307_, _12306_);
  and (_12309_, _12308_, _12305_);
  and (_12310_, _12309_, _12302_);
  and (_12311_, _12310_, _12295_);
  not (_12312_, _12311_);
  nor (_12313_, _12312_, _12268_);
  nor (_12314_, _12313_, _06296_);
  or (_12315_, _12314_, _06306_);
  or (_12316_, _12315_, _12267_);
  and (_12317_, _06306_, _04482_);
  nor (_12318_, _12317_, _04695_);
  and (_12319_, _12318_, _12316_);
  and (_12320_, _04695_, _06440_);
  or (_12321_, _12320_, _03483_);
  or (_12322_, _12321_, _12319_);
  and (_12323_, _03483_, \oc8051_golden_model_1.PC [1]);
  nor (_12324_, _12323_, _04704_);
  and (_12325_, _12324_, _12322_);
  or (_12326_, _12325_, _12208_);
  and (_12327_, _12326_, _06520_);
  and (_12328_, _08711_, _04702_);
  or (_12329_, _12328_, _12327_);
  and (_12330_, _12329_, _06519_);
  and (_12331_, _12206_, _04709_);
  or (_12332_, _12331_, _04707_);
  or (_12333_, _12332_, _12330_);
  or (_12334_, _08709_, _06030_);
  and (_12335_, _12334_, _12333_);
  or (_12336_, _12335_, _03477_);
  and (_12337_, _03477_, \oc8051_golden_model_1.PC [1]);
  nor (_12338_, _12337_, _06533_);
  and (_12339_, _12338_, _12336_);
  nor (_12340_, _12205_, _06539_);
  or (_12341_, _12340_, _06538_);
  or (_12342_, _12341_, _12339_);
  nand (_12343_, _08710_, _06538_);
  and (_12344_, _12343_, _06543_);
  and (_12345_, _12344_, _12342_);
  or (_12346_, _12345_, _12204_);
  and (_12347_, _12346_, _06550_);
  and (_12348_, _06554_, _06548_);
  not (_12349_, _12348_);
  nor (_12350_, _12216_, _06550_);
  or (_12351_, _12350_, _12349_);
  or (_12352_, _12351_, _12347_);
  nor (_12353_, _03420_, _03413_);
  and (_12354_, _12353_, _03254_);
  not (_12355_, _12354_);
  nand (_12356_, _12216_, _12349_);
  and (_12357_, _12356_, _12355_);
  and (_12358_, _12357_, _12352_);
  or (_12359_, _06936_, _06699_);
  and (_12360_, _12359_, _12354_);
  or (_12361_, _12360_, _12358_);
  and (_12362_, _12361_, _12203_);
  and (_12363_, _12359_, _12202_);
  or (_12364_, _12363_, _04726_);
  or (_12365_, _12364_, _12362_);
  nand (_12366_, _12225_, _04726_);
  and (_12367_, _12366_, _12365_);
  or (_12368_, _12367_, _03833_);
  nand (_12369_, _03833_, _10251_);
  and (_12370_, _12369_, _10904_);
  and (_12371_, _12370_, _12368_);
  and (_12372_, _03400_, _03100_);
  or (_12373_, _03672_, _12372_);
  or (_12374_, _12373_, _12371_);
  and (_12375_, _12374_, _12201_);
  or (_12376_, _12375_, _12199_);
  not (_12377_, _12199_);
  nor (_12378_, _12216_, _12377_);
  nor (_12379_, _12378_, _04904_);
  and (_12380_, _12379_, _12376_);
  and (_12381_, _12216_, _04904_);
  or (_12382_, _12381_, _05313_);
  or (_12383_, _12382_, _12380_);
  and (_12384_, _12353_, _03398_);
  not (_12385_, _12384_);
  not (_12386_, _12216_);
  nand (_12387_, _12386_, _05313_);
  and (_12388_, _12387_, _12385_);
  and (_12389_, _12388_, _12383_);
  and (_12390_, _12197_, _12384_);
  or (_12391_, _12390_, _12195_);
  or (_12392_, _12391_, _12389_);
  and (_12393_, _12392_, _12198_);
  or (_12394_, _12393_, _04742_);
  or (_12395_, _12225_, _04922_);
  and (_12396_, _12395_, _04993_);
  and (_12397_, _12396_, _12394_);
  or (_12398_, _12397_, _12010_);
  and (_12399_, _12398_, _12194_);
  nand (_12400_, _10218_, _03833_);
  or (_12401_, _10063_, _03833_);
  and (_12402_, _12401_, _12400_);
  and (_12403_, _12402_, _05334_);
  and (_12404_, _12403_, _12187_);
  or (_40487_, _12404_, _12399_);
  or (_12405_, _12000_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_12406_, _12405_, _12008_);
  nor (_12407_, _06936_, _06938_);
  nor (_12408_, _12407_, _08038_);
  or (_12409_, _12408_, _04744_);
  and (_12410_, _06131_, _05236_);
  nor (_12411_, _06131_, _05236_);
  nor (_12412_, _12411_, _12410_);
  nand (_12413_, _12412_, _06549_);
  nor (_12414_, _05699_, _04077_);
  and (_12415_, _12414_, _04709_);
  nand (_12416_, _05236_, _06291_);
  nand (_12417_, _05699_, _03808_);
  not (_12418_, _10696_);
  nand (_12419_, _10695_, _10693_);
  and (_12420_, _12419_, _03687_);
  and (_12421_, _12420_, _12418_);
  nor (_12422_, _10694_, _10693_);
  or (_12423_, _12422_, _06123_);
  or (_12424_, _06242_, _05700_);
  not (_12425_, _12424_);
  and (_12426_, _06242_, _05700_);
  nor (_12427_, _12426_, _12425_);
  nand (_12428_, _12427_, _04631_);
  nor (_12429_, _12412_, _06140_);
  and (_12430_, _04111_, _03405_);
  nor (_12431_, _04111_, _07740_);
  or (_12432_, _12431_, _12430_);
  and (_12433_, _12432_, _06140_);
  or (_12434_, _12433_, _04631_);
  or (_12435_, _12434_, _12429_);
  and (_12436_, _12435_, _06125_);
  and (_12437_, _12436_, _12428_);
  and (_12438_, _12419_, _04629_);
  or (_12439_, _12438_, _04933_);
  or (_12440_, _12439_, _12437_);
  nor (_12441_, _03445_, _03405_);
  nor (_12442_, _12441_, _04640_);
  and (_12443_, _12442_, _12440_);
  and (_12444_, _08217_, _04640_);
  or (_12445_, _12444_, _03694_);
  or (_12446_, _12445_, _12443_);
  and (_12447_, _12446_, _12423_);
  or (_12448_, _12447_, _03690_);
  nand (_12449_, _05699_, _03690_);
  and (_12450_, _12449_, _03688_);
  and (_12451_, _12450_, _12448_);
  or (_12452_, _12451_, _12421_);
  and (_12453_, _12452_, _03442_);
  or (_12454_, _03442_, _10089_);
  nand (_12455_, _03807_, _12454_);
  or (_12456_, _12455_, _12453_);
  and (_12457_, _12456_, _12417_);
  or (_12458_, _12457_, _04269_);
  and (_12459_, _06938_, _05351_);
  nand (_12460_, _05697_, _04269_);
  or (_12461_, _12460_, _12459_);
  and (_12462_, _12461_, _12458_);
  or (_12463_, _12462_, _04662_);
  and (_12464_, _10694_, \oc8051_golden_model_1.PSW [7]);
  nor (_12465_, _12464_, _12422_);
  nand (_12466_, _12465_, _04662_);
  and (_12467_, _12466_, _03418_);
  and (_12468_, _12467_, _12463_);
  or (_12469_, _03418_, _10089_);
  nand (_12470_, _04677_, _12469_);
  or (_12471_, _12470_, _12468_);
  and (_12472_, _12471_, _12416_);
  or (_12473_, _12472_, _04680_);
  or (_12474_, _06938_, _12070_);
  and (_12475_, _12474_, _12069_);
  and (_12476_, _12475_, _12473_);
  nor (_12477_, _06307_, _05236_);
  and (_12478_, _06420_, \oc8051_golden_model_1.IP [2]);
  and (_12479_, _06412_, \oc8051_golden_model_1.B [2]);
  nor (_12480_, _12479_, _12478_);
  and (_12481_, _06424_, \oc8051_golden_model_1.PSW [2]);
  and (_12482_, _06409_, \oc8051_golden_model_1.ACC [2]);
  nor (_12483_, _12482_, _12481_);
  and (_12484_, _12483_, _12480_);
  and (_12485_, _06482_, \oc8051_golden_model_1.IE [2]);
  and (_12486_, _06485_, \oc8051_golden_model_1.SBUF [2]);
  and (_12487_, _06487_, \oc8051_golden_model_1.SCON [2]);
  or (_12488_, _12487_, _12486_);
  nor (_12489_, _12488_, _12485_);
  and (_12490_, _06466_, \oc8051_golden_model_1.P0INREG [2]);
  not (_12491_, _12490_);
  and (_12492_, _06476_, \oc8051_golden_model_1.P3INREG [2]);
  and (_12493_, _06470_, \oc8051_golden_model_1.P1INREG [2]);
  and (_12494_, _06474_, \oc8051_golden_model_1.P2INREG [2]);
  or (_12495_, _12494_, _12493_);
  nor (_12496_, _12495_, _12492_);
  and (_12497_, _12496_, _12491_);
  and (_12498_, _12497_, _12489_);
  and (_12499_, _12498_, _12484_);
  and (_12500_, _06448_, \oc8051_golden_model_1.TH0 [2]);
  and (_12501_, _06452_, \oc8051_golden_model_1.TL1 [2]);
  nor (_12502_, _12501_, _12500_);
  and (_12503_, _06455_, \oc8051_golden_model_1.TCON [2]);
  and (_12504_, _06459_, \oc8051_golden_model_1.PCON [2]);
  nor (_12505_, _12504_, _12503_);
  and (_12506_, _12505_, _12502_);
  and (_12507_, _06491_, \oc8051_golden_model_1.DPH [2]);
  not (_12508_, _12507_);
  and (_12509_, _06434_, \oc8051_golden_model_1.TH1 [2]);
  and (_12510_, _06443_, \oc8051_golden_model_1.TL0 [2]);
  nor (_12511_, _12510_, _12509_);
  and (_12512_, _12511_, _12508_);
  and (_12513_, _06438_, \oc8051_golden_model_1.SP [2]);
  not (_12514_, _12513_);
  and (_12515_, _06463_, \oc8051_golden_model_1.DPL [2]);
  and (_12516_, _06493_, \oc8051_golden_model_1.TMOD [2]);
  nor (_12517_, _12516_, _12515_);
  and (_12518_, _12517_, _12514_);
  and (_12519_, _12518_, _12512_);
  and (_12520_, _12519_, _12506_);
  and (_12521_, _12520_, _12499_);
  not (_12522_, _12521_);
  nor (_12523_, _12522_, _12477_);
  nor (_12524_, _12523_, _06296_);
  or (_12525_, _12524_, _06306_);
  or (_12526_, _12525_, _12476_);
  and (_12527_, _06306_, _04165_);
  nor (_12528_, _12527_, _04695_);
  and (_12529_, _12528_, _12526_);
  and (_12530_, _04695_, _06457_);
  or (_12531_, _12530_, _03483_);
  or (_12532_, _12531_, _12529_);
  and (_12533_, _03483_, _10089_);
  nor (_12534_, _12533_, _04704_);
  and (_12535_, _12534_, _12532_);
  and (_12536_, _05699_, _04077_);
  nor (_12537_, _12536_, _12414_);
  nor (_12538_, _12537_, _04702_);
  nor (_12539_, _12538_, _04705_);
  or (_12540_, _12539_, _12535_);
  or (_12541_, _08707_, _06520_);
  and (_12542_, _12541_, _06519_);
  and (_12543_, _12542_, _12540_);
  or (_12544_, _12543_, _12415_);
  and (_12545_, _12544_, _06030_);
  and (_12546_, _08705_, _04707_);
  or (_12547_, _12546_, _03477_);
  or (_12548_, _12547_, _12545_);
  and (_12549_, _03477_, _10089_);
  nor (_12550_, _12549_, _06533_);
  and (_12551_, _12550_, _12548_);
  nor (_12552_, _12536_, _06539_);
  or (_12553_, _12552_, _06538_);
  or (_12554_, _12553_, _12551_);
  nand (_12555_, _08706_, _06538_);
  and (_12556_, _12555_, _06543_);
  and (_12557_, _12556_, _12554_);
  and (_12558_, _03474_, _03405_);
  or (_12559_, _06549_, _12558_);
  or (_12560_, _12559_, _12557_);
  nand (_12561_, _12560_, _12413_);
  and (_12562_, _12561_, _12348_);
  and (_12563_, _12412_, _12349_);
  or (_12564_, _12563_, _12354_);
  nor (_12565_, _12564_, _12562_);
  and (_12566_, _06699_, _06789_);
  nor (_12567_, _06699_, _06789_);
  nor (_12568_, _12567_, _12566_);
  nand (_12569_, _12568_, _04083_);
  and (_12570_, _12569_, _04727_);
  or (_12571_, _12570_, _12565_);
  nand (_12572_, _12568_, _12202_);
  and (_12573_, _12572_, _06562_);
  and (_12574_, _12573_, _12571_);
  nor (_12575_, _12427_, _06562_);
  or (_12576_, _12575_, _03833_);
  or (_12577_, _12576_, _12574_);
  nand (_12578_, _10249_, _03833_);
  and (_12579_, _12578_, _10904_);
  and (_12580_, _12579_, _12577_);
  and (_12581_, _03405_, _03400_);
  or (_12582_, _03672_, _12581_);
  or (_12583_, _12582_, _12580_);
  or (_12584_, _12422_, _03673_);
  and (_12585_, _12584_, _10909_);
  and (_12586_, _12585_, _12583_);
  not (_12587_, _10909_);
  nor (_12588_, _06915_, _08217_);
  nor (_12589_, _12588_, _08218_);
  and (_12590_, _12589_, _12587_);
  or (_12591_, _12590_, _04743_);
  or (_12592_, _12591_, _12586_);
  and (_12593_, _12592_, _12409_);
  or (_12594_, _12593_, _04742_);
  nor (_12595_, _05700_, _05653_);
  nor (_12596_, _12595_, _05701_);
  or (_12597_, _12596_, _04922_);
  and (_12598_, _12597_, _04993_);
  and (_12599_, _12598_, _12594_);
  or (_12600_, _12599_, _12010_);
  and (_12601_, _12600_, _12406_);
  nand (_12602_, _10211_, _03833_);
  or (_12603_, _10051_, _03833_);
  and (_12604_, _12603_, _12602_);
  and (_12605_, _12604_, _05334_);
  and (_12606_, _12605_, _12187_);
  or (_40489_, _12606_, _12601_);
  nor (_12607_, _12000_, _04998_);
  or (_12608_, _12607_, _12007_);
  and (_12609_, _12424_, _05554_);
  nor (_12610_, _12609_, _06245_);
  nor (_12611_, _12610_, _06562_);
  nor (_12612_, _12566_, _06744_);
  or (_12613_, _12612_, _06791_);
  and (_12614_, _12613_, _04727_);
  and (_12615_, _03516_, _03474_);
  nor (_12616_, _05553_, _03946_);
  and (_12617_, _12616_, _04709_);
  not (_12618_, _10832_);
  nand (_12619_, _10831_, _10829_);
  and (_12620_, _12619_, _03687_);
  and (_12621_, _12620_, _12618_);
  nor (_12622_, _10830_, _10829_);
  or (_12623_, _12622_, _06123_);
  or (_12624_, _12619_, _06125_);
  nor (_12625_, _12610_, _04816_);
  nor (_12626_, _12410_, _05050_);
  or (_12627_, _12626_, _06133_);
  or (_12628_, _12627_, _06140_);
  and (_12629_, _04111_, _03516_);
  nor (_12630_, _04111_, _07734_);
  or (_12631_, _12630_, _12629_);
  nor (_12632_, _12631_, _10320_);
  nor (_12633_, _12632_, _04631_);
  and (_12634_, _12633_, _12628_);
  or (_12635_, _12634_, _04629_);
  or (_12636_, _12635_, _12625_);
  and (_12637_, _12636_, _12624_);
  or (_12638_, _12637_, _04933_);
  nor (_12639_, _03516_, _03445_);
  nor (_12640_, _12639_, _04640_);
  and (_12641_, _12640_, _12638_);
  and (_12642_, _08216_, _04640_);
  or (_12643_, _12642_, _03694_);
  or (_12644_, _12643_, _12641_);
  and (_12645_, _12644_, _12623_);
  or (_12646_, _12645_, _03690_);
  nand (_12647_, _05553_, _03690_);
  and (_12648_, _12647_, _03688_);
  and (_12649_, _12648_, _12646_);
  or (_12650_, _12649_, _12621_);
  and (_12651_, _12650_, _03442_);
  or (_12652_, _03879_, _03442_);
  nand (_12653_, _03807_, _12652_);
  or (_12654_, _12653_, _12651_);
  nand (_12655_, _05553_, _03808_);
  and (_12657_, _12655_, _12654_);
  or (_12658_, _12657_, _04269_);
  and (_12659_, _06937_, _05351_);
  nand (_12660_, _05551_, _04269_);
  or (_12661_, _12660_, _12659_);
  and (_12662_, _12661_, _12658_);
  or (_12663_, _12662_, _04662_);
  and (_12664_, _10830_, \oc8051_golden_model_1.PSW [7]);
  nor (_12665_, _12622_, _12664_);
  nand (_12666_, _12665_, _04662_);
  and (_12667_, _12666_, _03418_);
  and (_12668_, _12667_, _12663_);
  or (_12669_, _03879_, _03418_);
  nand (_12670_, _04677_, _12669_);
  or (_12671_, _12670_, _12668_);
  nand (_12672_, _05050_, _06291_);
  and (_12673_, _12672_, _12671_);
  or (_12674_, _12673_, _04680_);
  or (_12675_, _06937_, _12070_);
  and (_12676_, _12675_, _12069_);
  and (_12678_, _12676_, _12674_);
  nor (_12679_, _06307_, _05050_);
  and (_12680_, _06470_, \oc8051_golden_model_1.P1INREG [3]);
  not (_12681_, _12680_);
  and (_12682_, _06466_, \oc8051_golden_model_1.P0INREG [3]);
  not (_12683_, _12682_);
  and (_12684_, _06474_, \oc8051_golden_model_1.P2INREG [3]);
  and (_12685_, _06476_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_12686_, _12685_, _12684_);
  and (_12687_, _12686_, _12683_);
  and (_12688_, _12687_, _12681_);
  and (_12689_, _06493_, \oc8051_golden_model_1.TMOD [3]);
  and (_12690_, _06443_, \oc8051_golden_model_1.TL0 [3]);
  nor (_12691_, _12690_, _12689_);
  and (_12692_, _12691_, _12688_);
  and (_12693_, _06482_, \oc8051_golden_model_1.IE [3]);
  and (_12694_, _06485_, \oc8051_golden_model_1.SBUF [3]);
  and (_12695_, _06487_, \oc8051_golden_model_1.SCON [3]);
  or (_12696_, _12695_, _12694_);
  nor (_12697_, _12696_, _12693_);
  and (_12698_, _06491_, \oc8051_golden_model_1.DPH [3]);
  and (_12699_, _06434_, \oc8051_golden_model_1.TH1 [3]);
  nor (_12700_, _12699_, _12698_);
  and (_12701_, _12700_, _12697_);
  and (_12702_, _12701_, _12692_);
  and (_12703_, _06412_, \oc8051_golden_model_1.B [3]);
  and (_12704_, _06409_, \oc8051_golden_model_1.ACC [3]);
  nor (_12705_, _12704_, _12703_);
  and (_12706_, _06420_, \oc8051_golden_model_1.IP [3]);
  and (_12707_, _06424_, \oc8051_golden_model_1.PSW [3]);
  nor (_12708_, _12707_, _12706_);
  and (_12709_, _12708_, _12705_);
  and (_12710_, _06438_, \oc8051_golden_model_1.SP [3]);
  and (_12711_, _06463_, \oc8051_golden_model_1.DPL [3]);
  nor (_12712_, _12711_, _12710_);
  and (_12713_, _12712_, _12709_);
  and (_12714_, _06455_, \oc8051_golden_model_1.TCON [3]);
  and (_12715_, _06448_, \oc8051_golden_model_1.TH0 [3]);
  nor (_12716_, _12715_, _12714_);
  and (_12717_, _06459_, \oc8051_golden_model_1.PCON [3]);
  and (_12718_, _06452_, \oc8051_golden_model_1.TL1 [3]);
  nor (_12719_, _12718_, _12717_);
  and (_12720_, _12719_, _12716_);
  and (_12721_, _12720_, _12713_);
  and (_12722_, _12721_, _12702_);
  not (_12723_, _12722_);
  nor (_12724_, _12723_, _12679_);
  nor (_12725_, _12724_, _06296_);
  or (_12726_, _12725_, _06306_);
  or (_12727_, _12726_, _12678_);
  and (_12728_, _06306_, _03669_);
  nor (_12729_, _12728_, _04695_);
  and (_12730_, _12729_, _12727_);
  and (_12731_, _04695_, _06415_);
  or (_12732_, _12731_, _03483_);
  or (_12733_, _12732_, _12730_);
  and (_12734_, _03879_, _03483_);
  nor (_12735_, _12734_, _04704_);
  and (_12736_, _12735_, _12733_);
  and (_12737_, _05553_, _03946_);
  nor (_12738_, _12737_, _12616_);
  nor (_12739_, _12738_, _04702_);
  nor (_12740_, _12739_, _04705_);
  or (_12741_, _12740_, _12736_);
  or (_12742_, _10455_, _06520_);
  and (_12743_, _12742_, _06519_);
  and (_12744_, _12743_, _12741_);
  or (_12745_, _12744_, _12617_);
  and (_12746_, _12745_, _06030_);
  and (_12747_, _08703_, _04707_);
  or (_12748_, _12747_, _03477_);
  or (_12749_, _12748_, _12746_);
  and (_12750_, _03879_, _03477_);
  nor (_12751_, _12750_, _06533_);
  and (_12752_, _12751_, _12749_);
  nor (_12753_, _12737_, _06539_);
  or (_12754_, _12753_, _06538_);
  or (_12755_, _12754_, _12752_);
  nand (_12756_, _08701_, _06538_);
  and (_12757_, _12756_, _06543_);
  and (_12758_, _12757_, _12755_);
  or (_12759_, _12758_, _12615_);
  and (_12760_, _12759_, _06555_);
  not (_12761_, _06555_);
  and (_12762_, _12627_, _12761_);
  or (_12763_, _12762_, _04891_);
  or (_12764_, _12763_, _12760_);
  or (_12765_, _12627_, _06548_);
  and (_12766_, _12765_, _04728_);
  and (_12767_, _12766_, _12764_);
  or (_12768_, _12767_, _12614_);
  and (_12769_, _12768_, _06562_);
  or (_12770_, _12769_, _12611_);
  and (_12771_, _12770_, _06956_);
  and (_12772_, _10243_, _03833_);
  or (_12773_, _12772_, _03400_);
  or (_12774_, _12773_, _12771_);
  and (_12775_, _03879_, _03400_);
  nor (_12776_, _12775_, _03672_);
  and (_12777_, _12776_, _12774_);
  and (_12778_, _12622_, _03672_);
  or (_12779_, _12778_, _12587_);
  or (_12780_, _12779_, _12777_);
  nor (_12781_, _08218_, _08216_);
  nor (_12782_, _12781_, _06917_);
  or (_12783_, _12782_, _10909_);
  and (_12784_, _12783_, _04744_);
  and (_12785_, _12784_, _12780_);
  or (_12786_, _08038_, _06937_);
  nor (_12787_, _06940_, _04744_);
  and (_12788_, _12787_, _12786_);
  or (_12789_, _12788_, _04742_);
  or (_12790_, _12789_, _12785_);
  nor (_12791_, _05701_, _05554_);
  nor (_12792_, _12791_, _05702_);
  or (_12793_, _12792_, _04922_);
  and (_12794_, _12793_, _04993_);
  and (_12795_, _12794_, _12790_);
  and (_12796_, _12795_, _11999_);
  or (_12797_, _12796_, _12608_);
  nand (_12798_, _10205_, _03833_);
  or (_12799_, _10055_, _03833_);
  and (_12800_, _12799_, _12798_);
  or (_12801_, _12800_, _12008_);
  and (_40490_, _12801_, _12797_);
  or (_12802_, _12000_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_12803_, _12802_, _12008_);
  nor (_12804_, _06940_, _06942_);
  nor (_12805_, _12804_, _08022_);
  or (_12806_, _12805_, _04744_);
  nand (_12807_, _10085_, _03483_);
  nor (_12808_, _10748_, _10747_);
  and (_12809_, _10748_, \oc8051_golden_model_1.PSW [7]);
  nor (_12810_, _12809_, _12808_);
  nor (_12811_, _12810_, _05114_);
  or (_12812_, _12808_, _06123_);
  and (_12813_, _10084_, _04111_);
  nor (_12814_, _04111_, _07640_);
  or (_12815_, _12814_, _12813_);
  and (_12816_, _12815_, _06140_);
  nor (_12817_, _06133_, _05898_);
  and (_12818_, _06133_, _05898_);
  or (_12819_, _12818_, _12817_);
  and (_12820_, _12819_, _10320_);
  or (_12821_, _12820_, _12816_);
  and (_12822_, _12821_, _04625_);
  and (_12823_, _06942_, _04624_);
  or (_12824_, _12823_, _12822_);
  and (_12825_, _12824_, _04816_);
  nor (_12826_, _06245_, _05900_);
  and (_12827_, _06245_, _05900_);
  nor (_12828_, _12827_, _12826_);
  nor (_12829_, _12828_, _04816_);
  or (_12830_, _12829_, _12825_);
  and (_12831_, _12830_, _06125_);
  nand (_12832_, _10749_, _10747_);
  and (_12833_, _12832_, _04629_);
  or (_12834_, _12833_, _04933_);
  or (_12835_, _12834_, _12831_);
  nor (_12836_, _10084_, _03445_);
  nor (_12837_, _12836_, _04640_);
  and (_12838_, _12837_, _12835_);
  and (_12839_, _08199_, _04640_);
  or (_12840_, _12839_, _03694_);
  or (_12841_, _12840_, _12838_);
  and (_12842_, _12841_, _12812_);
  or (_12843_, _12842_, _03690_);
  nand (_12844_, _05900_, _03690_);
  and (_12845_, _12844_, _03688_);
  and (_12846_, _12845_, _12843_);
  not (_12847_, _10750_);
  and (_12848_, _12832_, _12847_);
  and (_12849_, _12848_, _03687_);
  or (_12850_, _12849_, _12846_);
  and (_12851_, _12850_, _03442_);
  or (_12852_, _10085_, _03442_);
  nand (_12853_, _12852_, _03807_);
  or (_12854_, _12853_, _12851_);
  nand (_12855_, _05900_, _03808_);
  and (_12856_, _12855_, _12854_);
  or (_12857_, _12856_, _04269_);
  and (_12858_, _06942_, _05351_);
  nand (_12859_, _05845_, _04269_);
  or (_12860_, _12859_, _12858_);
  and (_12861_, _12860_, _05114_);
  and (_12862_, _12861_, _12857_);
  or (_12863_, _12862_, _12811_);
  and (_12864_, _12863_, _03418_);
  or (_12865_, _10085_, _03418_);
  nand (_12866_, _12865_, _04677_);
  or (_12867_, _12866_, _12864_);
  nand (_12868_, _05898_, _06291_);
  and (_12869_, _12868_, _12867_);
  or (_12870_, _12869_, _04680_);
  or (_12871_, _06942_, _06297_);
  and (_12872_, _12871_, _06296_);
  and (_12873_, _12872_, _12870_);
  nor (_12874_, _06307_, _05898_);
  and (_12875_, _06438_, \oc8051_golden_model_1.SP [4]);
  and (_12876_, _06443_, \oc8051_golden_model_1.TL0 [4]);
  nor (_12877_, _12876_, _12875_);
  and (_12878_, _06463_, \oc8051_golden_model_1.DPL [4]);
  and (_12879_, _06493_, \oc8051_golden_model_1.TMOD [4]);
  nor (_12880_, _12879_, _12878_);
  and (_12881_, _12880_, _12877_);
  and (_12882_, _06482_, \oc8051_golden_model_1.IE [4]);
  and (_12883_, _06485_, \oc8051_golden_model_1.SBUF [4]);
  and (_12884_, _06487_, \oc8051_golden_model_1.SCON [4]);
  or (_12885_, _12884_, _12883_);
  nor (_12886_, _12885_, _12882_);
  and (_12887_, _06470_, \oc8051_golden_model_1.P1INREG [4]);
  not (_12888_, _12887_);
  and (_12889_, _06466_, \oc8051_golden_model_1.P0INREG [4]);
  not (_12890_, _12889_);
  and (_12891_, _06474_, \oc8051_golden_model_1.P2INREG [4]);
  and (_12892_, _06476_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_12893_, _12892_, _12891_);
  and (_12894_, _12893_, _12890_);
  and (_12895_, _12894_, _12888_);
  and (_12896_, _12895_, _12886_);
  and (_12897_, _12896_, _12881_);
  and (_12898_, _06420_, \oc8051_golden_model_1.IP [4]);
  and (_12899_, _06409_, \oc8051_golden_model_1.ACC [4]);
  nor (_12900_, _12899_, _12898_);
  and (_12901_, _06424_, \oc8051_golden_model_1.PSW [4]);
  and (_12902_, _06412_, \oc8051_golden_model_1.B [4]);
  nor (_12903_, _12902_, _12901_);
  and (_12904_, _12903_, _12900_);
  and (_12905_, _06491_, \oc8051_golden_model_1.DPH [4]);
  and (_12906_, _06434_, \oc8051_golden_model_1.TH1 [4]);
  nor (_12907_, _12906_, _12905_);
  and (_12908_, _12907_, _12904_);
  and (_12909_, _06455_, \oc8051_golden_model_1.TCON [4]);
  and (_12910_, _06448_, \oc8051_golden_model_1.TH0 [4]);
  nor (_12911_, _12910_, _12909_);
  and (_12912_, _06459_, \oc8051_golden_model_1.PCON [4]);
  and (_12913_, _06452_, \oc8051_golden_model_1.TL1 [4]);
  nor (_12914_, _12913_, _12912_);
  and (_12915_, _12914_, _12911_);
  and (_12916_, _12915_, _12908_);
  and (_12917_, _12916_, _12897_);
  not (_12918_, _12917_);
  nor (_12919_, _12918_, _12874_);
  nor (_12920_, _12919_, _06296_);
  or (_12921_, _12920_, _06306_);
  or (_12922_, _12921_, _12873_);
  and (_12923_, _06306_, _04446_);
  nor (_12924_, _12923_, _04695_);
  and (_12925_, _12924_, _12922_);
  and (_12926_, _06422_, _04695_);
  or (_12927_, _12926_, _03483_);
  or (_12928_, _12927_, _12925_);
  and (_12929_, _12928_, _12807_);
  or (_12930_, _12929_, _04704_);
  and (_12931_, _06339_, _05900_);
  nor (_12932_, _06339_, _05900_);
  nor (_12933_, _12932_, _12931_);
  and (_12934_, _12933_, _06520_);
  or (_12935_, _12934_, _04705_);
  and (_12936_, _12935_, _12930_);
  and (_12937_, _08700_, _04702_);
  or (_12938_, _12937_, _04709_);
  or (_12939_, _12938_, _12936_);
  or (_12940_, _12932_, _06519_);
  and (_12941_, _12940_, _06030_);
  and (_12942_, _12941_, _12939_);
  and (_12943_, _08698_, _04707_);
  or (_12944_, _12943_, _03477_);
  or (_12945_, _12944_, _12942_);
  and (_12946_, _10085_, _03477_);
  nor (_12947_, _12946_, _06533_);
  and (_12948_, _12947_, _12945_);
  nor (_12949_, _12931_, _06539_);
  or (_12950_, _12949_, _06538_);
  or (_12951_, _12950_, _12948_);
  nand (_12952_, _08699_, _06538_);
  and (_12953_, _12952_, _06543_);
  and (_12954_, _12953_, _12951_);
  nand (_12955_, _10084_, _03474_);
  nand (_12956_, _12955_, _06556_);
  or (_12957_, _12956_, _12954_);
  or (_12958_, _12819_, _06556_);
  and (_12959_, _12958_, _12355_);
  and (_12960_, _12959_, _12957_);
  and (_12961_, _06791_, _06881_);
  nor (_12962_, _06791_, _06881_);
  nor (_12963_, _12962_, _12961_);
  nand (_12964_, _12963_, _04083_);
  and (_12965_, _12964_, _04727_);
  or (_12966_, _12965_, _12960_);
  nand (_12967_, _12963_, _12202_);
  and (_12968_, _12967_, _06562_);
  and (_12969_, _12968_, _12966_);
  nor (_12970_, _12828_, _06562_);
  or (_12971_, _12970_, _03833_);
  or (_12972_, _12971_, _12969_);
  nand (_12973_, _10240_, _03833_);
  and (_12974_, _12973_, _10904_);
  and (_12975_, _12974_, _12972_);
  and (_12976_, _10084_, _03400_);
  or (_12977_, _12976_, _03672_);
  or (_12978_, _12977_, _12975_);
  or (_12979_, _12808_, _03673_);
  and (_12980_, _12979_, _10909_);
  and (_12981_, _12980_, _12978_);
  nor (_12982_, _06917_, _08199_);
  nor (_12983_, _12982_, _08200_);
  and (_12984_, _12983_, _12587_);
  or (_12985_, _12984_, _04743_);
  or (_12986_, _12985_, _12981_);
  and (_12987_, _12986_, _12806_);
  or (_12988_, _12987_, _04742_);
  and (_12989_, _08303_, _05702_);
  nor (_12990_, _08303_, _05702_);
  nor (_12991_, _12990_, _12989_);
  or (_12992_, _12991_, _04922_);
  and (_12993_, _12992_, _04993_);
  and (_12994_, _12993_, _12988_);
  or (_12995_, _12994_, _12010_);
  and (_12996_, _12995_, _12803_);
  nand (_12997_, _10201_, _03833_);
  or (_12998_, _10048_, _03833_);
  and (_12999_, _12998_, _12997_);
  and (_13000_, _12999_, _05334_);
  and (_13001_, _13000_, _12187_);
  or (_40491_, _13001_, _12996_);
  or (_13002_, _12000_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_13003_, _13002_, _12008_);
  nor (_13004_, _12961_, _06836_);
  or (_13005_, _13004_, _06883_);
  and (_13006_, _13005_, _12202_);
  nor (_13007_, _10855_, _10854_);
  and (_13008_, _10855_, \oc8051_golden_model_1.PSW [7]);
  nor (_13009_, _13008_, _13007_);
  nor (_13010_, _13009_, _05114_);
  or (_13011_, _13007_, _06123_);
  nor (_13012_, _12818_, _05799_);
  or (_13013_, _13012_, _06134_);
  and (_13014_, _13013_, _10320_);
  nor (_13015_, _04111_, _07634_);
  and (_13016_, _10079_, _04111_);
  or (_13017_, _13016_, _13015_);
  and (_13018_, _13017_, _06140_);
  or (_13019_, _13018_, _13014_);
  and (_13020_, _13019_, _04625_);
  and (_13021_, _06941_, _04624_);
  or (_13022_, _13021_, _13020_);
  and (_13023_, _13022_, _04816_);
  nor (_13024_, _12827_, _05801_);
  nor (_13025_, _13024_, _06246_);
  nor (_13026_, _13025_, _04816_);
  or (_13027_, _13026_, _13023_);
  and (_13028_, _13027_, _06125_);
  nand (_13029_, _10856_, _10854_);
  and (_13030_, _13029_, _04629_);
  or (_13031_, _13030_, _04933_);
  or (_13032_, _13031_, _13028_);
  nor (_13033_, _10079_, _03445_);
  nor (_13034_, _13033_, _04640_);
  and (_13035_, _13034_, _13032_);
  and (_13036_, _08198_, _04640_);
  or (_13037_, _13036_, _03694_);
  or (_13038_, _13037_, _13035_);
  and (_13039_, _13038_, _13011_);
  or (_13040_, _13039_, _03690_);
  nand (_13041_, _05801_, _03690_);
  and (_13042_, _13041_, _03688_);
  and (_13043_, _13042_, _13040_);
  not (_13044_, _10857_);
  and (_13045_, _13029_, _13044_);
  and (_13046_, _13045_, _03687_);
  or (_13047_, _13046_, _13043_);
  and (_13048_, _13047_, _03442_);
  or (_13049_, _10080_, _03442_);
  nand (_13050_, _13049_, _03807_);
  or (_13051_, _13050_, _13048_);
  nand (_13052_, _05801_, _03808_);
  and (_13053_, _13052_, _13051_);
  or (_13054_, _13053_, _04269_);
  and (_13055_, _06941_, _05351_);
  nand (_13056_, _05746_, _04269_);
  or (_13057_, _13056_, _13055_);
  and (_13058_, _13057_, _05114_);
  and (_13059_, _13058_, _13054_);
  or (_13060_, _13059_, _13010_);
  and (_13061_, _13060_, _03418_);
  or (_13062_, _10080_, _03418_);
  nand (_13063_, _13062_, _04677_);
  or (_13064_, _13063_, _13061_);
  nand (_13065_, _05799_, _06291_);
  and (_13066_, _13065_, _13064_);
  or (_13067_, _13066_, _04680_);
  or (_13068_, _06941_, _12070_);
  and (_13069_, _13068_, _12069_);
  and (_13070_, _13069_, _13067_);
  nor (_13071_, _06307_, _05799_);
  and (_13072_, _06420_, \oc8051_golden_model_1.IP [5]);
  and (_13073_, _06412_, \oc8051_golden_model_1.B [5]);
  nor (_13074_, _13073_, _13072_);
  and (_13075_, _06424_, \oc8051_golden_model_1.PSW [5]);
  and (_13076_, _06409_, \oc8051_golden_model_1.ACC [5]);
  nor (_13077_, _13076_, _13075_);
  and (_13078_, _13077_, _13074_);
  and (_13079_, _06485_, \oc8051_golden_model_1.SBUF [5]);
  not (_13080_, _13079_);
  and (_13081_, _06487_, \oc8051_golden_model_1.SCON [5]);
  and (_13082_, _06482_, \oc8051_golden_model_1.IE [5]);
  nor (_13083_, _13082_, _13081_);
  and (_13084_, _13083_, _13080_);
  and (_13085_, _06466_, \oc8051_golden_model_1.P0INREG [5]);
  not (_13086_, _13085_);
  and (_13087_, _06476_, \oc8051_golden_model_1.P3INREG [5]);
  and (_13088_, _06470_, \oc8051_golden_model_1.P1INREG [5]);
  and (_13089_, _06474_, \oc8051_golden_model_1.P2INREG [5]);
  or (_13090_, _13089_, _13088_);
  nor (_13091_, _13090_, _13087_);
  and (_13092_, _13091_, _13086_);
  and (_13093_, _13092_, _13084_);
  and (_13094_, _13093_, _13078_);
  and (_13095_, _06448_, \oc8051_golden_model_1.TH0 [5]);
  and (_13096_, _06452_, \oc8051_golden_model_1.TL1 [5]);
  nor (_13097_, _13096_, _13095_);
  and (_13098_, _06455_, \oc8051_golden_model_1.TCON [5]);
  and (_13099_, _06459_, \oc8051_golden_model_1.PCON [5]);
  nor (_13100_, _13099_, _13098_);
  and (_13101_, _13100_, _13097_);
  and (_13102_, _06491_, \oc8051_golden_model_1.DPH [5]);
  not (_13103_, _13102_);
  and (_13104_, _06434_, \oc8051_golden_model_1.TH1 [5]);
  and (_13105_, _06443_, \oc8051_golden_model_1.TL0 [5]);
  nor (_13106_, _13105_, _13104_);
  and (_13107_, _13106_, _13103_);
  and (_13108_, _06438_, \oc8051_golden_model_1.SP [5]);
  not (_13109_, _13108_);
  and (_13110_, _06463_, \oc8051_golden_model_1.DPL [5]);
  and (_13111_, _06493_, \oc8051_golden_model_1.TMOD [5]);
  nor (_13112_, _13111_, _13110_);
  and (_13113_, _13112_, _13109_);
  and (_13114_, _13113_, _13107_);
  and (_13115_, _13114_, _13101_);
  and (_13116_, _13115_, _13094_);
  not (_13117_, _13116_);
  nor (_13118_, _13117_, _13071_);
  nor (_13119_, _13118_, _06296_);
  or (_13120_, _13119_, _06306_);
  or (_13121_, _13120_, _13070_);
  and (_13122_, _06306_, _04034_);
  nor (_13123_, _13122_, _04695_);
  and (_13124_, _13123_, _13121_);
  and (_13125_, _06371_, _04695_);
  or (_13126_, _13125_, _03483_);
  or (_13127_, _13126_, _13124_);
  and (_13128_, _10080_, _03483_);
  nor (_13129_, _13128_, _04704_);
  and (_13130_, _13129_, _13127_);
  and (_13131_, _06370_, _05801_);
  nor (_13132_, _06370_, _05801_);
  nor (_13133_, _13132_, _13131_);
  nor (_13134_, _13133_, _04702_);
  nor (_13135_, _13134_, _04705_);
  or (_13136_, _13135_, _13130_);
  or (_13137_, _10451_, _06520_);
  and (_13138_, _13137_, _06519_);
  and (_13139_, _13138_, _13136_);
  and (_13140_, _13132_, _04709_);
  or (_13141_, _13140_, _13139_);
  and (_13142_, _13141_, _06030_);
  and (_13143_, _08696_, _04707_);
  or (_13144_, _13143_, _03477_);
  or (_13145_, _13144_, _13142_);
  and (_13146_, _10080_, _03477_);
  nor (_13147_, _13146_, _06533_);
  and (_13148_, _13147_, _13145_);
  nor (_13149_, _13131_, _06539_);
  or (_13150_, _13149_, _06538_);
  or (_13151_, _13150_, _13148_);
  nand (_13152_, _08697_, _06538_);
  and (_13153_, _13152_, _06543_);
  and (_13154_, _13153_, _13151_);
  and (_13155_, _03786_, _03254_);
  nor (_13156_, _12761_, _13155_);
  and (_13157_, _03789_, _03254_);
  and (_13158_, _10079_, _03474_);
  nor (_13159_, _13158_, _13157_);
  nand (_13160_, _13159_, _13156_);
  or (_13161_, _13160_, _13154_);
  or (_13162_, _13013_, _06556_);
  and (_13163_, _13162_, _12355_);
  and (_13164_, _13163_, _13161_);
  and (_13165_, _13005_, _12354_);
  or (_13166_, _13165_, _13164_);
  and (_13167_, _13166_, _12203_);
  or (_13168_, _13167_, _13006_);
  and (_13169_, _13168_, _06562_);
  nor (_13170_, _13025_, _06562_);
  or (_13171_, _13170_, _03833_);
  or (_13172_, _13171_, _13169_);
  nand (_13173_, _10235_, _03833_);
  and (_13174_, _13173_, _10904_);
  and (_13175_, _13174_, _13172_);
  and (_13176_, _10079_, _03400_);
  or (_13177_, _13176_, _03672_);
  or (_13178_, _13177_, _13175_);
  or (_13179_, _13007_, _03673_);
  and (_13180_, _13179_, _10909_);
  and (_13181_, _13180_, _13178_);
  or (_13182_, _08200_, _08198_);
  nor (_13183_, _10909_, _06919_);
  and (_13184_, _13183_, _13182_);
  or (_13185_, _13184_, _13181_);
  and (_13186_, _13185_, _04744_);
  or (_13187_, _08022_, _06941_);
  nor (_13188_, _06944_, _04744_);
  and (_13189_, _13188_, _13187_);
  or (_13190_, _13189_, _04742_);
  or (_13191_, _13190_, _13186_);
  nor (_13192_, _12989_, _08302_);
  nor (_13193_, _13192_, _05902_);
  or (_13194_, _13193_, _04922_);
  and (_13195_, _13194_, _04993_);
  and (_13196_, _13195_, _13191_);
  or (_13197_, _13196_, _12010_);
  and (_13198_, _13197_, _13003_);
  or (_13199_, _10195_, _06956_);
  or (_13200_, _10044_, _03833_);
  and (_13201_, _13200_, _13199_);
  and (_13202_, _13201_, _05334_);
  and (_13203_, _13202_, _12187_);
  or (_40493_, _13203_, _13198_);
  or (_13204_, _12000_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_13205_, _13204_, _12008_);
  nor (_13206_, _06944_, _06933_);
  nor (_13207_, _13206_, _06945_);
  and (_13208_, _13207_, _12384_);
  nor (_13209_, _06919_, _06013_);
  and (_13210_, _06919_, _06013_);
  or (_13211_, _13210_, _13209_);
  and (_13212_, _13211_, _12587_);
  nor (_13213_, _06134_, _06013_);
  nor (_13214_, _13213_, _06135_);
  nand (_13215_, _13214_, _12761_);
  nor (_13216_, _06406_, _06015_);
  and (_13217_, _13216_, _04709_);
  nor (_13218_, _10803_, _10802_);
  and (_13219_, _10803_, \oc8051_golden_model_1.PSW [7]);
  nor (_13220_, _13219_, _13218_);
  nor (_13221_, _13220_, _05114_);
  or (_13222_, _13218_, _06123_);
  nand (_13223_, _13214_, _10320_);
  nor (_13224_, _04111_, _07586_);
  and (_13225_, _10071_, _04111_);
  or (_13226_, _13225_, _13224_);
  or (_13227_, _13226_, _10320_);
  and (_13228_, _13227_, _13223_);
  or (_13229_, _13228_, _04624_);
  or (_13230_, _06933_, _04625_);
  and (_13231_, _13230_, _13229_);
  and (_13232_, _13231_, _04816_);
  nor (_13233_, _06246_, _06015_);
  nor (_13234_, _13233_, _06247_);
  nor (_13235_, _13234_, _04816_);
  or (_13236_, _13235_, _13232_);
  and (_13237_, _13236_, _06125_);
  nand (_13238_, _10804_, _10802_);
  and (_13239_, _13238_, _04629_);
  or (_13240_, _13239_, _04933_);
  or (_13241_, _13240_, _13237_);
  nor (_13242_, _10071_, _03445_);
  nor (_13243_, _13242_, _04640_);
  and (_13244_, _13243_, _13241_);
  and (_13245_, _08185_, _04640_);
  or (_13246_, _13245_, _03694_);
  or (_13247_, _13246_, _13244_);
  and (_13248_, _13247_, _13222_);
  or (_13249_, _13248_, _03690_);
  nand (_13250_, _06015_, _03690_);
  and (_13251_, _13250_, _03688_);
  and (_13252_, _13251_, _13249_);
  not (_13253_, _10805_);
  and (_13254_, _13238_, _13253_);
  and (_13255_, _13254_, _03687_);
  or (_13256_, _13255_, _13252_);
  and (_13257_, _13256_, _03442_);
  or (_13258_, _10072_, _03442_);
  nand (_13259_, _13258_, _03807_);
  or (_13260_, _13259_, _13257_);
  nand (_13261_, _06015_, _03808_);
  and (_13262_, _13261_, _13260_);
  or (_13263_, _13262_, _04269_);
  and (_13264_, _06933_, _05351_);
  nand (_13265_, _05947_, _04269_);
  or (_13266_, _13265_, _13264_);
  and (_13267_, _13266_, _05114_);
  and (_13268_, _13267_, _13263_);
  or (_13269_, _13268_, _13221_);
  and (_13270_, _13269_, _03418_);
  or (_13271_, _10072_, _03418_);
  nand (_13272_, _13271_, _04677_);
  or (_13273_, _13272_, _13270_);
  nand (_13274_, _06013_, _06291_);
  and (_13275_, _13274_, _13273_);
  or (_13276_, _13275_, _04680_);
  or (_13277_, _06933_, _12070_);
  and (_13278_, _13277_, _12069_);
  and (_13279_, _13278_, _13276_);
  nor (_13280_, _06307_, _06013_);
  and (_13281_, _06412_, \oc8051_golden_model_1.B [6]);
  and (_13282_, _06409_, \oc8051_golden_model_1.ACC [6]);
  nor (_13283_, _13282_, _13281_);
  and (_13284_, _06420_, \oc8051_golden_model_1.IP [6]);
  and (_13285_, _06424_, \oc8051_golden_model_1.PSW [6]);
  nor (_13286_, _13285_, _13284_);
  and (_13287_, _13286_, _13283_);
  and (_13288_, _06493_, \oc8051_golden_model_1.TMOD [6]);
  and (_13289_, _06491_, \oc8051_golden_model_1.DPH [6]);
  nor (_13290_, _13289_, _13288_);
  and (_13291_, _06443_, \oc8051_golden_model_1.TL0 [6]);
  and (_13292_, _06434_, \oc8051_golden_model_1.TH1 [6]);
  nor (_13293_, _13292_, _13291_);
  and (_13294_, _13293_, _13290_);
  and (_13295_, _13294_, _13287_);
  and (_13296_, _06476_, \oc8051_golden_model_1.P3INREG [6]);
  not (_13297_, _13296_);
  and (_13298_, _06470_, \oc8051_golden_model_1.P1INREG [6]);
  and (_13299_, _06474_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_13300_, _13299_, _13298_);
  and (_13301_, _13300_, _13297_);
  and (_13302_, _06482_, \oc8051_golden_model_1.IE [6]);
  not (_13303_, _13302_);
  and (_13304_, _06487_, \oc8051_golden_model_1.SCON [6]);
  and (_13305_, _06485_, \oc8051_golden_model_1.SBUF [6]);
  nor (_13306_, _13305_, _13304_);
  and (_13307_, _13306_, _13303_);
  and (_13308_, _13307_, _13301_);
  and (_13309_, _06448_, \oc8051_golden_model_1.TH0 [6]);
  and (_13310_, _06452_, \oc8051_golden_model_1.TL1 [6]);
  nor (_13311_, _13310_, _13309_);
  and (_13312_, _06455_, \oc8051_golden_model_1.TCON [6]);
  and (_13313_, _06459_, \oc8051_golden_model_1.PCON [6]);
  nor (_13314_, _13313_, _13312_);
  and (_13315_, _13314_, _13311_);
  and (_13316_, _06463_, \oc8051_golden_model_1.DPL [6]);
  not (_13317_, _13316_);
  and (_13318_, _06438_, \oc8051_golden_model_1.SP [6]);
  and (_13319_, _06466_, \oc8051_golden_model_1.P0INREG [6]);
  nor (_13320_, _13319_, _13318_);
  and (_13321_, _13320_, _13317_);
  and (_13322_, _13321_, _13315_);
  and (_13323_, _13322_, _13308_);
  and (_13324_, _13323_, _13295_);
  not (_13325_, _13324_);
  nor (_13326_, _13325_, _13280_);
  nor (_13327_, _13326_, _06296_);
  or (_13328_, _13327_, _06306_);
  or (_13329_, _13328_, _13279_);
  and (_13330_, _06306_, _03740_);
  nor (_13331_, _13330_, _04695_);
  and (_13332_, _13331_, _13329_);
  not (_13333_, _06406_);
  and (_13334_, _13333_, _04695_);
  or (_13335_, _13334_, _03483_);
  or (_13336_, _13335_, _13332_);
  and (_13337_, _10072_, _03483_);
  nor (_13338_, _13337_, _04704_);
  and (_13339_, _13338_, _13336_);
  and (_13340_, _06406_, _06015_);
  nor (_13341_, _13340_, _13216_);
  nor (_13342_, _13341_, _04702_);
  nor (_13343_, _13342_, _04705_);
  or (_13344_, _13343_, _13339_);
  or (_13345_, _08695_, _06520_);
  and (_13346_, _13345_, _06519_);
  and (_13347_, _13346_, _13344_);
  or (_13348_, _13347_, _13217_);
  and (_13349_, _13348_, _06030_);
  and (_13350_, _08693_, _04707_);
  or (_13351_, _13350_, _03477_);
  or (_13352_, _13351_, _13349_);
  and (_13353_, _10072_, _03477_);
  nor (_13354_, _13353_, _06533_);
  and (_13355_, _13354_, _13352_);
  nor (_13356_, _13340_, _06539_);
  or (_13357_, _13356_, _06538_);
  or (_13358_, _13357_, _13355_);
  nand (_13359_, _08694_, _06538_);
  and (_13360_, _13359_, _06543_);
  and (_13361_, _13360_, _13358_);
  nand (_13362_, _10071_, _03474_);
  nand (_13363_, _13362_, _06555_);
  or (_13364_, _13363_, _13361_);
  nand (_13365_, _13364_, _13215_);
  and (_13366_, _13365_, _06548_);
  and (_13367_, _13214_, _04891_);
  or (_13368_, _13367_, _12354_);
  nor (_13369_, _13368_, _13366_);
  nor (_13370_, _06883_, _06607_);
  nor (_13371_, _13370_, _06884_);
  nand (_13372_, _13371_, _04083_);
  and (_13373_, _13372_, _04727_);
  or (_13374_, _13373_, _13369_);
  nand (_13375_, _13371_, _12202_);
  and (_13376_, _13375_, _06562_);
  and (_13377_, _13376_, _13374_);
  nor (_13378_, _13234_, _06562_);
  or (_13379_, _13378_, _03833_);
  or (_13380_, _13379_, _13377_);
  nand (_13381_, _10227_, _03833_);
  and (_13382_, _13381_, _10904_);
  and (_13383_, _13382_, _13380_);
  and (_13384_, _10071_, _03400_);
  or (_13385_, _13384_, _03672_);
  or (_13386_, _13385_, _13383_);
  or (_13387_, _13218_, _03673_);
  and (_13388_, _13387_, _10909_);
  and (_13389_, _13388_, _13386_);
  or (_13390_, _13389_, _13212_);
  and (_13391_, _13390_, _12385_);
  or (_13392_, _13391_, _13208_);
  and (_13393_, _13392_, _12196_);
  and (_13394_, _13207_, _12195_);
  or (_13395_, _13394_, _04742_);
  or (_13396_, _13395_, _13393_);
  nor (_13397_, _06015_, _05902_);
  and (_13398_, _06015_, _05902_);
  nor (_13399_, _13398_, _13397_);
  nand (_13400_, _13399_, _04742_);
  and (_13401_, _13400_, _04993_);
  and (_13402_, _13401_, _13396_);
  or (_13403_, _13402_, _12010_);
  and (_13404_, _13403_, _13205_);
  or (_13405_, _10188_, _06956_);
  or (_13406_, _10038_, _03833_);
  and (_13407_, _13406_, _13405_);
  and (_13408_, _13407_, _05334_);
  and (_13409_, _13408_, _12187_);
  or (_40494_, _13409_, _13404_);
  or (_13410_, _12000_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_13411_, _13410_, _12008_);
  nand (_13412_, _12000_, _06952_);
  and (_13413_, _13412_, _13411_);
  and (_13414_, _12187_, _06980_);
  or (_40495_, _13414_, _13413_);
  nor (_13415_, _05331_, _04992_);
  not (_13416_, _13415_);
  nor (_13417_, _13416_, _05173_);
  nor (_13418_, _13416_, _05318_);
  nor (_13419_, _13418_, _13417_);
  nor (_13420_, _13416_, _04749_);
  and (_13421_, _13420_, _04914_);
  and (_13422_, _13421_, _13419_);
  or (_13423_, _13422_, \oc8051_golden_model_1.IRAM[1] [0]);
  not (_13424_, _12002_);
  nand (_13425_, _12005_, _05055_);
  or (_13426_, _13425_, _13424_);
  and (_13427_, _13426_, _13423_);
  and (_13428_, _12179_, _13415_);
  and (_13429_, _13428_, _12178_);
  not (_13430_, _13422_);
  or (_13431_, _13430_, _13429_);
  and (_13432_, _13431_, _13427_);
  and (_13433_, _05334_, _05055_);
  and (_13434_, _13433_, _12185_);
  and (_13435_, _13434_, _12191_);
  or (_40500_, _13435_, _13432_);
  or (_13436_, _13422_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_13437_, _13436_, _13426_);
  and (_13438_, _12395_, _13415_);
  and (_13439_, _13438_, _12394_);
  or (_13440_, _13430_, _13439_);
  and (_13441_, _13440_, _13437_);
  and (_13442_, _13434_, _12403_);
  or (_40501_, _13442_, _13441_);
  or (_13443_, _13422_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_13444_, _13443_, _13426_);
  and (_13445_, _12597_, _13415_);
  and (_13446_, _13445_, _12594_);
  or (_13447_, _13430_, _13446_);
  and (_13448_, _13447_, _13444_);
  and (_13449_, _13434_, _12605_);
  or (_40502_, _13449_, _13448_);
  or (_13450_, _13422_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_13451_, _13450_, _13426_);
  and (_13452_, _12793_, _13415_);
  and (_13453_, _13452_, _12790_);
  or (_13454_, _13430_, _13453_);
  and (_13455_, _13454_, _13451_);
  and (_13456_, _12800_, _05334_);
  and (_13457_, _13434_, _13456_);
  or (_40503_, _13457_, _13455_);
  or (_13458_, _13422_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_13459_, _13458_, _13426_);
  and (_13460_, _12992_, _13415_);
  and (_13461_, _13460_, _12988_);
  or (_13462_, _13430_, _13461_);
  and (_13463_, _13462_, _13459_);
  and (_13464_, _13434_, _13000_);
  or (_40505_, _13464_, _13463_);
  or (_13465_, _13422_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_13466_, _13465_, _13426_);
  and (_13467_, _13194_, _13415_);
  and (_13468_, _13467_, _13191_);
  or (_13469_, _13430_, _13468_);
  and (_13470_, _13469_, _13466_);
  and (_13471_, _13434_, _13202_);
  or (_40506_, _13471_, _13470_);
  or (_13472_, _13422_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_13473_, _13472_, _13426_);
  and (_13474_, _13400_, _13415_);
  and (_13475_, _13474_, _13396_);
  or (_13476_, _13430_, _13475_);
  and (_13477_, _13476_, _13473_);
  and (_13478_, _13434_, _13408_);
  or (_40507_, _13478_, _13477_);
  or (_13479_, _13422_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_13480_, _13479_, _13426_);
  nor (_13481_, _06952_, _13416_);
  or (_13482_, _13430_, _13481_);
  and (_13483_, _13482_, _13480_);
  and (_13484_, _13434_, _06980_);
  or (_40508_, _13484_, _13483_);
  and (_13485_, _04995_, _04749_);
  and (_13486_, _13485_, _11998_);
  or (_13487_, _13486_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_13488_, _12005_, _06151_);
  or (_13489_, _13488_, _13424_);
  and (_13490_, _13489_, _13487_);
  not (_13491_, _13486_);
  or (_13492_, _13491_, _12181_);
  and (_13493_, _13492_, _13490_);
  and (_13494_, _06151_, _05334_);
  and (_13495_, _13494_, _12185_);
  and (_13496_, _13495_, _12191_);
  or (_40512_, _13496_, _13493_);
  or (_13497_, _13486_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_13498_, _13497_, _13489_);
  or (_13499_, _13491_, _12397_);
  and (_13500_, _13499_, _13498_);
  and (_13501_, _13495_, _12403_);
  or (_40514_, _13501_, _13500_);
  or (_13502_, _13486_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_13503_, _13502_, _13489_);
  or (_13504_, _13491_, _12599_);
  and (_13505_, _13504_, _13503_);
  and (_13506_, _13495_, _12605_);
  or (_40515_, _13506_, _13505_);
  or (_13507_, _13486_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_13508_, _13507_, _13489_);
  or (_13509_, _13491_, _12795_);
  and (_13510_, _13509_, _13508_);
  and (_13511_, _13495_, _13456_);
  or (_40516_, _13511_, _13510_);
  or (_13512_, _13486_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_13513_, _13512_, _13489_);
  or (_13514_, _13491_, _12994_);
  and (_13515_, _13514_, _13513_);
  and (_13516_, _13495_, _13000_);
  or (_40517_, _13516_, _13515_);
  or (_13517_, _13491_, _13196_);
  or (_13518_, _13486_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_13519_, _13518_, _13489_);
  and (_13520_, _13519_, _13517_);
  and (_13521_, _13495_, _13202_);
  or (_40518_, _13521_, _13520_);
  or (_13522_, _13486_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_13523_, _13522_, _13489_);
  or (_13524_, _13491_, _13402_);
  and (_13525_, _13524_, _13523_);
  and (_13526_, _13495_, _13408_);
  or (_40520_, _13526_, _13525_);
  or (_13527_, _13486_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_13528_, _13527_, _13489_);
  or (_13529_, _13491_, _06953_);
  and (_13530_, _13529_, _13528_);
  and (_13531_, _13495_, _06980_);
  or (_40521_, _13531_, _13530_);
  and (_13532_, _11998_, _04997_);
  or (_13533_, _13532_, \oc8051_golden_model_1.IRAM[3] [0]);
  nand (_13534_, _12005_, _04752_);
  or (_13535_, _13534_, _13424_);
  and (_13536_, _13535_, _13533_);
  not (_13537_, _13532_);
  or (_13538_, _13537_, _12181_);
  and (_13539_, _13538_, _13536_);
  and (_13540_, _05334_, _04752_);
  and (_13541_, _13540_, _12185_);
  and (_13542_, _13541_, _12191_);
  or (_40525_, _13542_, _13539_);
  or (_13543_, _13532_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_13544_, _13543_, _13535_);
  or (_13545_, _13537_, _12397_);
  and (_13546_, _13545_, _13544_);
  and (_13547_, _13541_, _12403_);
  or (_40526_, _13547_, _13546_);
  or (_13548_, _13532_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_13549_, _13548_, _13535_);
  or (_13550_, _13537_, _12599_);
  and (_13551_, _13550_, _13549_);
  and (_13552_, _13541_, _12605_);
  or (_40527_, _13552_, _13551_);
  or (_13553_, _13532_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_13554_, _13553_, _13535_);
  or (_13555_, _13537_, _12795_);
  and (_13556_, _13555_, _13554_);
  and (_13557_, _13541_, _13456_);
  or (_40528_, _13557_, _13556_);
  or (_13558_, _13532_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_13559_, _13558_, _13535_);
  or (_13560_, _13537_, _12994_);
  and (_13561_, _13560_, _13559_);
  and (_13562_, _13541_, _13000_);
  or (_40530_, _13562_, _13561_);
  or (_13563_, _13532_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_13564_, _13563_, _13535_);
  or (_13565_, _13537_, _13196_);
  and (_13566_, _13565_, _13564_);
  and (_13567_, _13541_, _13202_);
  or (_40531_, _13567_, _13566_);
  or (_13568_, _13532_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_13569_, _13568_, _13535_);
  or (_13570_, _13537_, _13402_);
  and (_13572_, _13570_, _13569_);
  and (_13573_, _13541_, _13408_);
  or (_40532_, _13573_, _13572_);
  or (_13574_, _13532_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_13575_, _13574_, _13535_);
  or (_13576_, _13537_, _06953_);
  and (_13577_, _13576_, _13575_);
  and (_13578_, _13541_, _06980_);
  or (_40533_, _13578_, _13577_);
  not (_13579_, _05329_);
  and (_13581_, _12003_, _13579_);
  nand (_13582_, _13581_, _04753_);
  and (_13583_, _12190_, _12002_);
  or (_13584_, _13583_, _13582_);
  and (_13585_, _05319_, _05173_);
  and (_13586_, _13585_, _11996_);
  and (_13587_, _13586_, _12181_);
  or (_13588_, _13586_, _04575_);
  nand (_13589_, _13588_, _13582_);
  or (_13590_, _13589_, _13587_);
  and (_40537_, _13590_, _13584_);
  or (_13592_, _13586_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_13593_, _13592_, _13582_);
  not (_13594_, _13586_);
  or (_13595_, _13594_, _12397_);
  and (_13596_, _13595_, _13593_);
  and (_13597_, _12184_, _13579_);
  and (_13598_, _13597_, _04753_);
  and (_13599_, _13598_, _12403_);
  or (_40539_, _13599_, _13596_);
  or (_13601_, _13586_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_13602_, _13601_, _13582_);
  or (_13603_, _13594_, _12599_);
  and (_13604_, _13603_, _13602_);
  and (_13605_, _13598_, _12605_);
  or (_40540_, _13605_, _13604_);
  or (_13606_, _13586_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_13607_, _13606_, _13582_);
  or (_13608_, _13594_, _12795_);
  and (_13609_, _13608_, _13607_);
  and (_13611_, _13598_, _13456_);
  or (_40541_, _13611_, _13609_);
  or (_13612_, _13586_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_13613_, _13612_, _13582_);
  or (_13614_, _13594_, _12994_);
  and (_13615_, _13614_, _13613_);
  and (_13616_, _13598_, _13000_);
  or (_40542_, _13616_, _13615_);
  or (_13617_, _13594_, _13196_);
  or (_13618_, _13586_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_13620_, _13618_, _13582_);
  and (_13621_, _13620_, _13617_);
  and (_13622_, _13598_, _13202_);
  or (_40543_, _13622_, _13621_);
  or (_13623_, _13586_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_13624_, _13623_, _13582_);
  or (_13625_, _13594_, _13402_);
  and (_13626_, _13625_, _13624_);
  and (_13627_, _13598_, _13408_);
  or (_40545_, _13627_, _13626_);
  or (_13629_, _13586_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_13630_, _13629_, _13582_);
  or (_13631_, _13594_, _06953_);
  and (_13632_, _13631_, _13630_);
  and (_13633_, _13598_, _06980_);
  or (_40546_, _13633_, _13632_);
  and (_13634_, _13581_, _05055_);
  not (_13635_, _13634_);
  or (_13636_, _13635_, _13583_);
  and (_13637_, _11995_, _04914_);
  and (_13639_, _13585_, _13637_);
  and (_13640_, _13639_, _12181_);
  nor (_13641_, _13639_, _04577_);
  or (_13642_, _13641_, _13634_);
  or (_13643_, _13642_, _13640_);
  and (_40550_, _13643_, _13636_);
  not (_13644_, _13639_);
  or (_13645_, _13644_, _12397_);
  or (_13646_, _13639_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_13647_, _13646_, _13635_);
  and (_13649_, _13647_, _13645_);
  and (_13650_, _13597_, _05055_);
  and (_13651_, _13650_, _12403_);
  or (_40551_, _13651_, _13649_);
  or (_13652_, _13639_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_13653_, _13652_, _13635_);
  or (_13654_, _13644_, _12599_);
  and (_13655_, _13654_, _13653_);
  and (_13656_, _13650_, _12605_);
  or (_40552_, _13656_, _13655_);
  or (_13658_, _13639_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_13659_, _13658_, _13635_);
  or (_13660_, _13644_, _12795_);
  and (_13661_, _13660_, _13659_);
  and (_13662_, _13650_, _13456_);
  or (_40553_, _13662_, _13661_);
  or (_13663_, _13644_, _12994_);
  or (_13664_, _13639_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_13665_, _13664_, _13635_);
  and (_13666_, _13665_, _13663_);
  and (_13668_, _13650_, _13000_);
  or (_40554_, _13668_, _13666_);
  and (_13669_, _13650_, _13202_);
  or (_13670_, _13639_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_13671_, _13670_, _13635_);
  or (_13672_, _13644_, _13196_);
  and (_13673_, _13672_, _13671_);
  or (_40556_, _13673_, _13669_);
  or (_13674_, _13639_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_13675_, _13674_, _13635_);
  or (_13677_, _13644_, _13402_);
  and (_13678_, _13677_, _13675_);
  and (_13679_, _13650_, _13408_);
  or (_40557_, _13679_, _13678_);
  and (_13680_, _13639_, _06953_);
  nor (_13681_, _13639_, _05468_);
  or (_13682_, _13681_, _13634_);
  or (_13683_, _13682_, _13680_);
  not (_13684_, _13650_);
  or (_13685_, _13684_, _06980_);
  and (_40558_, _13685_, _13683_);
  nor (_13687_, _13416_, _04914_);
  and (_13688_, _13687_, _04749_);
  and (_13689_, _13418_, _05173_);
  and (_13690_, _13689_, _13688_);
  not (_13691_, _13690_);
  or (_13692_, _13691_, _13429_);
  and (_13693_, _13581_, _06151_);
  not (_13694_, _13693_);
  or (_13695_, _13690_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_13697_, _13695_, _13694_);
  and (_13698_, _13697_, _13692_);
  and (_13699_, _13693_, _12191_);
  or (_40562_, _13699_, _13698_);
  or (_13700_, _13690_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_13701_, _13700_, _13694_);
  or (_13702_, _13691_, _13439_);
  and (_13703_, _13702_, _13701_);
  and (_13704_, _13693_, _12403_);
  or (_40563_, _13704_, _13703_);
  or (_13705_, _13690_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_13706_, _13705_, _13694_);
  or (_13707_, _13691_, _13446_);
  and (_13708_, _13707_, _13706_);
  and (_13709_, _13693_, _12605_);
  or (_40564_, _13709_, _13708_);
  or (_13710_, _13690_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_13711_, _13710_, _13694_);
  or (_13712_, _13691_, _13453_);
  and (_13713_, _13712_, _13711_);
  and (_13714_, _13693_, _13456_);
  or (_40565_, _13714_, _13713_);
  or (_13715_, _13691_, _13461_);
  or (_13716_, _13690_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_13717_, _13716_, _13694_);
  and (_13718_, _13717_, _13715_);
  and (_13719_, _13693_, _13000_);
  or (_40566_, _13719_, _13718_);
  or (_13720_, _13690_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_13721_, _13720_, _13694_);
  or (_13722_, _13691_, _13468_);
  and (_13723_, _13722_, _13721_);
  and (_13724_, _13693_, _13202_);
  or (_40568_, _13724_, _13723_);
  or (_13725_, _13690_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_13726_, _13725_, _13694_);
  or (_13727_, _13691_, _13475_);
  and (_13728_, _13727_, _13726_);
  and (_13729_, _13693_, _13408_);
  or (_40569_, _13729_, _13728_);
  or (_13730_, _13690_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_13731_, _13730_, _13694_);
  or (_13732_, _13691_, _13481_);
  and (_13733_, _13732_, _13731_);
  and (_13734_, _13693_, _06980_);
  or (_40570_, _13734_, _13733_);
  nand (_13735_, _13581_, _04752_);
  or (_13736_, _13735_, _13583_);
  and (_13737_, _13585_, _04997_);
  and (_13738_, _13737_, _12181_);
  or (_13739_, _13737_, _04569_);
  nand (_13740_, _13739_, _13735_);
  or (_13741_, _13740_, _13738_);
  and (_40574_, _13741_, _13736_);
  or (_13742_, _13737_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_13743_, _13742_, _13735_);
  not (_13744_, _13737_);
  or (_13745_, _13744_, _12397_);
  and (_13746_, _13745_, _13743_);
  and (_13747_, _13597_, _04752_);
  and (_13748_, _13747_, _12403_);
  or (_40575_, _13748_, _13746_);
  or (_13749_, _13737_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_13750_, _13749_, _13735_);
  or (_13751_, _13744_, _12599_);
  and (_13752_, _13751_, _13750_);
  and (_13753_, _13747_, _12605_);
  or (_40576_, _13753_, _13752_);
  or (_13754_, _13737_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_13755_, _13754_, _13735_);
  or (_13756_, _13744_, _12795_);
  and (_13757_, _13756_, _13755_);
  and (_13758_, _13747_, _13456_);
  or (_40577_, _13758_, _13757_);
  or (_13759_, _13737_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_13760_, _13759_, _13735_);
  or (_13761_, _13744_, _12994_);
  and (_13762_, _13761_, _13760_);
  and (_13763_, _13747_, _13000_);
  or (_40579_, _13763_, _13762_);
  or (_13764_, _13737_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_13765_, _13764_, _13735_);
  or (_13766_, _13744_, _13196_);
  and (_13767_, _13766_, _13765_);
  and (_13768_, _13747_, _13202_);
  or (_40580_, _13768_, _13767_);
  or (_13769_, _13737_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_13770_, _13769_, _13735_);
  or (_13771_, _13744_, _13402_);
  and (_13772_, _13771_, _13770_);
  and (_13773_, _13747_, _13408_);
  or (_40581_, _13773_, _13772_);
  or (_13774_, _13737_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_13775_, _13774_, _13735_);
  or (_13776_, _13744_, _06953_);
  and (_13777_, _13776_, _13775_);
  and (_13778_, _13747_, _06980_);
  or (_40582_, _13778_, _13777_);
  nor (_13779_, _13687_, _13420_);
  and (_13780_, _13417_, _05318_);
  and (_13781_, _13780_, _13779_);
  not (_13782_, _13781_);
  or (_13783_, _13782_, _13429_);
  or (_13784_, _13781_, \oc8051_golden_model_1.IRAM[8] [0]);
  not (_13785_, _05326_);
  and (_13786_, _05335_, _13785_);
  and (_13787_, _13786_, _04753_);
  not (_13788_, _13787_);
  and (_13789_, _13788_, _13784_);
  and (_13790_, _13789_, _13783_);
  and (_13791_, _13787_, _12191_);
  or (_40586_, _13791_, _13790_);
  or (_13792_, _13781_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_13793_, _13792_, _13788_);
  or (_13794_, _13782_, _13439_);
  and (_13795_, _13794_, _13793_);
  and (_13796_, _13787_, _12403_);
  or (_40588_, _13796_, _13795_);
  or (_13797_, _13781_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_13798_, _13797_, _13788_);
  or (_13799_, _13782_, _13446_);
  and (_13800_, _13799_, _13798_);
  and (_13801_, _13787_, _12605_);
  or (_40589_, _13801_, _13800_);
  or (_13802_, _13781_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_13803_, _13802_, _13788_);
  or (_13804_, _13782_, _13453_);
  and (_13805_, _13804_, _13803_);
  and (_13806_, _13787_, _13456_);
  or (_40590_, _13806_, _13805_);
  or (_13807_, _13781_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_13808_, _13807_, _13788_);
  or (_13809_, _13782_, _13461_);
  and (_13810_, _13809_, _13808_);
  and (_13811_, _13787_, _13000_);
  or (_40591_, _13811_, _13810_);
  or (_13812_, _13781_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_13813_, _13812_, _13788_);
  or (_13814_, _13782_, _13468_);
  and (_13815_, _13814_, _13813_);
  and (_13816_, _13787_, _13202_);
  or (_40592_, _13816_, _13815_);
  or (_13817_, _13781_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_13818_, _13817_, _13788_);
  or (_13819_, _13782_, _13475_);
  and (_13820_, _13819_, _13818_);
  and (_13821_, _13787_, _13408_);
  or (_40594_, _13821_, _13820_);
  or (_13822_, _13781_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_13823_, _13822_, _13788_);
  or (_13824_, _13782_, _13481_);
  and (_13825_, _13824_, _13823_);
  and (_13826_, _13787_, _06980_);
  or (_40595_, _13826_, _13825_);
  and (_13827_, _13780_, _13421_);
  not (_13828_, _13827_);
  or (_13829_, _13828_, _13429_);
  or (_13830_, _13827_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_13831_, _13830_, _13829_);
  and (_13832_, _13786_, _05055_);
  or (_13833_, _13832_, _13831_);
  nand (_13834_, _12004_, _05056_);
  or (_13835_, _13834_, _12190_);
  and (_40599_, _13835_, _13833_);
  or (_13836_, _13828_, _13439_);
  or (_13837_, _13827_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_13838_, _13837_, _13834_);
  and (_13839_, _13838_, _13836_);
  and (_13840_, _13832_, _12403_);
  or (_40600_, _13840_, _13839_);
  or (_13841_, _13827_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_13842_, _13841_, _13834_);
  or (_13843_, _13828_, _13446_);
  and (_13844_, _13843_, _13842_);
  and (_13845_, _13832_, _12605_);
  or (_40601_, _13845_, _13844_);
  or (_13846_, _13828_, _13453_);
  or (_13847_, _13827_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_13848_, _13847_, _13834_);
  and (_13849_, _13848_, _13846_);
  and (_13850_, _13832_, _13456_);
  or (_40602_, _13850_, _13849_);
  or (_13851_, _13828_, _13461_);
  or (_13852_, _13827_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_13853_, _13852_, _13834_);
  and (_13854_, _13853_, _13851_);
  and (_13855_, _13832_, _13000_);
  or (_40603_, _13855_, _13854_);
  or (_13856_, _13827_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_13857_, _13856_, _13834_);
  or (_13858_, _13828_, _13468_);
  and (_13859_, _13858_, _13857_);
  and (_13860_, _13832_, _13202_);
  or (_40605_, _13860_, _13859_);
  or (_13861_, _13827_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_13862_, _13861_, _13834_);
  or (_13863_, _13828_, _13475_);
  and (_13864_, _13863_, _13862_);
  and (_13865_, _13832_, _13408_);
  or (_40606_, _13865_, _13864_);
  or (_13866_, _13828_, _13481_);
  or (_13867_, _13827_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_13868_, _13867_, _13834_);
  and (_13869_, _13868_, _13866_);
  and (_13870_, _13832_, _06980_);
  or (_40607_, _13870_, _13869_);
  and (_13871_, _13780_, _13688_);
  or (_13872_, _13871_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_13873_, _13786_, _06151_);
  not (_13874_, _13873_);
  and (_13875_, _13874_, _13872_);
  not (_13876_, _13871_);
  or (_13877_, _13876_, _13429_);
  and (_13878_, _13877_, _13875_);
  and (_13879_, _13873_, _12191_);
  or (_40611_, _13879_, _13878_);
  or (_13880_, _13871_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_13881_, _13880_, _13874_);
  or (_13882_, _13876_, _13439_);
  and (_13883_, _13882_, _13881_);
  and (_13884_, _13873_, _12403_);
  or (_40612_, _13884_, _13883_);
  or (_13885_, _13871_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_13886_, _13885_, _13874_);
  or (_13887_, _13876_, _13446_);
  and (_13888_, _13887_, _13886_);
  and (_13889_, _13873_, _12605_);
  or (_40613_, _13889_, _13888_);
  or (_13890_, _13871_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_13891_, _13890_, _13874_);
  or (_13892_, _13876_, _13453_);
  and (_13893_, _13892_, _13891_);
  and (_13894_, _13873_, _13456_);
  or (_40614_, _13894_, _13893_);
  or (_13895_, _13871_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_13896_, _13895_, _13874_);
  or (_13897_, _13876_, _13461_);
  and (_13898_, _13897_, _13896_);
  and (_13899_, _13873_, _13000_);
  or (_40615_, _13899_, _13898_);
  or (_13900_, _13871_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_13901_, _13900_, _13874_);
  or (_13902_, _13876_, _13468_);
  and (_13903_, _13902_, _13901_);
  and (_13904_, _13873_, _13202_);
  or (_40617_, _13904_, _13903_);
  or (_13905_, _13871_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_13906_, _13905_, _13874_);
  or (_13907_, _13876_, _13475_);
  and (_13908_, _13907_, _13906_);
  and (_13909_, _13873_, _13408_);
  or (_40618_, _13909_, _13908_);
  or (_13910_, _13871_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_13911_, _13910_, _13874_);
  or (_13912_, _13876_, _13481_);
  and (_13913_, _13912_, _13911_);
  and (_13914_, _13873_, _06980_);
  or (_40619_, _13914_, _13913_);
  not (_13915_, _04914_);
  and (_13916_, _13420_, _13915_);
  and (_13917_, _13780_, _13916_);
  not (_13918_, _13917_);
  or (_13919_, _13918_, _13429_);
  and (_13920_, _13786_, _04752_);
  not (_13921_, _13920_);
  or (_13922_, _13917_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_13923_, _13922_, _13921_);
  and (_13924_, _13923_, _13919_);
  and (_13925_, _13920_, _12191_);
  or (_40623_, _13925_, _13924_);
  or (_13926_, _13917_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_13927_, _13926_, _13921_);
  or (_13928_, _13918_, _13439_);
  and (_13929_, _13928_, _13927_);
  and (_13930_, _13920_, _12403_);
  or (_40624_, _13930_, _13929_);
  or (_13931_, _13917_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_13932_, _13931_, _13921_);
  or (_13933_, _13918_, _13446_);
  and (_13934_, _13933_, _13932_);
  and (_13935_, _13920_, _12605_);
  or (_40625_, _13935_, _13934_);
  or (_13936_, _13917_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_13937_, _13936_, _13921_);
  or (_13938_, _13918_, _13453_);
  and (_13939_, _13938_, _13937_);
  and (_13940_, _13920_, _13456_);
  or (_40626_, _13940_, _13939_);
  or (_13941_, _13917_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_13942_, _13941_, _13921_);
  or (_13943_, _13918_, _13461_);
  and (_13944_, _13943_, _13942_);
  and (_13945_, _13920_, _13000_);
  or (_40628_, _13945_, _13944_);
  or (_13946_, _13917_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_13947_, _13946_, _13921_);
  or (_13948_, _13918_, _13468_);
  and (_13949_, _13948_, _13947_);
  and (_13950_, _13920_, _13202_);
  or (_40629_, _13950_, _13949_);
  or (_13951_, _13917_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_13952_, _13951_, _13921_);
  or (_13953_, _13918_, _13475_);
  and (_13954_, _13953_, _13952_);
  and (_13955_, _13920_, _13408_);
  or (_40630_, _13955_, _13954_);
  or (_13956_, _13917_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_13957_, _13956_, _13921_);
  or (_13958_, _13918_, _13481_);
  and (_13959_, _13958_, _13957_);
  and (_13960_, _13920_, _06980_);
  or (_40631_, _13960_, _13959_);
  not (_13961_, _05318_);
  and (_13962_, _13417_, _13961_);
  and (_13963_, _13779_, _13962_);
  not (_13964_, _13963_);
  or (_13965_, _13964_, _13429_);
  and (_13966_, _05336_, _04753_);
  not (_13967_, _13966_);
  or (_13968_, _13963_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_13969_, _13968_, _13967_);
  and (_13970_, _13969_, _13965_);
  and (_13971_, _13966_, _12191_);
  or (_40635_, _13971_, _13970_);
  and (_13972_, _11996_, _05321_);
  or (_13973_, _13972_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_13974_, _13973_, _13967_);
  or (_13975_, _13964_, _13439_);
  and (_13976_, _13975_, _13974_);
  and (_13977_, _13966_, _12403_);
  or (_40636_, _13977_, _13976_);
  or (_13978_, _13972_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_13979_, _13978_, _13967_);
  or (_13980_, _13964_, _13446_);
  and (_13981_, _13980_, _13979_);
  and (_13982_, _13966_, _12605_);
  or (_40637_, _13982_, _13981_);
  or (_13983_, _13972_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_13984_, _13983_, _13967_);
  or (_13985_, _13964_, _13453_);
  and (_13986_, _13985_, _13984_);
  and (_13987_, _13966_, _13456_);
  or (_40639_, _13987_, _13986_);
  or (_13988_, _13972_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_13989_, _13988_, _13967_);
  or (_13990_, _13964_, _13461_);
  and (_13991_, _13990_, _13989_);
  and (_13992_, _13966_, _13000_);
  or (_40640_, _13992_, _13991_);
  or (_13993_, _13972_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_13994_, _13993_, _13967_);
  or (_13995_, _13964_, _13468_);
  and (_13996_, _13995_, _13994_);
  and (_13997_, _13966_, _13202_);
  or (_40641_, _13997_, _13996_);
  or (_13998_, _13972_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_13999_, _13998_, _13967_);
  or (_14000_, _13964_, _13475_);
  and (_14001_, _14000_, _13999_);
  and (_14002_, _13966_, _13408_);
  or (_40642_, _14002_, _14001_);
  or (_14003_, _13972_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_14004_, _14003_, _13967_);
  or (_14005_, _13964_, _13481_);
  and (_14006_, _14005_, _14004_);
  and (_14007_, _13966_, _06980_);
  or (_40643_, _14007_, _14006_);
  and (_14008_, _13421_, _13962_);
  not (_14009_, _14008_);
  or (_14010_, _14009_, _13429_);
  or (_14011_, _14008_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_14012_, _14011_, _14010_);
  and (_14013_, _05336_, _05055_);
  or (_14014_, _14013_, _14012_);
  not (_14015_, _14013_);
  or (_14016_, _14015_, _12191_);
  and (_40647_, _14016_, _14014_);
  and (_14017_, _13637_, _05321_);
  or (_14018_, _14017_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_14019_, _14018_, _14015_);
  or (_14020_, _14009_, _13439_);
  and (_14021_, _14020_, _14019_);
  and (_14022_, _14013_, _12403_);
  or (_40648_, _14022_, _14021_);
  or (_14023_, _14017_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_14024_, _14023_, _14015_);
  or (_14025_, _14009_, _13446_);
  and (_14026_, _14025_, _14024_);
  and (_14027_, _14013_, _12605_);
  or (_40650_, _14027_, _14026_);
  or (_14028_, _14017_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_14029_, _14028_, _14015_);
  or (_14030_, _14009_, _13453_);
  and (_14031_, _14030_, _14029_);
  and (_14032_, _14013_, _13456_);
  or (_40651_, _14032_, _14031_);
  or (_14033_, _14017_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_14034_, _14033_, _14015_);
  or (_14035_, _14009_, _13461_);
  and (_14036_, _14035_, _14034_);
  and (_14037_, _14013_, _13000_);
  or (_40652_, _14037_, _14036_);
  or (_14038_, _14017_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_14039_, _14038_, _14015_);
  or (_14040_, _14009_, _13468_);
  and (_14041_, _14040_, _14039_);
  and (_14042_, _14013_, _13202_);
  or (_40653_, _14042_, _14041_);
  or (_14043_, _14017_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_14044_, _14043_, _14015_);
  or (_14045_, _14009_, _13475_);
  and (_14046_, _14045_, _14044_);
  and (_14047_, _14013_, _13408_);
  or (_40654_, _14047_, _14046_);
  nor (_14048_, _14008_, \oc8051_golden_model_1.IRAM[13] [7]);
  nor (_14049_, _14009_, _13481_);
  or (_14050_, _14049_, _14048_);
  nand (_14051_, _14050_, _14015_);
  or (_14052_, _14015_, _06980_);
  and (_40656_, _14052_, _14051_);
  and (_14053_, _13485_, _05321_);
  or (_14054_, _14053_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_14055_, _06151_, _05336_);
  not (_14056_, _14055_);
  and (_14057_, _14056_, _14054_);
  not (_14058_, _14053_);
  or (_14059_, _14058_, _12181_);
  and (_14060_, _14059_, _14057_);
  and (_14061_, _14055_, _12191_);
  or (_40659_, _14061_, _14060_);
  or (_14062_, _14053_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_14063_, _14062_, _14056_);
  or (_14064_, _14058_, _12397_);
  and (_14065_, _14064_, _14063_);
  and (_14066_, _14055_, _12403_);
  or (_40660_, _14066_, _14065_);
  or (_14067_, _14053_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_14068_, _14067_, _14056_);
  or (_14069_, _14058_, _12599_);
  and (_14070_, _14069_, _14068_);
  and (_14071_, _14055_, _12605_);
  or (_40662_, _14071_, _14070_);
  or (_14072_, _14053_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_14073_, _14072_, _14056_);
  or (_14074_, _14058_, _12795_);
  and (_14075_, _14074_, _14073_);
  and (_14076_, _14055_, _13456_);
  or (_40663_, _14076_, _14075_);
  or (_14077_, _14053_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_14078_, _14077_, _14056_);
  or (_14079_, _14058_, _12994_);
  and (_14080_, _14079_, _14078_);
  and (_14081_, _14055_, _13000_);
  or (_40664_, _14081_, _14080_);
  or (_14082_, _14053_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_14083_, _14082_, _14056_);
  or (_14084_, _14058_, _13196_);
  and (_14085_, _14084_, _14083_);
  and (_14086_, _14055_, _13202_);
  or (_40665_, _14086_, _14085_);
  or (_14087_, _14053_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_14088_, _14087_, _14056_);
  or (_14089_, _14058_, _13402_);
  and (_14090_, _14089_, _14088_);
  and (_14091_, _14055_, _13408_);
  or (_40666_, _14091_, _14090_);
  or (_14092_, _14053_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_14093_, _14092_, _14056_);
  or (_14094_, _14058_, _06953_);
  and (_14095_, _14094_, _14093_);
  and (_14096_, _14055_, _06980_);
  or (_40668_, _14096_, _14095_);
  and (_14097_, _13962_, _13916_);
  not (_14098_, _14097_);
  or (_14099_, _13429_, _14098_);
  or (_14100_, _14097_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_14101_, _14100_, _05338_);
  and (_14102_, _14101_, _14099_);
  and (_14103_, _12191_, _05337_);
  or (_40671_, _14103_, _14102_);
  or (_14104_, _12397_, _05340_);
  or (_14105_, _05322_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_14106_, _14105_, _05338_);
  and (_14107_, _14106_, _14104_);
  and (_14108_, _12403_, _05337_);
  or (_40672_, _14108_, _14107_);
  or (_14109_, _05322_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_14110_, _14109_, _05338_);
  or (_14111_, _12599_, _05340_);
  and (_14112_, _14111_, _14110_);
  and (_14113_, _12605_, _05337_);
  or (_40674_, _14113_, _14112_);
  or (_14114_, _05322_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_14115_, _14114_, _05338_);
  or (_14116_, _12795_, _05340_);
  and (_14117_, _14116_, _14115_);
  and (_14118_, _13456_, _05337_);
  or (_40675_, _14118_, _14117_);
  or (_14119_, _05322_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_14120_, _14119_, _05338_);
  or (_14121_, _12994_, _05340_);
  and (_14122_, _14121_, _14120_);
  and (_14123_, _13000_, _05337_);
  or (_40676_, _14123_, _14122_);
  or (_14124_, _13196_, _05340_);
  or (_14125_, _05322_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_14126_, _14125_, _05338_);
  and (_14127_, _14126_, _14124_);
  and (_14128_, _13202_, _05337_);
  or (_40677_, _14128_, _14127_);
  or (_14129_, _13402_, _05340_);
  or (_14130_, _05322_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_14131_, _14130_, _05338_);
  and (_14132_, _14131_, _14129_);
  and (_14133_, _13408_, _05337_);
  or (_40678_, _14133_, _14132_);
  nor (_14134_, _42908_, _07604_);
  nand (_14135_, _08712_, _05354_);
  nor (_14136_, _05354_, _07604_);
  nor (_14137_, _14136_, _04706_);
  nand (_14138_, _14137_, _14135_);
  and (_14139_, _05354_, _04608_);
  or (_14140_, _14139_, _14136_);
  or (_14141_, _14140_, _04537_);
  nor (_14142_, _05652_, _06988_);
  or (_14143_, _14142_, _14136_);
  or (_14144_, _14143_, _04630_);
  and (_14145_, _05354_, \oc8051_golden_model_1.ACC [0]);
  or (_14146_, _14145_, _14136_);
  and (_14147_, _14146_, _04615_);
  nor (_14148_, _04615_, _07604_);
  or (_14149_, _14148_, _03757_);
  or (_14150_, _14149_, _14147_);
  and (_14151_, _14150_, _03697_);
  and (_14152_, _14151_, _14144_);
  nor (_14153_, _06094_, _07604_);
  and (_14154_, _12032_, _06094_);
  or (_14155_, _14154_, _14153_);
  and (_14156_, _14155_, _03696_);
  or (_14157_, _14156_, _14152_);
  or (_14158_, _14157_, _03755_);
  and (_14159_, _14158_, _14141_);
  or (_14160_, _14159_, _03750_);
  or (_14161_, _14146_, _03751_);
  and (_14162_, _14161_, _03692_);
  and (_14163_, _14162_, _14160_);
  and (_14164_, _14136_, _03691_);
  or (_14165_, _14164_, _03684_);
  or (_14166_, _14165_, _14163_);
  or (_14167_, _14143_, _03685_);
  and (_14168_, _14167_, _14166_);
  or (_14169_, _14168_, _07024_);
  nor (_14170_, _07505_, _07503_);
  nor (_14171_, _14170_, _07506_);
  or (_14172_, _14171_, _07030_);
  and (_14173_, _14172_, _03680_);
  and (_14174_, _14173_, _14169_);
  nand (_14175_, _10753_, _08059_);
  or (_14176_, _14153_, _14175_);
  and (_14177_, _14176_, _03679_);
  and (_14178_, _14177_, _14155_);
  or (_14179_, _14178_, _07544_);
  or (_14180_, _14179_, _14174_);
  or (_14181_, _14140_, _06994_);
  and (_14182_, _14181_, _04679_);
  and (_14183_, _14182_, _14180_);
  and (_14184_, _06935_, _05354_);
  or (_14185_, _14184_, _14136_);
  and (_14186_, _14185_, _04678_);
  or (_14187_, _14186_, _07559_);
  or (_14188_, _14187_, _14183_);
  nor (_14189_, _12119_, _06988_);
  or (_14190_, _14136_, _03415_);
  or (_14191_, _14190_, _14189_);
  and (_14192_, _14191_, _07565_);
  and (_14193_, _14192_, _14188_);
  or (_14194_, _07908_, _07883_);
  or (_14195_, _07914_, _14194_);
  nand (_14196_, _07914_, _03558_);
  and (_14197_, _14196_, _07558_);
  and (_14198_, _14197_, _14195_);
  or (_14199_, _14198_, _08854_);
  or (_14200_, _14199_, _14193_);
  and (_14201_, _12133_, _05354_);
  or (_14202_, _14136_, _04703_);
  or (_14203_, _14202_, _14201_);
  and (_14204_, _05354_, _06428_);
  or (_14205_, _14204_, _14136_);
  or (_14206_, _14205_, _04694_);
  and (_14207_, _14206_, _04701_);
  and (_14208_, _14207_, _14203_);
  and (_14209_, _14208_, _14200_);
  nor (_14210_, _10458_, _06988_);
  or (_14211_, _14210_, _14136_);
  and (_14212_, _14135_, _03959_);
  and (_14213_, _14212_, _14211_);
  or (_14214_, _14213_, _14209_);
  and (_14215_, _14214_, _04708_);
  nand (_14216_, _14205_, _03866_);
  nor (_14217_, _14216_, _14142_);
  or (_14218_, _14217_, _03967_);
  or (_14219_, _14218_, _14215_);
  and (_14220_, _14219_, _14138_);
  or (_14221_, _14220_, _03835_);
  nor (_14222_, _12132_, _06988_);
  or (_14223_, _14136_, _06532_);
  or (_14224_, _14223_, _14222_);
  and (_14225_, _14224_, _06537_);
  and (_14226_, _14225_, _14221_);
  and (_14227_, _14211_, _03954_);
  or (_14228_, _14227_, _03703_);
  or (_14229_, _14228_, _14226_);
  or (_14230_, _14143_, _03704_);
  and (_14231_, _14230_, _14229_);
  or (_14232_, _14231_, _03384_);
  or (_14233_, _14136_, _03385_);
  and (_14234_, _14233_, _14232_);
  or (_14235_, _14234_, _03701_);
  or (_14236_, _14143_, _03702_);
  and (_14237_, _14236_, _42908_);
  and (_14238_, _14237_, _14235_);
  or (_14239_, _14238_, _14134_);
  and (_43136_, _14239_, _41654_);
  nor (_14240_, _42908_, _07568_);
  nor (_14241_, _05354_, _07568_);
  nor (_14242_, _08710_, _06988_);
  or (_14243_, _14242_, _14241_);
  or (_14244_, _14243_, _06537_);
  or (_14245_, _05354_, \oc8051_golden_model_1.B [1]);
  nand (_14246_, _05354_, _04515_);
  and (_14247_, _14246_, _03839_);
  and (_14248_, _14247_, _14245_);
  nor (_14249_, _06094_, _07568_);
  and (_14250_, _12200_, _06094_);
  or (_14251_, _14250_, _14249_);
  and (_14252_, _14251_, _03691_);
  and (_14253_, _05354_, _04813_);
  or (_14254_, _14253_, _14241_);
  or (_14255_, _14254_, _04537_);
  and (_14256_, _12225_, _05354_);
  not (_14257_, _14256_);
  and (_14258_, _14257_, _14245_);
  or (_14259_, _14258_, _04630_);
  and (_14260_, _05354_, \oc8051_golden_model_1.ACC [1]);
  or (_14261_, _14260_, _14241_);
  and (_14262_, _14261_, _04615_);
  nor (_14263_, _04615_, _07568_);
  or (_14264_, _14263_, _03757_);
  or (_14265_, _14264_, _14262_);
  and (_14266_, _14265_, _03697_);
  and (_14267_, _14266_, _14259_);
  and (_14268_, _12212_, _06094_);
  or (_14269_, _14268_, _14249_);
  and (_14270_, _14269_, _03696_);
  or (_14271_, _14270_, _03755_);
  or (_14272_, _14271_, _14267_);
  and (_14273_, _14272_, _14255_);
  or (_14274_, _14273_, _03750_);
  or (_14275_, _14261_, _03751_);
  and (_14276_, _14275_, _03692_);
  and (_14277_, _14276_, _14274_);
  or (_14278_, _14277_, _14252_);
  and (_14279_, _14278_, _03685_);
  and (_14280_, _14268_, _12211_);
  or (_14281_, _14280_, _14249_);
  and (_14282_, _14281_, _03684_);
  or (_14283_, _14282_, _07024_);
  or (_14284_, _14283_, _14279_);
  nor (_14285_, _07508_, _07451_);
  nor (_14286_, _14285_, _07509_);
  or (_14287_, _14286_, _07030_);
  and (_14288_, _14287_, _03680_);
  and (_14289_, _14288_, _14284_);
  nor (_14290_, _12256_, _07545_);
  or (_14291_, _14290_, _14249_);
  and (_14292_, _14291_, _03679_);
  or (_14293_, _14292_, _07544_);
  or (_14294_, _14293_, _14289_);
  or (_14295_, _14254_, _06994_);
  and (_14296_, _14295_, _14294_);
  or (_14297_, _14296_, _04678_);
  and (_14298_, _06934_, _05354_);
  or (_14299_, _14241_, _04679_);
  or (_14300_, _14299_, _14298_);
  and (_14301_, _14300_, _03415_);
  and (_14302_, _14301_, _14297_);
  nand (_14303_, _12313_, _05354_);
  and (_14304_, _14245_, _07559_);
  and (_14305_, _14304_, _14303_);
  or (_14306_, _14305_, _07558_);
  or (_14307_, _14306_, _14302_);
  nor (_14308_, _07909_, _07907_);
  or (_14309_, _14308_, _07910_);
  nor (_14310_, _14309_, _07914_);
  and (_14311_, _07914_, _07880_);
  or (_14312_, _14311_, _14310_);
  or (_14313_, _14312_, _07565_);
  and (_14314_, _14313_, _04694_);
  and (_14315_, _14314_, _14307_);
  or (_14316_, _14315_, _14248_);
  and (_14317_, _14316_, _04703_);
  or (_14318_, _12207_, _06988_);
  and (_14319_, _14245_, _03838_);
  and (_14320_, _14319_, _14318_);
  or (_14321_, _14320_, _03959_);
  or (_14322_, _14321_, _14317_);
  nand (_14323_, _08709_, _05354_);
  and (_14324_, _14323_, _14243_);
  or (_14325_, _14324_, _04701_);
  and (_14326_, _14325_, _04708_);
  and (_14327_, _14326_, _14322_);
  or (_14328_, _12206_, _06988_);
  and (_14329_, _14245_, _03866_);
  and (_14330_, _14329_, _14328_);
  or (_14331_, _14330_, _03967_);
  or (_14332_, _14331_, _14327_);
  nor (_14333_, _14241_, _04706_);
  nand (_14334_, _14333_, _14323_);
  and (_14335_, _14334_, _06532_);
  and (_14336_, _14335_, _14332_);
  or (_14337_, _14246_, _05603_);
  and (_14338_, _14245_, _03835_);
  and (_14339_, _14338_, _14337_);
  or (_14340_, _14339_, _03954_);
  or (_14341_, _14340_, _14336_);
  and (_14342_, _14341_, _14244_);
  or (_14343_, _14342_, _03703_);
  or (_14344_, _14258_, _03704_);
  and (_14345_, _14344_, _03385_);
  and (_14346_, _14345_, _14343_);
  and (_14347_, _14251_, _03384_);
  or (_14348_, _14347_, _03701_);
  or (_14349_, _14348_, _14346_);
  or (_14350_, _14241_, _03702_);
  or (_14351_, _14350_, _14256_);
  and (_14352_, _14351_, _42908_);
  and (_14353_, _14352_, _14349_);
  or (_14354_, _14353_, _14240_);
  and (_43137_, _14354_, _41654_);
  nor (_14355_, _42908_, _07580_);
  nor (_14356_, _05354_, _07580_);
  nor (_14357_, _06988_, _05236_);
  or (_14358_, _14357_, _14356_);
  or (_14359_, _14358_, _06994_);
  and (_14360_, _12419_, _06094_);
  and (_14361_, _14360_, _12418_);
  nor (_14362_, _06094_, _07580_);
  or (_14363_, _14362_, _03685_);
  or (_14364_, _14363_, _14361_);
  or (_14365_, _14358_, _04537_);
  nor (_14366_, _12427_, _06988_);
  or (_14367_, _14366_, _14356_);
  or (_14368_, _14367_, _04630_);
  and (_14369_, _05354_, \oc8051_golden_model_1.ACC [2]);
  or (_14370_, _14369_, _14356_);
  and (_14371_, _14370_, _04615_);
  nor (_14372_, _04615_, _07580_);
  or (_14373_, _14372_, _03757_);
  or (_14374_, _14373_, _14371_);
  and (_14375_, _14374_, _03697_);
  and (_14376_, _14375_, _14368_);
  or (_14377_, _14362_, _14360_);
  and (_14378_, _14377_, _03696_);
  or (_14379_, _14378_, _03755_);
  or (_14380_, _14379_, _14376_);
  and (_14381_, _14380_, _14365_);
  or (_14382_, _14381_, _03750_);
  or (_14383_, _14370_, _03751_);
  and (_14384_, _14383_, _03692_);
  and (_14385_, _14384_, _14382_);
  and (_14386_, _12422_, _06094_);
  or (_14387_, _14386_, _14362_);
  and (_14388_, _14387_, _03691_);
  or (_14389_, _14388_, _03684_);
  or (_14390_, _14389_, _14385_);
  and (_14391_, _14390_, _14364_);
  or (_14392_, _14391_, _07024_);
  or (_14393_, _07510_, _07406_);
  and (_14394_, _14393_, _07511_);
  or (_14395_, _14394_, _07030_);
  and (_14396_, _14395_, _03680_);
  and (_14397_, _14396_, _14392_);
  nor (_14398_, _12465_, _07545_);
  or (_14399_, _14398_, _14362_);
  and (_14400_, _14399_, _03679_);
  or (_14401_, _14400_, _07544_);
  or (_14402_, _14401_, _14397_);
  and (_14403_, _14402_, _14359_);
  or (_14404_, _14403_, _04678_);
  and (_14405_, _06938_, _05354_);
  or (_14406_, _14356_, _04679_);
  or (_14407_, _14406_, _14405_);
  and (_14408_, _14407_, _14404_);
  or (_14409_, _14408_, _07559_);
  nor (_14410_, _12523_, _06988_);
  or (_14411_, _14356_, _03415_);
  or (_14412_, _14411_, _14410_);
  and (_14413_, _14412_, _07565_);
  and (_14414_, _14413_, _14409_);
  nor (_14415_, _07910_, _07881_);
  not (_14416_, _14415_);
  and (_14417_, _14416_, _07873_);
  nor (_14418_, _14416_, _07873_);
  nor (_14419_, _14418_, _14417_);
  or (_14420_, _14419_, _07914_);
  not (_14421_, _07914_);
  or (_14422_, _14421_, _07870_);
  and (_14423_, _14422_, _07558_);
  and (_14424_, _14423_, _14420_);
  or (_14425_, _14424_, _08854_);
  or (_14426_, _14425_, _14414_);
  and (_14427_, _12537_, _05354_);
  or (_14428_, _14356_, _04703_);
  or (_14429_, _14428_, _14427_);
  and (_14430_, _05354_, _06457_);
  or (_14431_, _14430_, _14356_);
  or (_14432_, _14431_, _04694_);
  and (_14433_, _14432_, _04701_);
  and (_14434_, _14433_, _14429_);
  and (_14435_, _14434_, _14426_);
  and (_14436_, _08707_, _05354_);
  or (_14437_, _14436_, _14356_);
  and (_14438_, _14437_, _03959_);
  or (_14439_, _14438_, _14435_);
  and (_14440_, _14439_, _04708_);
  or (_14441_, _14356_, _05700_);
  and (_14442_, _14431_, _03866_);
  and (_14443_, _14442_, _14441_);
  or (_14444_, _14443_, _14440_);
  and (_14445_, _14444_, _04706_);
  and (_14446_, _14370_, _03967_);
  and (_14447_, _14446_, _14441_);
  or (_14448_, _14447_, _03835_);
  or (_14449_, _14448_, _14445_);
  nor (_14450_, _12536_, _06988_);
  or (_14451_, _14356_, _06532_);
  or (_14452_, _14451_, _14450_);
  and (_14453_, _14452_, _06537_);
  and (_14454_, _14453_, _14449_);
  nor (_14455_, _08706_, _06988_);
  or (_14456_, _14455_, _14356_);
  and (_14457_, _14456_, _03954_);
  or (_14458_, _14457_, _03703_);
  or (_14459_, _14458_, _14454_);
  or (_14460_, _14367_, _03704_);
  and (_14461_, _14460_, _03385_);
  and (_14462_, _14461_, _14459_);
  and (_14463_, _14387_, _03384_);
  or (_14464_, _14463_, _03701_);
  or (_14465_, _14464_, _14462_);
  and (_14466_, _12596_, _05354_);
  or (_14467_, _14356_, _03702_);
  or (_14468_, _14467_, _14466_);
  and (_14469_, _14468_, _42908_);
  and (_14470_, _14469_, _14465_);
  or (_14471_, _14470_, _14355_);
  and (_43138_, _14471_, _41654_);
  nor (_14472_, _42908_, _07581_);
  nor (_14473_, _05354_, _07581_);
  nor (_14474_, _12724_, _06988_);
  or (_14475_, _14474_, _14473_);
  and (_14476_, _14475_, _07559_);
  nor (_14477_, _06094_, _07581_);
  and (_14478_, _12619_, _06094_);
  or (_14479_, _14478_, _14477_);
  or (_14480_, _14477_, _12618_);
  and (_14481_, _14480_, _14479_);
  or (_14482_, _14481_, _03685_);
  nor (_14483_, _12610_, _06988_);
  or (_14484_, _14483_, _14473_);
  or (_14485_, _14484_, _04630_);
  and (_14486_, _05354_, \oc8051_golden_model_1.ACC [3]);
  or (_14487_, _14486_, _14473_);
  and (_14488_, _14487_, _04615_);
  nor (_14489_, _04615_, _07581_);
  or (_14490_, _14489_, _03757_);
  or (_14491_, _14490_, _14488_);
  and (_14492_, _14491_, _03697_);
  and (_14493_, _14492_, _14485_);
  and (_14494_, _14479_, _03696_);
  or (_14495_, _14494_, _03755_);
  or (_14496_, _14495_, _14493_);
  nor (_14497_, _06988_, _05050_);
  or (_14498_, _14497_, _14473_);
  or (_14499_, _14498_, _04537_);
  and (_14500_, _14499_, _14496_);
  or (_14501_, _14500_, _03750_);
  or (_14502_, _14487_, _03751_);
  and (_14503_, _14502_, _03692_);
  and (_14504_, _14503_, _14501_);
  and (_14505_, _12622_, _06094_);
  or (_14506_, _14505_, _14477_);
  and (_14507_, _14506_, _03691_);
  or (_14508_, _14507_, _03684_);
  or (_14509_, _14508_, _14504_);
  and (_14510_, _14509_, _14482_);
  or (_14511_, _14510_, _07024_);
  nor (_14512_, _07513_, _07348_);
  nor (_14513_, _14512_, _07514_);
  or (_14514_, _14513_, _07030_);
  and (_14515_, _14514_, _03680_);
  and (_14516_, _14515_, _14511_);
  nor (_14517_, _12665_, _07545_);
  or (_14518_, _14517_, _14477_);
  and (_14519_, _14518_, _03679_);
  or (_14520_, _14519_, _07544_);
  or (_14521_, _14520_, _14516_);
  or (_14522_, _14498_, _06994_);
  and (_14523_, _14522_, _14521_);
  or (_14524_, _14523_, _04678_);
  and (_14525_, _06937_, _05354_);
  or (_14526_, _14473_, _04679_);
  or (_14527_, _14526_, _14525_);
  and (_14528_, _14527_, _03415_);
  and (_14529_, _14528_, _14524_);
  or (_14530_, _14529_, _14476_);
  and (_14531_, _14530_, _07565_);
  nor (_14532_, _14417_, _07872_);
  nor (_14533_, _14532_, _07865_);
  and (_14534_, _14532_, _07865_);
  or (_14535_, _14534_, _14533_);
  or (_14536_, _14535_, _07914_);
  or (_14537_, _14421_, _07862_);
  and (_14538_, _14537_, _07558_);
  and (_14539_, _14538_, _14536_);
  or (_14540_, _14539_, _08854_);
  or (_14541_, _14540_, _14531_);
  and (_14542_, _12738_, _05354_);
  or (_14543_, _14473_, _04703_);
  or (_14544_, _14543_, _14542_);
  and (_14545_, _05354_, _06415_);
  or (_14546_, _14545_, _14473_);
  or (_14547_, _14546_, _04694_);
  and (_14548_, _14547_, _04701_);
  and (_14549_, _14548_, _14544_);
  and (_14550_, _14549_, _14541_);
  and (_14551_, _10455_, _05354_);
  or (_14552_, _14551_, _14473_);
  and (_14553_, _14552_, _03959_);
  or (_14554_, _14553_, _14550_);
  and (_14555_, _14554_, _04708_);
  or (_14556_, _14473_, _05554_);
  and (_14557_, _14546_, _03866_);
  and (_14558_, _14557_, _14556_);
  or (_14559_, _14558_, _14555_);
  and (_14560_, _14559_, _04706_);
  and (_14561_, _14487_, _03967_);
  and (_14562_, _14561_, _14556_);
  or (_14563_, _14562_, _03835_);
  or (_14564_, _14563_, _14560_);
  nor (_14565_, _12737_, _06988_);
  or (_14566_, _14473_, _06532_);
  or (_14567_, _14566_, _14565_);
  and (_14568_, _14567_, _06537_);
  and (_14569_, _14568_, _14564_);
  nor (_14570_, _08701_, _06988_);
  or (_14571_, _14570_, _14473_);
  and (_14572_, _14571_, _03954_);
  or (_14573_, _14572_, _03703_);
  or (_14574_, _14573_, _14569_);
  or (_14575_, _14484_, _03704_);
  and (_14576_, _14575_, _03385_);
  and (_14577_, _14576_, _14574_);
  and (_14578_, _14506_, _03384_);
  or (_14579_, _14578_, _03701_);
  or (_14580_, _14579_, _14577_);
  and (_14581_, _12792_, _05354_);
  or (_14582_, _14473_, _03702_);
  or (_14583_, _14582_, _14581_);
  and (_14584_, _14583_, _42908_);
  and (_14585_, _14584_, _14580_);
  or (_14586_, _14585_, _14472_);
  and (_43139_, _14586_, _41654_);
  nor (_14587_, _42908_, _07706_);
  nor (_14588_, _05354_, _07706_);
  nor (_14589_, _12919_, _06988_);
  or (_14590_, _14589_, _14588_);
  and (_14591_, _14590_, _07559_);
  nor (_14592_, _05898_, _06988_);
  or (_14593_, _14592_, _14588_);
  or (_14594_, _14593_, _06994_);
  nor (_14595_, _06094_, _07706_);
  and (_14596_, _12808_, _06094_);
  or (_14597_, _14596_, _14595_);
  and (_14598_, _14597_, _03691_);
  nor (_14599_, _12828_, _06988_);
  or (_14600_, _14599_, _14588_);
  or (_14601_, _14600_, _04630_);
  and (_14602_, _05354_, \oc8051_golden_model_1.ACC [4]);
  or (_14603_, _14602_, _14588_);
  and (_14604_, _14603_, _04615_);
  nor (_14605_, _04615_, _07706_);
  or (_14606_, _14605_, _03757_);
  or (_14607_, _14606_, _14604_);
  and (_14608_, _14607_, _03697_);
  and (_14609_, _14608_, _14601_);
  and (_14610_, _12832_, _06094_);
  or (_14611_, _14610_, _14595_);
  and (_14612_, _14611_, _03696_);
  or (_14613_, _14612_, _03755_);
  or (_14614_, _14613_, _14609_);
  or (_14615_, _14593_, _04537_);
  and (_14616_, _14615_, _14614_);
  or (_14617_, _14616_, _03750_);
  or (_14618_, _14603_, _03751_);
  and (_14619_, _14618_, _03692_);
  and (_14620_, _14619_, _14617_);
  or (_14621_, _14620_, _14598_);
  and (_14622_, _14621_, _03685_);
  or (_14623_, _14595_, _12847_);
  and (_14624_, _14623_, _03684_);
  and (_14625_, _14624_, _14611_);
  or (_14626_, _14625_, _07024_);
  or (_14627_, _14626_, _14622_);
  or (_14628_, _07517_, _07515_);
  and (_14629_, _14628_, _07518_);
  or (_14630_, _14629_, _07030_);
  and (_14631_, _14630_, _03680_);
  and (_14632_, _14631_, _14627_);
  nor (_14633_, _12810_, _07545_);
  or (_14634_, _14633_, _14595_);
  and (_14635_, _14634_, _03679_);
  or (_14636_, _14635_, _07544_);
  or (_14637_, _14636_, _14632_);
  and (_14638_, _14637_, _14594_);
  or (_14639_, _14638_, _04678_);
  and (_14640_, _06942_, _05354_);
  or (_14641_, _14588_, _04679_);
  or (_14642_, _14641_, _14640_);
  and (_14643_, _14642_, _03415_);
  and (_14644_, _14643_, _14639_);
  or (_14645_, _14644_, _14591_);
  and (_14646_, _14645_, _07565_);
  or (_14647_, _14421_, _07854_);
  nor (_14648_, _14532_, _07864_);
  or (_14649_, _14648_, _07863_);
  nand (_14650_, _14649_, _07901_);
  or (_14651_, _14649_, _07901_);
  and (_14652_, _14651_, _14650_);
  or (_14653_, _14652_, _07914_);
  and (_14654_, _14653_, _07558_);
  and (_14655_, _14654_, _14647_);
  or (_14656_, _14655_, _08854_);
  or (_14657_, _14656_, _14646_);
  and (_14658_, _12933_, _05354_);
  or (_14659_, _14588_, _04703_);
  or (_14660_, _14659_, _14658_);
  and (_14661_, _06422_, _05354_);
  or (_14662_, _14661_, _14588_);
  or (_14663_, _14662_, _04694_);
  and (_14664_, _14663_, _04701_);
  and (_14665_, _14664_, _14660_);
  and (_14666_, _14665_, _14657_);
  and (_14667_, _08700_, _05354_);
  or (_14668_, _14667_, _14588_);
  and (_14669_, _14668_, _03959_);
  or (_14670_, _14669_, _14666_);
  and (_14671_, _14670_, _04708_);
  or (_14672_, _14588_, _08303_);
  and (_14673_, _14662_, _03866_);
  and (_14674_, _14673_, _14672_);
  or (_14675_, _14674_, _14671_);
  and (_14676_, _14675_, _04706_);
  and (_14677_, _14603_, _03967_);
  and (_14678_, _14677_, _14672_);
  or (_14679_, _14678_, _03835_);
  or (_14680_, _14679_, _14676_);
  nor (_14681_, _12931_, _06988_);
  or (_14682_, _14588_, _06532_);
  or (_14683_, _14682_, _14681_);
  and (_14684_, _14683_, _06537_);
  and (_14685_, _14684_, _14680_);
  nor (_14686_, _08699_, _06988_);
  or (_14687_, _14686_, _14588_);
  and (_14688_, _14687_, _03954_);
  or (_14689_, _14688_, _03703_);
  or (_14690_, _14689_, _14685_);
  or (_14691_, _14600_, _03704_);
  and (_14692_, _14691_, _03385_);
  and (_14693_, _14692_, _14690_);
  and (_14694_, _14597_, _03384_);
  or (_14695_, _14694_, _03701_);
  or (_14696_, _14695_, _14693_);
  and (_14697_, _12991_, _05354_);
  or (_14698_, _14588_, _03702_);
  or (_14699_, _14698_, _14697_);
  and (_14700_, _14699_, _42908_);
  and (_14701_, _14700_, _14696_);
  or (_14702_, _14701_, _14587_);
  and (_43140_, _14702_, _41654_);
  nor (_14703_, _42908_, _07697_);
  nor (_14704_, _05354_, _07697_);
  nor (_14705_, _13118_, _06988_);
  or (_14706_, _14705_, _14704_);
  and (_14707_, _14706_, _07559_);
  nor (_14708_, _05799_, _06988_);
  or (_14709_, _14708_, _14704_);
  or (_14710_, _14709_, _06994_);
  nor (_14711_, _06094_, _07697_);
  and (_14712_, _13007_, _06094_);
  or (_14713_, _14712_, _14711_);
  and (_14714_, _14713_, _03691_);
  nor (_14715_, _13025_, _06988_);
  or (_14716_, _14715_, _14704_);
  or (_14717_, _14716_, _04630_);
  and (_14718_, _05354_, \oc8051_golden_model_1.ACC [5]);
  or (_14719_, _14718_, _14704_);
  and (_14720_, _14719_, _04615_);
  nor (_14721_, _04615_, _07697_);
  or (_14722_, _14721_, _03757_);
  or (_14723_, _14722_, _14720_);
  and (_14724_, _14723_, _03697_);
  and (_14725_, _14724_, _14717_);
  and (_14726_, _13029_, _06094_);
  or (_14727_, _14726_, _14711_);
  and (_14728_, _14727_, _03696_);
  or (_14729_, _14728_, _03755_);
  or (_14730_, _14729_, _14725_);
  or (_14731_, _14709_, _04537_);
  and (_14732_, _14731_, _14730_);
  or (_14733_, _14732_, _03750_);
  or (_14734_, _14719_, _03751_);
  and (_14735_, _14734_, _03692_);
  and (_14736_, _14735_, _14733_);
  or (_14737_, _14736_, _14714_);
  and (_14738_, _14737_, _03685_);
  or (_14739_, _14711_, _13044_);
  and (_14740_, _14739_, _03684_);
  and (_14741_, _14740_, _14727_);
  or (_14742_, _14741_, _07024_);
  or (_14743_, _14742_, _14738_);
  or (_14744_, _07221_, _07222_);
  and (_14745_, _14744_, _07519_);
  nor (_14746_, _14745_, _07520_);
  or (_14747_, _14746_, _07030_);
  and (_14748_, _14747_, _03680_);
  and (_14749_, _14748_, _14743_);
  nor (_14750_, _13009_, _07545_);
  or (_14751_, _14750_, _14711_);
  and (_14752_, _14751_, _03679_);
  or (_14753_, _14752_, _07544_);
  or (_14754_, _14753_, _14749_);
  and (_14755_, _14754_, _14710_);
  or (_14756_, _14755_, _04678_);
  and (_14757_, _06941_, _05354_);
  or (_14758_, _14704_, _04679_);
  or (_14759_, _14758_, _14757_);
  and (_14760_, _14759_, _03415_);
  and (_14761_, _14760_, _14756_);
  or (_14762_, _14761_, _14707_);
  and (_14763_, _14762_, _07565_);
  not (_14764_, _07892_);
  and (_14765_, _14650_, _14764_);
  nor (_14766_, _14765_, _07902_);
  and (_14767_, _14765_, _07902_);
  or (_14768_, _14767_, _14766_);
  nor (_14769_, _07914_, _07565_);
  and (_14770_, _14769_, _14768_);
  and (_14771_, _07846_, _07558_);
  and (_14772_, _14771_, _07914_);
  or (_14773_, _14772_, _08854_);
  or (_14774_, _14773_, _14770_);
  or (_14775_, _14774_, _14763_);
  and (_14776_, _13133_, _05354_);
  or (_14777_, _14704_, _04703_);
  or (_14778_, _14777_, _14776_);
  and (_14779_, _06371_, _05354_);
  or (_14780_, _14779_, _14704_);
  or (_14781_, _14780_, _04694_);
  and (_14782_, _14781_, _04701_);
  and (_14783_, _14782_, _14778_);
  and (_14784_, _14783_, _14775_);
  and (_14785_, _10451_, _05354_);
  or (_14786_, _14785_, _14704_);
  and (_14787_, _14786_, _03959_);
  or (_14788_, _14787_, _14784_);
  and (_14789_, _14788_, _04708_);
  or (_14790_, _14704_, _08302_);
  and (_14791_, _14780_, _03866_);
  and (_14792_, _14791_, _14790_);
  or (_14793_, _14792_, _14789_);
  and (_14794_, _14793_, _04706_);
  and (_14795_, _14719_, _03967_);
  and (_14796_, _14795_, _14790_);
  or (_14797_, _14796_, _03835_);
  or (_14798_, _14797_, _14794_);
  nor (_14799_, _13131_, _06988_);
  or (_14800_, _14704_, _06532_);
  or (_14801_, _14800_, _14799_);
  and (_14802_, _14801_, _06537_);
  and (_14803_, _14802_, _14798_);
  nor (_14804_, _08697_, _06988_);
  or (_14805_, _14804_, _14704_);
  and (_14806_, _14805_, _03954_);
  or (_14807_, _14806_, _03703_);
  or (_14808_, _14807_, _14803_);
  or (_14809_, _14716_, _03704_);
  and (_14810_, _14809_, _03385_);
  and (_14811_, _14810_, _14808_);
  and (_14812_, _14713_, _03384_);
  or (_14813_, _14812_, _03701_);
  or (_14814_, _14813_, _14811_);
  and (_14815_, _13193_, _05354_);
  or (_14816_, _14704_, _03702_);
  or (_14817_, _14816_, _14815_);
  and (_14818_, _14817_, _42908_);
  and (_14819_, _14818_, _14814_);
  or (_14820_, _14819_, _14703_);
  and (_43141_, _14820_, _41654_);
  nor (_14821_, _42908_, _07831_);
  nor (_14822_, _05354_, _07831_);
  nor (_14823_, _13326_, _06988_);
  or (_14824_, _14823_, _14822_);
  and (_14825_, _14824_, _07559_);
  nor (_14826_, _06013_, _06988_);
  or (_14827_, _14826_, _14822_);
  or (_14828_, _14827_, _06994_);
  nor (_14829_, _06094_, _07831_);
  and (_14830_, _13218_, _06094_);
  or (_14831_, _14830_, _14829_);
  and (_14832_, _14831_, _03691_);
  nor (_14833_, _13234_, _06988_);
  or (_14834_, _14833_, _14822_);
  or (_14835_, _14834_, _04630_);
  and (_14836_, _05354_, \oc8051_golden_model_1.ACC [6]);
  or (_14837_, _14836_, _14822_);
  and (_14838_, _14837_, _04615_);
  nor (_14839_, _04615_, _07831_);
  or (_14840_, _14839_, _03757_);
  or (_14841_, _14840_, _14838_);
  and (_14842_, _14841_, _03697_);
  and (_14843_, _14842_, _14835_);
  and (_14844_, _13238_, _06094_);
  or (_14845_, _14844_, _14829_);
  and (_14846_, _14845_, _03696_);
  or (_14847_, _14846_, _03755_);
  or (_14848_, _14847_, _14843_);
  or (_14849_, _14827_, _04537_);
  and (_14850_, _14849_, _14848_);
  or (_14851_, _14850_, _03750_);
  or (_14852_, _14837_, _03751_);
  and (_14853_, _14852_, _03692_);
  and (_14854_, _14853_, _14851_);
  or (_14855_, _14854_, _14832_);
  and (_14856_, _14855_, _03685_);
  or (_14857_, _14829_, _13253_);
  and (_14858_, _14845_, _03684_);
  and (_14859_, _14858_, _14857_);
  or (_14860_, _14859_, _07024_);
  or (_14861_, _14860_, _14856_);
  nor (_14862_, _07533_, _07521_);
  nor (_14863_, _14862_, _07534_);
  or (_14864_, _14863_, _07030_);
  and (_14865_, _14864_, _03680_);
  and (_14866_, _14865_, _14861_);
  nor (_14867_, _13220_, _07545_);
  or (_14868_, _14867_, _14829_);
  and (_14869_, _14868_, _03679_);
  or (_14870_, _14869_, _07544_);
  or (_14871_, _14870_, _14866_);
  and (_14872_, _14871_, _14828_);
  or (_14873_, _14872_, _04678_);
  and (_14874_, _06933_, _05354_);
  or (_14875_, _14822_, _04679_);
  or (_14876_, _14875_, _14874_);
  and (_14877_, _14876_, _03415_);
  and (_14878_, _14877_, _14873_);
  or (_14879_, _14878_, _14825_);
  and (_14880_, _14879_, _07565_);
  nor (_14881_, _14765_, _07847_);
  or (_14882_, _14881_, _07848_);
  or (_14883_, _14882_, _07904_);
  nand (_14884_, _14882_, _07904_);
  and (_14885_, _14884_, _14883_);
  or (_14886_, _14885_, _07914_);
  and (_14887_, _07837_, _07558_);
  or (_14888_, _14887_, _14769_);
  and (_14889_, _14888_, _14886_);
  or (_14890_, _14889_, _08854_);
  or (_14891_, _14890_, _14880_);
  and (_14892_, _13341_, _05354_);
  or (_14893_, _14822_, _04703_);
  or (_14894_, _14893_, _14892_);
  and (_14895_, _13333_, _05354_);
  or (_14896_, _14895_, _14822_);
  or (_14897_, _14896_, _04694_);
  and (_14898_, _14897_, _04701_);
  and (_14899_, _14898_, _14894_);
  and (_14900_, _14899_, _14891_);
  and (_14901_, _08695_, _05354_);
  or (_14902_, _14901_, _14822_);
  and (_14903_, _14902_, _03959_);
  or (_14904_, _14903_, _14900_);
  and (_14905_, _14904_, _04708_);
  or (_14906_, _14822_, _08289_);
  and (_14907_, _14896_, _03866_);
  and (_14908_, _14907_, _14906_);
  or (_14909_, _14908_, _14905_);
  and (_14910_, _14909_, _04706_);
  and (_14911_, _14837_, _03967_);
  and (_14912_, _14911_, _14906_);
  or (_14913_, _14912_, _03835_);
  or (_14914_, _14913_, _14910_);
  nor (_14915_, _13340_, _06988_);
  or (_14916_, _14822_, _06532_);
  or (_14917_, _14916_, _14915_);
  and (_14918_, _14917_, _06537_);
  and (_14919_, _14918_, _14914_);
  nor (_14920_, _08694_, _06988_);
  or (_14921_, _14920_, _14822_);
  and (_14922_, _14921_, _03954_);
  or (_14923_, _14922_, _03703_);
  or (_14924_, _14923_, _14919_);
  or (_14925_, _14834_, _03704_);
  and (_14926_, _14925_, _03385_);
  and (_14927_, _14926_, _14924_);
  and (_14928_, _14831_, _03384_);
  or (_14929_, _14928_, _03701_);
  or (_14930_, _14929_, _14927_);
  nor (_14931_, _13399_, _06988_);
  or (_14932_, _14822_, _03702_);
  or (_14933_, _14932_, _14931_);
  and (_14934_, _14933_, _42908_);
  and (_14935_, _14934_, _14930_);
  or (_14936_, _14935_, _14821_);
  and (_43142_, _14936_, _41654_);
  nor (_14937_, _42908_, _03558_);
  and (_14938_, _08777_, \oc8051_golden_model_1.ACC [1]);
  nand (_14939_, _07964_, _06142_);
  and (_14940_, _06698_, _03558_);
  nor (_14941_, _14940_, _07989_);
  or (_14942_, _14941_, _10004_);
  nand (_14943_, _08521_, _14940_);
  nor (_14944_, _08087_, _04353_);
  nor (_14945_, _04608_, \oc8051_golden_model_1.ACC [0]);
  nor (_14946_, _08089_, _04353_);
  nand (_14947_, _14946_, _14945_);
  and (_14948_, _03858_, _03476_);
  and (_14949_, _14948_, _08667_);
  not (_14950_, _14948_);
  and (_14951_, _03799_, _03476_);
  or (_14952_, _04525_, _14951_);
  and (_14953_, _14952_, _08667_);
  nor (_14954_, _05365_, _03558_);
  and (_14955_, _12133_, _05365_);
  nor (_14956_, _14955_, _14954_);
  nand (_14957_, _14956_, _03838_);
  nand (_14958_, _04211_, _03466_);
  nor (_14959_, _12119_, _08094_);
  nor (_14960_, _14959_, _14954_);
  nor (_14961_, _14960_, _03415_);
  and (_14962_, _05365_, _04608_);
  nor (_14963_, _14962_, _14954_);
  nand (_14964_, _14963_, _07544_);
  nor (_14965_, _08061_, _03558_);
  nor (_14966_, _14965_, _08270_);
  nand (_14967_, _14966_, _08260_);
  not (_14968_, _04839_);
  or (_14969_, _14968_, _04608_);
  or (_14970_, _10342_, _04608_);
  nor (_14971_, _04234_, _03558_);
  and (_14972_, _04234_, _03558_);
  or (_14973_, _14972_, _14971_);
  or (_14974_, _14973_, _08105_);
  and (_14975_, _14974_, _08108_);
  and (_14976_, _14975_, _14970_);
  and (_14977_, _14976_, _04625_);
  or (_14978_, _14977_, _06935_);
  or (_14979_, _14976_, _08107_);
  and (_14980_, _14979_, _03450_);
  or (_14981_, _14980_, _04624_);
  and (_14982_, _14981_, _04630_);
  and (_14983_, _14982_, _14978_);
  nor (_14984_, _05652_, _08094_);
  nor (_14985_, _14984_, _14954_);
  nor (_14986_, _14985_, _04630_);
  or (_14987_, _14986_, _03696_);
  or (_14988_, _14987_, _14983_);
  nor (_14989_, _06086_, _03558_);
  and (_14990_, _12032_, _06086_);
  nor (_14991_, _14990_, _14989_);
  nand (_14992_, _14991_, _03696_);
  and (_14993_, _14992_, _04537_);
  and (_14994_, _14993_, _14988_);
  nor (_14995_, _14963_, _04537_);
  or (_14996_, _14995_, _04839_);
  or (_14997_, _14996_, _14994_);
  and (_14998_, _14997_, _14969_);
  or (_14999_, _14998_, _04645_);
  or (_15000_, _06935_, _04646_);
  and (_15001_, _15000_, _03751_);
  and (_15002_, _15001_, _14999_);
  and (_15003_, _05652_, _03750_);
  or (_15004_, _15003_, _08098_);
  or (_15005_, _15004_, _15002_);
  nand (_15006_, _08098_, _07640_);
  and (_15007_, _15006_, _15005_);
  or (_15008_, _15007_, _03691_);
  or (_15009_, _14954_, _03692_);
  and (_15010_, _15009_, _03685_);
  nand (_15011_, _15010_, _15008_);
  or (_15012_, _14985_, _03685_);
  and (_15013_, _15012_, _07030_);
  and (_15014_, _15013_, _15011_);
  not (_15015_, _07484_);
  and (_15016_, _15015_, _07024_);
  or (_15017_, _15016_, _08182_);
  nor (_15018_, _15017_, _15014_);
  nor (_15019_, _08237_, _03558_);
  nor (_15020_, _15019_, _08238_);
  or (_15021_, _15020_, _08181_);
  nand (_15022_, _15021_, _08261_);
  or (_15023_, _15022_, _15018_);
  and (_15024_, _15023_, _14967_);
  or (_15025_, _15024_, _03818_);
  nor (_15026_, _08337_, _03558_);
  nor (_15027_, _15026_, _08338_);
  nand (_15028_, _15027_, _03818_);
  and (_15029_, _15028_, _08288_);
  and (_15030_, _15029_, _15025_);
  nor (_15031_, _08405_, _03558_);
  nor (_15032_, _15031_, _08406_);
  nor (_15033_, _15032_, _08288_);
  or (_15034_, _15033_, _03547_);
  or (_15035_, _15034_, _15030_);
  nand (_15036_, _04211_, _03547_);
  and (_15037_, _15036_, _03680_);
  and (_15038_, _15037_, _15035_);
  nor (_15039_, _12060_, _08432_);
  or (_15040_, _15039_, _14989_);
  and (_15041_, _15040_, _03679_);
  or (_15042_, _15041_, _07544_);
  or (_15043_, _15042_, _15038_);
  and (_15044_, _15043_, _14964_);
  or (_15045_, _15044_, _04678_);
  and (_15046_, _06935_, _05365_);
  nor (_15047_, _15046_, _14954_);
  nand (_15048_, _15047_, _04678_);
  and (_15049_, _15048_, _03415_);
  and (_15050_, _15049_, _15045_);
  or (_15051_, _15050_, _14961_);
  and (_15052_, _15051_, _07565_);
  or (_15053_, _14769_, _03466_);
  or (_15054_, _15053_, _15052_);
  and (_15055_, _15054_, _14958_);
  or (_15056_, _15055_, _03839_);
  and (_15057_, _05365_, _06428_);
  nor (_15058_, _15057_, _14954_);
  nand (_15059_, _15058_, _03839_);
  and (_15060_, _15059_, _08457_);
  and (_15061_, _15060_, _15056_);
  nor (_15062_, _08457_, _04211_);
  or (_15063_, _15062_, _08464_);
  or (_15064_, _15063_, _15061_);
  nor (_15065_, _08667_, _14945_);
  and (_15066_, _08472_, _15065_);
  or (_15067_, _15066_, _10585_);
  and (_15068_, _15067_, _15064_);
  and (_15069_, _08471_, _14941_);
  or (_15070_, _15069_, _03957_);
  or (_15071_, _15070_, _15068_);
  nand (_15072_, _10459_, _03957_);
  and (_15073_, _15072_, _08479_);
  and (_15074_, _15073_, _15071_);
  and (_15075_, _08478_, _10442_);
  or (_15076_, _15075_, _03838_);
  or (_15077_, _15076_, _15074_);
  and (_15078_, _15077_, _14957_);
  or (_15079_, _15078_, _03959_);
  not (_15080_, _14952_);
  or (_15081_, _14954_, _04701_);
  and (_15082_, _15081_, _15080_);
  and (_15083_, _15082_, _15079_);
  or (_15084_, _15083_, _14953_);
  and (_15085_, _15084_, _14950_);
  or (_15086_, _15085_, _14949_);
  and (_15087_, _15086_, _08503_);
  and (_15088_, _08502_, _07989_);
  or (_15089_, _15088_, _03965_);
  or (_15090_, _15089_, _15087_);
  or (_15091_, _08712_, _03966_);
  and (_15092_, _15091_, _08509_);
  and (_15093_, _15092_, _15090_);
  and (_15094_, _08508_, _08748_);
  or (_15095_, _15094_, _15093_);
  and (_15096_, _15095_, _04708_);
  nor (_15097_, _15058_, _14984_);
  and (_15098_, _15097_, _03866_);
  or (_15099_, _15098_, _14946_);
  or (_15100_, _15099_, _15096_);
  and (_15101_, _15100_, _14947_);
  or (_15102_, _15101_, _14944_);
  and (_15103_, _03789_, _03480_);
  or (_15104_, _14945_, _15103_);
  nand (_15105_, _15104_, _10023_);
  and (_15106_, _15105_, _15102_);
  not (_15107_, _15103_);
  nor (_15108_, _14945_, _15107_);
  or (_15109_, _15108_, _08521_);
  or (_15110_, _15109_, _15106_);
  and (_15111_, _15110_, _14943_);
  or (_15112_, _15111_, _03952_);
  nand (_15113_, _10458_, _03952_);
  and (_15114_, _15113_, _08529_);
  and (_15115_, _15114_, _15112_);
  nor (_15116_, _08529_, _10441_);
  or (_15117_, _15116_, _03835_);
  or (_15118_, _15117_, _15115_);
  nor (_15119_, _08540_, _04366_);
  nor (_15120_, _12132_, _08094_);
  nor (_15121_, _15120_, _14954_);
  nand (_15122_, _15121_, _03835_);
  and (_15123_, _15122_, _15119_);
  and (_15124_, _15123_, _15118_);
  nor (_15125_, _15119_, _15020_);
  and (_15126_, _03858_, _03473_);
  or (_15127_, _15126_, _15125_);
  or (_15128_, _15127_, _15124_);
  nand (_15129_, _15126_, _15020_);
  and (_15130_, _15129_, _08080_);
  and (_15131_, _15130_, _15128_);
  nor (_15132_, _14966_, _08080_);
  or (_15133_, _15132_, _03963_);
  or (_15134_, _15133_, _15131_);
  nand (_15135_, _15027_, _03963_);
  and (_15136_, _15135_, _08581_);
  and (_15137_, _15136_, _15134_);
  nor (_15138_, _08581_, _15032_);
  or (_15139_, _15138_, _08006_);
  or (_15140_, _15139_, _15137_);
  nand (_15141_, _08006_, _08059_);
  and (_15142_, _15141_, _08647_);
  and (_15143_, _15142_, _08644_);
  and (_15144_, _15143_, _15140_);
  not (_15145_, _10007_);
  and (_15146_, _15145_, _15065_);
  or (_15147_, _15146_, _07966_);
  or (_15148_, _15147_, _15144_);
  and (_15149_, _15148_, _14942_);
  or (_15150_, _15149_, _03709_);
  nand (_15151_, _10459_, _03709_);
  and (_15152_, _15151_, _08692_);
  and (_15153_, _15152_, _15150_);
  and (_15154_, _08691_, _10442_);
  or (_15155_, _15154_, _07964_);
  or (_15156_, _15155_, _15153_);
  and (_15157_, _15156_, _14939_);
  or (_15158_, _15157_, _03703_);
  nand (_15159_, _14985_, _03703_);
  and (_15160_, _15159_, _08773_);
  and (_15161_, _15160_, _15158_);
  and (_15162_, _08772_, _03558_);
  or (_15163_, _15162_, _15161_);
  and (_15164_, _15163_, _11972_);
  or (_15165_, _15164_, _14938_);
  and (_15166_, _15165_, _03385_);
  and (_15167_, _14954_, _03384_);
  or (_15168_, _15167_, _03701_);
  or (_15169_, _15168_, _15166_);
  nand (_15170_, _14985_, _03701_);
  and (_15171_, _15170_, _08795_);
  and (_15172_, _15171_, _15169_);
  nor (_15173_, _08801_, _03558_);
  nor (_15174_, _15173_, _10917_);
  or (_15175_, _15174_, _15172_);
  nand (_15176_, _08801_, _03491_);
  and (_15177_, _15176_, _42908_);
  and (_15178_, _15177_, _15175_);
  or (_15179_, _15178_, _14937_);
  and (_43143_, _15179_, _41654_);
  nor (_15180_, _42908_, _03491_);
  nand (_15181_, _07964_, _03558_);
  nor (_15182_, _07989_, _07988_);
  nor (_15183_, _15182_, _07990_);
  or (_15184_, _15183_, _10004_);
  and (_15185_, _08617_, _08615_);
  nor (_15186_, _15185_, _08618_);
  or (_15187_, _15186_, _08581_);
  nand (_15188_, _08665_, _08083_);
  and (_15189_, _08664_, _10611_);
  nor (_15190_, _05365_, _03491_);
  and (_15191_, _12207_, _05365_);
  nor (_15192_, _15191_, _15190_);
  nand (_15193_, _15192_, _03838_);
  nand (_15194_, _04482_, _03466_);
  and (_15195_, _05365_, _04813_);
  nor (_15196_, _15195_, _15190_);
  nand (_15197_, _15196_, _07544_);
  and (_15198_, \oc8051_golden_model_1.PSW [7], _03558_);
  and (_15199_, _08059_, \oc8051_golden_model_1.ACC [0]);
  not (_15200_, _15199_);
  and (_15201_, _15200_, _06935_);
  nor (_15202_, _15201_, _15198_);
  and (_15203_, _15202_, _07988_);
  nor (_15204_, _15202_, _07988_);
  or (_15205_, _15204_, _15203_);
  or (_15206_, _15205_, _08261_);
  or (_15207_, _14968_, _04813_);
  or (_15208_, _10342_, _04813_);
  nor (_15209_, _04234_, _03491_);
  and (_15210_, _04234_, _03491_);
  or (_15211_, _15210_, _15209_);
  or (_15212_, _15211_, _08105_);
  and (_15213_, _15212_, _08108_);
  and (_15214_, _15213_, _15208_);
  or (_15215_, _15214_, _08107_);
  and (_15216_, _15215_, _03450_);
  or (_15217_, _15216_, _04624_);
  and (_15218_, _15214_, _04625_);
  or (_15219_, _15218_, _06934_);
  and (_15220_, _15219_, _15217_);
  or (_15221_, _15220_, _03757_);
  nor (_15222_, _05365_, \oc8051_golden_model_1.ACC [1]);
  and (_15223_, _12225_, _05365_);
  nor (_15224_, _15223_, _15222_);
  or (_15225_, _15224_, _04630_);
  and (_15226_, _15225_, _15221_);
  or (_15227_, _15226_, _08120_);
  nor (_15228_, _08128_, \oc8051_golden_model_1.PSW [6]);
  nor (_15229_, _15228_, \oc8051_golden_model_1.ACC [1]);
  and (_15230_, _15228_, \oc8051_golden_model_1.ACC [1]);
  nor (_15231_, _15230_, _15229_);
  nand (_15232_, _15231_, _08120_);
  and (_15233_, _15232_, _03761_);
  and (_15234_, _15233_, _15227_);
  nor (_15235_, _06086_, _03491_);
  and (_15236_, _12212_, _06086_);
  nor (_15237_, _15236_, _15235_);
  nor (_15238_, _15237_, _03697_);
  nor (_15239_, _15196_, _04537_);
  or (_15240_, _15239_, _04839_);
  or (_15241_, _15240_, _15238_);
  or (_15242_, _15241_, _15234_);
  and (_15243_, _15242_, _15207_);
  or (_15244_, _15243_, _04645_);
  or (_15245_, _06934_, _04646_);
  and (_15246_, _15245_, _03751_);
  and (_15247_, _15246_, _15244_);
  nor (_15248_, _05602_, _03751_);
  or (_15249_, _15248_, _08098_);
  or (_15250_, _15249_, _15247_);
  nand (_15251_, _08098_, _07634_);
  and (_15252_, _15251_, _15250_);
  or (_15253_, _15252_, _03691_);
  and (_15254_, _12200_, _06086_);
  nor (_15255_, _15254_, _15235_);
  nand (_15256_, _15255_, _03691_);
  and (_15257_, _15256_, _03685_);
  and (_15258_, _15257_, _15253_);
  and (_15259_, _15236_, _12211_);
  nor (_15260_, _15259_, _15235_);
  nor (_15261_, _15260_, _03685_);
  or (_15262_, _15261_, _07024_);
  or (_15263_, _15262_, _15258_);
  and (_15264_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_15265_, _15264_, _07876_);
  nor (_15266_, _15265_, _07485_);
  or (_15267_, _15266_, _07030_);
  and (_15268_, _15267_, _08181_);
  and (_15269_, _15268_, _15263_);
  and (_15270_, _15200_, _04608_);
  nor (_15271_, _15270_, _15198_);
  and (_15272_, _15271_, _08666_);
  nor (_15273_, _15271_, _08666_);
  or (_15274_, _15273_, _15272_);
  and (_15275_, _15274_, _08182_);
  or (_15276_, _15275_, _08260_);
  or (_15277_, _15276_, _15269_);
  and (_15278_, _15277_, _15206_);
  or (_15279_, _15278_, _03818_);
  and (_15280_, _15200_, _05652_);
  nor (_15281_, _15280_, _15198_);
  and (_15282_, _15281_, _08711_);
  nor (_15283_, _15281_, _08711_);
  or (_15284_, _15283_, _15282_);
  or (_15285_, _15284_, _03823_);
  and (_15286_, _15285_, _08288_);
  and (_15287_, _15286_, _15279_);
  nor (_15288_, _15199_, _04211_);
  nor (_15289_, _15288_, _15198_);
  and (_15290_, _15289_, _08751_);
  nor (_15291_, _15289_, _08751_);
  nor (_15292_, _15291_, _15290_);
  and (_15293_, _15292_, _08287_);
  or (_15294_, _15293_, _03547_);
  or (_15295_, _15294_, _15287_);
  nand (_15296_, _04482_, _03547_);
  and (_15297_, _15296_, _03680_);
  and (_15298_, _15297_, _15295_);
  nor (_15299_, _12256_, _08432_);
  nor (_15300_, _15299_, _15235_);
  nor (_15301_, _15300_, _03680_);
  or (_15302_, _15301_, _07544_);
  or (_15303_, _15302_, _15298_);
  and (_15304_, _15303_, _15197_);
  or (_15305_, _15304_, _04678_);
  and (_15306_, _06934_, _05365_);
  nor (_15307_, _15306_, _15190_);
  nand (_15308_, _15307_, _04678_);
  and (_15309_, _15308_, _03415_);
  and (_15310_, _15309_, _15305_);
  nor (_15311_, _12313_, _08094_);
  nor (_15312_, _15311_, _15190_);
  nor (_15313_, _15312_, _03415_);
  or (_15314_, _15313_, _07558_);
  or (_15315_, _15314_, _15310_);
  nand (_15316_, _07824_, _07558_);
  and (_15317_, _15316_, _15315_);
  or (_15318_, _15317_, _03466_);
  and (_15319_, _15318_, _15194_);
  or (_15320_, _15319_, _03839_);
  and (_15321_, _05365_, _04515_);
  nor (_15322_, _15321_, _15222_);
  or (_15323_, _15322_, _04694_);
  and (_15324_, _15323_, _08457_);
  nand (_15325_, _15324_, _15320_);
  or (_15326_, _08457_, _04482_);
  and (_15327_, _15326_, _08469_);
  nand (_15328_, _15327_, _15325_);
  and (_15329_, _08472_, _08666_);
  or (_15330_, _15329_, _10585_);
  and (_15331_, _15330_, _15328_);
  and (_15332_, _08471_, _07988_);
  or (_15333_, _15332_, _03957_);
  or (_15334_, _15333_, _15331_);
  or (_15335_, _08711_, _03958_);
  and (_15336_, _15335_, _08479_);
  and (_15337_, _15336_, _15334_);
  nor (_15338_, _08479_, _08751_);
  or (_15339_, _15338_, _03838_);
  or (_15340_, _15339_, _15337_);
  and (_15341_, _15340_, _15193_);
  or (_15342_, _15341_, _03959_);
  not (_15343_, _10611_);
  or (_15344_, _15190_, _04701_);
  and (_15345_, _15344_, _15343_);
  and (_15346_, _15345_, _15342_);
  or (_15347_, _15346_, _15189_);
  and (_15348_, _15347_, _08503_);
  and (_15349_, _08502_, _07986_);
  or (_15350_, _15349_, _03965_);
  or (_15351_, _15350_, _15348_);
  or (_15352_, _08709_, _03966_);
  and (_15353_, _15352_, _08509_);
  and (_15354_, _15353_, _15351_);
  and (_15355_, _08508_, _08747_);
  or (_15356_, _15355_, _15354_);
  and (_15357_, _15356_, _04708_);
  and (_15358_, _12206_, _05365_);
  nor (_15359_, _15358_, _15190_);
  nor (_15360_, _15359_, _04708_);
  or (_15361_, _15360_, _08083_);
  or (_15362_, _15361_, _15357_);
  and (_15363_, _15362_, _15188_);
  or (_15364_, _15363_, _08521_);
  nand (_15365_, _08521_, _07987_);
  and (_15366_, _15365_, _03953_);
  and (_15367_, _15366_, _15364_);
  nor (_15368_, _08710_, _03953_);
  or (_15369_, _15368_, _08526_);
  or (_15370_, _15369_, _15367_);
  nand (_15371_, _08526_, _08750_);
  and (_15372_, _15371_, _15370_);
  or (_15373_, _15372_, _03835_);
  nor (_15374_, _12205_, _08094_);
  or (_15375_, _15374_, _15190_);
  or (_15376_, _15375_, _06532_);
  and (_15377_, _15376_, _08547_);
  and (_15378_, _15377_, _15373_);
  not (_15379_, _08547_);
  and (_15380_, _08556_, _08554_);
  nor (_15381_, _15380_, _08557_);
  and (_15382_, _15381_, _15379_);
  or (_15383_, _15382_, _08079_);
  or (_15384_, _15383_, _15378_);
  and (_15385_, _08063_, _08058_);
  nor (_15386_, _15385_, _08064_);
  or (_15387_, _15386_, _08080_);
  and (_15388_, _15387_, _03964_);
  and (_15389_, _15388_, _15384_);
  and (_15390_, _08590_, _08588_);
  nor (_15391_, _15390_, _08591_);
  and (_15392_, _15391_, _03963_);
  or (_15393_, _15392_, _08580_);
  or (_15394_, _15393_, _15389_);
  and (_15395_, _15394_, _15187_);
  or (_15396_, _15395_, _08006_);
  nand (_15397_, _08006_, _03558_);
  and (_15398_, _15397_, _10007_);
  and (_15399_, _15398_, _15396_);
  nor (_15400_, _08667_, _08666_);
  nor (_15401_, _15400_, _08668_);
  and (_15402_, _15401_, _15145_);
  or (_15403_, _15402_, _07966_);
  or (_15404_, _15403_, _15399_);
  and (_15405_, _15404_, _15184_);
  or (_15406_, _15405_, _03709_);
  nor (_15407_, _08712_, _08711_);
  nor (_15408_, _15407_, _08713_);
  or (_15409_, _15408_, _04166_);
  and (_15410_, _15409_, _08692_);
  and (_15411_, _15410_, _15406_);
  and (_15412_, _08751_, _08749_);
  nor (_15413_, _15412_, _08752_);
  and (_15414_, _15413_, _08691_);
  or (_15415_, _15414_, _07964_);
  or (_15416_, _15415_, _15411_);
  and (_15417_, _15416_, _15181_);
  or (_15418_, _15417_, _03703_);
  or (_15419_, _15224_, _03704_);
  and (_15420_, _15419_, _08773_);
  and (_15421_, _15420_, _15418_);
  nor (_15422_, _08802_, _08778_);
  not (_15423_, _15422_);
  and (_15424_, _15423_, _08772_);
  or (_15425_, _15424_, _08777_);
  or (_15426_, _15425_, _15421_);
  nand (_15427_, _08777_, _07740_);
  and (_15428_, _15427_, _03385_);
  and (_15429_, _15428_, _15426_);
  nor (_15430_, _15255_, _03385_);
  or (_15431_, _15430_, _03701_);
  or (_15432_, _15431_, _15429_);
  nor (_15433_, _15223_, _15190_);
  nand (_15434_, _15433_, _03701_);
  and (_15435_, _15434_, _08795_);
  and (_15436_, _15435_, _15432_);
  and (_15437_, _15422_, _08794_);
  or (_15438_, _15437_, _08801_);
  or (_15439_, _15438_, _15436_);
  nand (_15440_, _08801_, _07740_);
  and (_15441_, _15440_, _42908_);
  and (_15442_, _15441_, _15439_);
  or (_15443_, _15442_, _15180_);
  and (_43144_, _15443_, _41654_);
  nor (_15444_, _42908_, _07740_);
  nand (_15445_, _07964_, _03491_);
  nor (_15446_, _05365_, _07740_);
  and (_15447_, _15446_, _03959_);
  or (_15448_, _08479_, _08745_);
  and (_15449_, _03858_, _03485_);
  not (_15450_, _15449_);
  or (_15451_, _15450_, _08662_);
  nand (_15452_, _04165_, _03466_);
  nor (_15453_, _08094_, _05236_);
  nor (_15454_, _15453_, _15446_);
  nand (_15455_, _15454_, _07544_);
  nand (_15456_, _05236_, _04839_);
  nand (_15457_, _08105_, _05236_);
  nor (_15458_, _04234_, _07740_);
  and (_15459_, _04234_, _07740_);
  or (_15460_, _15459_, _15458_);
  or (_15461_, _15460_, _08105_);
  and (_15462_, _15461_, _08108_);
  and (_15463_, _15462_, _15457_);
  or (_15464_, _15463_, _08107_);
  and (_15465_, _15464_, _03450_);
  or (_15466_, _15465_, _04624_);
  and (_15467_, _15463_, _04625_);
  or (_15468_, _15467_, _06938_);
  and (_15469_, _15468_, _15466_);
  and (_15470_, _15469_, _04630_);
  nor (_15471_, _12427_, _08094_);
  nor (_15472_, _15471_, _15446_);
  nor (_15473_, _15472_, _04630_);
  or (_15474_, _15473_, _08120_);
  or (_15475_, _15474_, _15470_);
  and (_15476_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_15477_, _15476_, _08127_);
  nor (_15478_, _15477_, _15228_);
  and (_15479_, _15228_, \oc8051_golden_model_1.ACC [2]);
  nor (_15480_, _15479_, _15478_);
  nand (_15481_, _15480_, _08120_);
  and (_15482_, _15481_, _03761_);
  and (_15483_, _15482_, _15475_);
  nor (_15484_, _06086_, _07740_);
  and (_15485_, _12419_, _06086_);
  nor (_15486_, _15485_, _15484_);
  nor (_15487_, _15486_, _03697_);
  nor (_15488_, _15454_, _04537_);
  or (_15489_, _15488_, _04839_);
  or (_15490_, _15489_, _15487_);
  or (_15491_, _15490_, _15483_);
  and (_15492_, _15491_, _15456_);
  or (_15493_, _15492_, _04645_);
  or (_15494_, _06938_, _04646_);
  and (_15495_, _15494_, _03751_);
  and (_15496_, _15495_, _15493_);
  nor (_15497_, _05699_, _03751_);
  or (_15498_, _15497_, _08098_);
  or (_15499_, _15498_, _15496_);
  nand (_15500_, _08098_, _07586_);
  and (_15501_, _15500_, _15499_);
  or (_15502_, _15501_, _03691_);
  and (_15503_, _12422_, _06086_);
  nor (_15504_, _15503_, _15484_);
  nand (_15505_, _15504_, _03691_);
  and (_15506_, _15505_, _03685_);
  and (_15507_, _15506_, _15502_);
  and (_15508_, _15485_, _12418_);
  nor (_15509_, _15508_, _15484_);
  nor (_15510_, _15509_, _03685_);
  or (_15511_, _15510_, _07024_);
  or (_15512_, _15511_, _15507_);
  nor (_15513_, _07487_, _07485_);
  nor (_15514_, _15513_, _07488_);
  or (_15515_, _15514_, _07030_);
  and (_15516_, _15515_, _08181_);
  and (_15517_, _15516_, _15512_);
  and (_15518_, _04842_, \oc8051_golden_model_1.ACC [1]);
  and (_15519_, _04608_, _03558_);
  nor (_15520_, _15519_, _08666_);
  nor (_15521_, _15520_, _15518_);
  nor (_15522_, _08662_, _15521_);
  and (_15523_, _08662_, _15521_);
  nor (_15524_, _15523_, _15522_);
  nor (_15525_, _15065_, _08666_);
  not (_15526_, _15525_);
  or (_15527_, _15526_, _15524_);
  and (_15528_, _15527_, \oc8051_golden_model_1.PSW [7]);
  nor (_15529_, _15524_, \oc8051_golden_model_1.PSW [7]);
  or (_15530_, _15529_, _15528_);
  nand (_15531_, _15526_, _15524_);
  and (_15532_, _15531_, _15530_);
  nand (_15533_, _15532_, _08261_);
  and (_15534_, _15533_, _10494_);
  or (_15535_, _15534_, _15517_);
  and (_15536_, _06653_, \oc8051_golden_model_1.ACC [1]);
  and (_15537_, _06935_, _03558_);
  nor (_15538_, _15537_, _07988_);
  nor (_15539_, _15538_, _15536_);
  nor (_15540_, _15539_, _07984_);
  and (_15541_, _15539_, _07984_);
  nor (_15542_, _15541_, _15540_);
  nor (_15543_, _14941_, _07988_);
  not (_15544_, _15543_);
  or (_15545_, _15544_, _15542_);
  and (_15546_, _15545_, \oc8051_golden_model_1.PSW [7]);
  nor (_15547_, _15542_, \oc8051_golden_model_1.PSW [7]);
  or (_15548_, _15547_, _15546_);
  nand (_15549_, _15544_, _15542_);
  and (_15550_, _15549_, _15548_);
  nand (_15551_, _15550_, _08260_);
  and (_15552_, _15551_, _15535_);
  or (_15553_, _15552_, _03818_);
  and (_15554_, _05602_, \oc8051_golden_model_1.ACC [1]);
  and (_15555_, _05652_, _03558_);
  nor (_15556_, _11675_, _15555_);
  nor (_15557_, _15556_, _15554_);
  nor (_15558_, _08707_, _15557_);
  and (_15559_, _08707_, _15557_);
  nor (_15560_, _15559_, _15558_);
  not (_15561_, _15560_);
  and (_15562_, _10460_, \oc8051_golden_model_1.PSW [7]);
  and (_15563_, _15562_, _15561_);
  nor (_15564_, _15562_, _15561_);
  nor (_15565_, _15564_, _15563_);
  nand (_15566_, _15565_, _03818_);
  and (_15567_, _15566_, _08288_);
  and (_15568_, _15567_, _15553_);
  nor (_15569_, _04211_, \oc8051_golden_model_1.ACC [0]);
  not (_15570_, _15569_);
  and (_15571_, _08751_, _15570_);
  nor (_15572_, _15571_, _11697_);
  nor (_15573_, _08745_, _15572_);
  and (_15574_, _08745_, _15572_);
  nor (_15575_, _15574_, _15573_);
  not (_15576_, _10444_);
  or (_15577_, _15576_, _15575_);
  and (_15578_, _15577_, \oc8051_golden_model_1.PSW [7]);
  nor (_15579_, _15575_, \oc8051_golden_model_1.PSW [7]);
  or (_15580_, _15579_, _15578_);
  nand (_15581_, _15576_, _15575_);
  and (_15582_, _15581_, _15580_);
  nor (_15583_, _15582_, _08288_);
  or (_15584_, _15583_, _03547_);
  or (_15585_, _15584_, _15568_);
  nand (_15586_, _04165_, _03547_);
  and (_15587_, _15586_, _03680_);
  and (_15588_, _15587_, _15585_);
  nor (_15589_, _12465_, _08432_);
  nor (_15590_, _15589_, _15484_);
  nor (_15591_, _15590_, _03680_);
  or (_15592_, _15591_, _07544_);
  or (_15593_, _15592_, _15588_);
  and (_15594_, _15593_, _15455_);
  or (_15595_, _15594_, _04678_);
  and (_15596_, _06938_, _05365_);
  nor (_15597_, _15596_, _15446_);
  nand (_15598_, _15597_, _04678_);
  and (_15599_, _15598_, _03415_);
  and (_15600_, _15599_, _15595_);
  nor (_15601_, _12523_, _08094_);
  nor (_15602_, _15601_, _15446_);
  nor (_15603_, _15602_, _03415_);
  or (_15604_, _15603_, _07558_);
  or (_15605_, _15604_, _15600_);
  or (_15606_, _07760_, _07565_);
  and (_15607_, _15606_, _15605_);
  or (_15608_, _15607_, _03466_);
  and (_15609_, _15608_, _15452_);
  or (_15610_, _15609_, _03839_);
  and (_15611_, _05365_, _06457_);
  nor (_15612_, _15611_, _15446_);
  nand (_15613_, _15612_, _03839_);
  and (_15614_, _15613_, _08457_);
  and (_15615_, _15614_, _15610_);
  and (_15616_, _04671_, _03485_);
  nor (_15617_, _08457_, _04165_);
  or (_15618_, _15617_, _15616_);
  or (_15619_, _15618_, _15615_);
  not (_15620_, _03485_);
  or (_15621_, _08641_, _15620_);
  not (_15622_, _15616_);
  or (_15623_, _15622_, _08662_);
  and (_15624_, _15623_, _15621_);
  and (_15625_, _15624_, _15619_);
  nor (_15626_, _04674_, _15620_);
  and (_15627_, _15626_, _08662_);
  or (_15628_, _15627_, _15625_);
  and (_15629_, _15628_, _15451_);
  or (_15630_, _15629_, _08471_);
  or (_15631_, _08472_, _07984_);
  and (_15632_, _15631_, _03958_);
  and (_15633_, _15632_, _15630_);
  or (_15634_, _08478_, _08707_);
  and (_15635_, _15634_, _10590_);
  or (_15636_, _15635_, _15633_);
  and (_15637_, _15636_, _15448_);
  or (_15638_, _15637_, _03838_);
  and (_15639_, _12537_, _05365_);
  nor (_15640_, _15639_, _15446_);
  nand (_15641_, _15640_, _03838_);
  and (_15642_, _15641_, _04701_);
  and (_15643_, _15642_, _15638_);
  or (_15644_, _15643_, _15447_);
  and (_15645_, _15644_, _15343_);
  and (_15646_, _08660_, _10611_);
  or (_15647_, _15646_, _15645_);
  and (_15648_, _15647_, _08503_);
  and (_15649_, _08502_, _07982_);
  or (_15650_, _15649_, _03965_);
  or (_15651_, _15650_, _15648_);
  or (_15652_, _08705_, _03966_);
  and (_15653_, _15652_, _08509_);
  and (_15654_, _15653_, _15651_);
  and (_15655_, _08508_, _08743_);
  or (_15656_, _15655_, _15654_);
  and (_15657_, _15656_, _04708_);
  and (_15658_, _03799_, _03480_);
  or (_15659_, _15612_, _08706_);
  nor (_15660_, _15659_, _04708_);
  or (_15661_, _15660_, _15658_);
  or (_15662_, _15661_, _15657_);
  not (_15663_, _08083_);
  nor (_15664_, _08661_, _10022_);
  or (_15665_, _15664_, _15663_);
  and (_15666_, _15665_, _15662_);
  not (_15667_, _08661_);
  and (_15668_, _15667_, _10022_);
  or (_15669_, _15668_, _08521_);
  or (_15670_, _15669_, _15666_);
  nand (_15671_, _08521_, _07983_);
  and (_15672_, _15671_, _03953_);
  and (_15673_, _15672_, _15670_);
  nor (_15674_, _08706_, _03953_);
  or (_15675_, _15674_, _08526_);
  or (_15676_, _15675_, _15673_);
  nand (_15677_, _08526_, _08744_);
  and (_15678_, _15677_, _15676_);
  or (_15679_, _15678_, _03835_);
  nor (_15680_, _12536_, _08094_);
  nor (_15681_, _15680_, _15446_);
  nand (_15682_, _15681_, _03835_);
  and (_15683_, _15682_, _08547_);
  and (_15684_, _15683_, _15679_);
  and (_15685_, _08558_, _08229_);
  nor (_15686_, _15685_, _08559_);
  and (_15687_, _15686_, _15379_);
  or (_15688_, _15687_, _08079_);
  or (_15689_, _15688_, _15684_);
  and (_15690_, _08065_, _08051_);
  nor (_15691_, _15690_, _08066_);
  or (_15692_, _15691_, _08080_);
  and (_15693_, _15692_, _03964_);
  and (_15694_, _15693_, _15689_);
  and (_15695_, _08592_, _08330_);
  nor (_15696_, _15695_, _08593_);
  and (_15697_, _15696_, _03963_);
  or (_15698_, _15697_, _15694_);
  and (_15699_, _15698_, _08581_);
  and (_15700_, _08619_, _08397_);
  nor (_15701_, _15700_, _08620_);
  and (_15702_, _15701_, _08580_);
  or (_15703_, _15702_, _08006_);
  or (_15704_, _15703_, _15699_);
  nand (_15705_, _08006_, _03491_);
  and (_15706_, _15705_, _10007_);
  and (_15707_, _15706_, _15704_);
  and (_15708_, _08669_, _08663_);
  nor (_15709_, _15708_, _08670_);
  and (_15710_, _15709_, _15145_);
  or (_15711_, _15710_, _15707_);
  and (_15712_, _15711_, _10004_);
  and (_15713_, _07991_, _07985_);
  nor (_15714_, _15713_, _07992_);
  and (_15715_, _15714_, _07966_);
  or (_15716_, _15715_, _03709_);
  or (_15717_, _15716_, _15712_);
  and (_15718_, _08714_, _08708_);
  nor (_15719_, _15718_, _08715_);
  or (_15720_, _15719_, _04166_);
  and (_15721_, _15720_, _08692_);
  and (_15722_, _15721_, _15717_);
  and (_15723_, _08753_, _08746_);
  nor (_15724_, _15723_, _08754_);
  and (_15725_, _15724_, _08691_);
  or (_15726_, _15725_, _07964_);
  or (_15727_, _15726_, _15722_);
  and (_15728_, _15727_, _15445_);
  or (_15729_, _15728_, _03703_);
  nand (_15730_, _15472_, _03703_);
  and (_15731_, _15730_, _08773_);
  and (_15732_, _15731_, _15729_);
  and (_15733_, _08127_, _03558_);
  nor (_15734_, _08778_, _07740_);
  or (_15735_, _15734_, _15733_);
  and (_15736_, _15735_, _08772_);
  or (_15737_, _15736_, _08777_);
  or (_15738_, _15737_, _15732_);
  nand (_15739_, _08777_, _07734_);
  and (_15740_, _15739_, _03385_);
  and (_15741_, _15740_, _15738_);
  nor (_15742_, _15504_, _03385_);
  or (_15743_, _15742_, _03701_);
  or (_15744_, _15743_, _15741_);
  and (_15745_, _12596_, _05365_);
  nor (_15746_, _15745_, _15446_);
  nand (_15747_, _15746_, _03701_);
  and (_15748_, _15747_, _08795_);
  and (_15749_, _15748_, _15744_);
  and (_15750_, _08802_, \oc8051_golden_model_1.ACC [2]);
  nor (_15751_, _08802_, \oc8051_golden_model_1.ACC [2]);
  nor (_15752_, _15751_, _15750_);
  and (_15753_, _15752_, _08794_);
  or (_15754_, _15753_, _08801_);
  or (_15755_, _15754_, _15749_);
  nand (_15756_, _08801_, _07734_);
  and (_15757_, _15756_, _42908_);
  and (_15758_, _15757_, _15755_);
  or (_15759_, _15758_, _15444_);
  and (_43145_, _15759_, _41654_);
  nor (_15760_, _42908_, _07734_);
  nor (_15761_, _08658_, _08659_);
  nor (_15762_, _08671_, _15761_);
  and (_15763_, _08671_, _15761_);
  nor (_15764_, _15763_, _15762_);
  nand (_15765_, _15764_, _15145_);
  and (_15766_, _08560_, _08224_);
  nor (_15767_, _15766_, _08561_);
  or (_15768_, _15767_, _08547_);
  nand (_15769_, _08659_, _08083_);
  nor (_15770_, _05365_, _07734_);
  and (_15771_, _12738_, _05365_);
  or (_15772_, _15771_, _15770_);
  or (_15773_, _15772_, _04703_);
  and (_15774_, _03789_, _03485_);
  and (_15775_, _03786_, _03485_);
  nor (_15776_, _15775_, _15616_);
  and (_15777_, _15776_, _15621_);
  or (_15778_, _15777_, _15761_);
  nand (_15779_, _03669_, _03466_);
  nor (_15780_, _08094_, _05050_);
  nor (_15781_, _15780_, _15770_);
  nand (_15782_, _15781_, _07544_);
  and (_15783_, _04165_, \oc8051_golden_model_1.ACC [2]);
  nor (_15784_, _15573_, _15783_);
  nor (_15785_, _10439_, _15784_);
  and (_15786_, _10439_, _15784_);
  nor (_15787_, _15786_, _15785_);
  and (_15788_, _15787_, \oc8051_golden_model_1.PSW [7]);
  nor (_15789_, _15787_, \oc8051_golden_model_1.PSW [7]);
  nor (_15790_, _15789_, _15788_);
  and (_15791_, _15790_, _15578_);
  nor (_15792_, _15790_, _15578_);
  or (_15793_, _15792_, _15791_);
  nand (_15794_, _15793_, _08287_);
  and (_15795_, _05236_, \oc8051_golden_model_1.ACC [2]);
  nor (_15796_, _15522_, _15795_);
  nor (_15797_, _15761_, _15796_);
  and (_15798_, _15761_, _15796_);
  nor (_15799_, _15798_, _15797_);
  and (_15800_, _15799_, \oc8051_golden_model_1.PSW [7]);
  nor (_15801_, _15799_, \oc8051_golden_model_1.PSW [7]);
  nor (_15802_, _15801_, _15800_);
  and (_15803_, _15802_, _15528_);
  nor (_15804_, _15802_, _15528_);
  or (_15805_, _15804_, _15803_);
  nand (_15806_, _15805_, _08182_);
  nor (_15807_, _06086_, _07734_);
  and (_15808_, _12619_, _06086_);
  and (_15809_, _15808_, _12618_);
  nor (_15810_, _15809_, _15807_);
  nor (_15811_, _15810_, _03685_);
  nand (_15812_, _05050_, _04839_);
  nand (_15813_, _08105_, _05050_);
  nor (_15814_, _04234_, _07734_);
  and (_15815_, _04234_, _07734_);
  or (_15816_, _15815_, _15814_);
  or (_15817_, _15816_, _08105_);
  and (_15818_, _15817_, _08108_);
  and (_15819_, _15818_, _15813_);
  and (_15820_, _15819_, _04625_);
  or (_15821_, _15820_, _06937_);
  or (_15822_, _15819_, _08107_);
  and (_15823_, _15822_, _03450_);
  or (_15824_, _15823_, _04624_);
  and (_15825_, _15824_, _04630_);
  and (_15826_, _15825_, _15821_);
  nor (_15827_, _12610_, _08094_);
  nor (_15828_, _15827_, _15770_);
  nor (_15829_, _15828_, _04630_);
  or (_15830_, _15829_, _08120_);
  or (_15831_, _15830_, _15826_);
  not (_15832_, \oc8051_golden_model_1.PSW [6]);
  nor (_15833_, _08127_, _15832_);
  nor (_15834_, _15833_, \oc8051_golden_model_1.ACC [3]);
  nor (_15835_, _15834_, _08128_);
  or (_15836_, _15835_, _11746_);
  and (_15837_, _15836_, _15831_);
  or (_15838_, _15837_, _03696_);
  nor (_15839_, _15808_, _15807_);
  nand (_15840_, _15839_, _03696_);
  and (_15841_, _15840_, _04537_);
  and (_15842_, _15841_, _15838_);
  nor (_15843_, _15781_, _04537_);
  or (_15844_, _15843_, _04839_);
  or (_15845_, _15844_, _15842_);
  and (_15846_, _15845_, _15812_);
  or (_15847_, _15846_, _04645_);
  or (_15848_, _06937_, _04646_);
  and (_15849_, _15848_, _03751_);
  and (_15850_, _15849_, _15847_);
  nor (_15851_, _05553_, _03751_);
  or (_15852_, _15851_, _08098_);
  or (_15853_, _15852_, _15850_);
  nand (_15854_, _08098_, _06142_);
  and (_15855_, _15854_, _15853_);
  or (_15856_, _15855_, _03691_);
  and (_15857_, _12622_, _06086_);
  nor (_15858_, _15857_, _15807_);
  nand (_15859_, _15858_, _03691_);
  and (_15860_, _15859_, _03685_);
  and (_15861_, _15860_, _15856_);
  or (_15862_, _15861_, _15811_);
  and (_15863_, _15862_, _07030_);
  nor (_15864_, _07490_, _07488_);
  nor (_15865_, _15864_, _07491_);
  and (_15866_, _15865_, _07024_);
  or (_15867_, _15866_, _08182_);
  or (_15868_, _15867_, _15863_);
  and (_15869_, _15868_, _15806_);
  or (_15870_, _15869_, _08260_);
  nor (_15871_, _07981_, _07980_);
  and (_15872_, _06789_, \oc8051_golden_model_1.ACC [2]);
  nor (_15873_, _15540_, _15872_);
  nor (_15874_, _15873_, _15871_);
  and (_15875_, _15873_, _15871_);
  nor (_15876_, _15875_, _15874_);
  and (_15877_, _15876_, \oc8051_golden_model_1.PSW [7]);
  nor (_15878_, _15876_, \oc8051_golden_model_1.PSW [7]);
  nor (_15879_, _15878_, _15877_);
  and (_15880_, _15879_, _15546_);
  nor (_15881_, _15879_, _15546_);
  nor (_15882_, _15881_, _15880_);
  or (_15883_, _15882_, _08261_);
  and (_15884_, _15883_, _03823_);
  and (_15885_, _15884_, _15870_);
  nand (_15886_, _10460_, _15561_);
  and (_15887_, _15886_, \oc8051_golden_model_1.PSW [7]);
  and (_15888_, _05699_, \oc8051_golden_model_1.ACC [2]);
  nor (_15889_, _15558_, _15888_);
  nor (_15890_, _10455_, _15889_);
  and (_15891_, _10455_, _15889_);
  nor (_15892_, _15891_, _15890_);
  and (_15893_, _15892_, \oc8051_golden_model_1.PSW [7]);
  nor (_15894_, _15892_, \oc8051_golden_model_1.PSW [7]);
  nor (_15895_, _15894_, _15893_);
  and (_15896_, _15895_, _15887_);
  nor (_15897_, _15895_, _15887_);
  or (_15898_, _15897_, _15896_);
  nor (_15899_, _15898_, _03823_);
  or (_15900_, _15899_, _08287_);
  or (_15901_, _15900_, _15885_);
  and (_15902_, _15901_, _15794_);
  or (_15903_, _15902_, _03547_);
  nand (_15904_, _03669_, _03547_);
  and (_15905_, _15904_, _03680_);
  and (_15906_, _15905_, _15903_);
  nor (_15907_, _12665_, _08432_);
  nor (_15908_, _15907_, _15807_);
  nor (_15909_, _15908_, _03680_);
  or (_15910_, _15909_, _07544_);
  or (_15911_, _15910_, _15906_);
  and (_15912_, _15911_, _15782_);
  or (_15913_, _15912_, _04678_);
  and (_15914_, _06937_, _05365_);
  nor (_15915_, _15914_, _15770_);
  nand (_15916_, _15915_, _04678_);
  and (_15917_, _15916_, _03415_);
  and (_15918_, _15917_, _15913_);
  nor (_15919_, _12724_, _08094_);
  nor (_15920_, _15919_, _15770_);
  nor (_15921_, _15920_, _03415_);
  or (_15922_, _15921_, _07558_);
  or (_15923_, _15922_, _15918_);
  or (_15924_, _07703_, _07565_);
  and (_15925_, _15924_, _15923_);
  or (_15926_, _15925_, _03466_);
  and (_15927_, _15926_, _15779_);
  or (_15928_, _15927_, _03839_);
  and (_15929_, _05365_, _06415_);
  nor (_15930_, _15929_, _15770_);
  nand (_15931_, _15930_, _03839_);
  and (_15932_, _15931_, _08457_);
  and (_15933_, _15932_, _15928_);
  or (_15934_, _08457_, _03669_);
  nand (_15935_, _15934_, _15777_);
  or (_15936_, _15935_, _15933_);
  and (_15937_, _15936_, _15778_);
  or (_15938_, _15937_, _15774_);
  not (_15939_, _15774_);
  or (_15940_, _15761_, _15939_);
  and (_15941_, _15940_, _08472_);
  and (_15942_, _15941_, _15938_);
  and (_15943_, _08471_, _15871_);
  or (_15944_, _15943_, _03957_);
  or (_15945_, _15944_, _15942_);
  or (_15946_, _10455_, _03958_);
  and (_15947_, _15946_, _08479_);
  and (_15948_, _15947_, _15945_);
  and (_15949_, _08478_, _10439_);
  or (_15950_, _15949_, _03838_);
  or (_15951_, _15950_, _15948_);
  and (_15952_, _15951_, _15773_);
  or (_15953_, _15952_, _03959_);
  nor (_15954_, _15770_, _04701_);
  nor (_15955_, _15954_, _08090_);
  and (_15956_, _15955_, _15953_);
  and (_15957_, _08658_, _08496_);
  or (_15958_, _15957_, _15956_);
  not (_15959_, _08658_);
  nand (_15960_, _15959_, _08088_);
  and (_15961_, _15960_, _15958_);
  or (_15962_, _15961_, _08085_);
  or (_15963_, _08658_, _08086_);
  and (_15964_, _15963_, _08503_);
  and (_15965_, _15964_, _15962_);
  and (_15966_, _08502_, _07980_);
  or (_15967_, _15966_, _03965_);
  or (_15968_, _15967_, _15965_);
  or (_15969_, _08703_, _03966_);
  and (_15970_, _15969_, _15968_);
  or (_15971_, _15970_, _08508_);
  or (_15972_, _08509_, _08741_);
  and (_15973_, _15972_, _04708_);
  and (_15974_, _15973_, _15971_);
  or (_15975_, _15930_, _08701_);
  nor (_15976_, _15975_, _04708_);
  or (_15977_, _15976_, _08083_);
  or (_15978_, _15977_, _15974_);
  and (_15979_, _15978_, _15769_);
  or (_15980_, _15979_, _08521_);
  nand (_15981_, _08521_, _07981_);
  and (_15982_, _15981_, _03953_);
  and (_15983_, _15982_, _15980_);
  nor (_15984_, _08701_, _03953_);
  or (_15985_, _15984_, _08526_);
  or (_15986_, _15985_, _15983_);
  nand (_15987_, _08526_, _08742_);
  and (_15988_, _15987_, _06532_);
  and (_15989_, _15988_, _15986_);
  nor (_15990_, _12737_, _08094_);
  nor (_15991_, _15990_, _15770_);
  nor (_15992_, _15991_, _06532_);
  or (_15993_, _15992_, _15379_);
  or (_15994_, _15993_, _15989_);
  and (_15995_, _15994_, _15768_);
  or (_15996_, _15995_, _08079_);
  and (_15997_, _08067_, _08045_);
  nor (_15998_, _15997_, _08068_);
  or (_15999_, _15998_, _08080_);
  and (_16000_, _15999_, _03964_);
  and (_16001_, _16000_, _15996_);
  and (_16002_, _08594_, _08325_);
  nor (_16003_, _16002_, _08595_);
  and (_16004_, _16003_, _03963_);
  or (_16005_, _16004_, _08580_);
  or (_16006_, _16005_, _16001_);
  and (_16007_, _08621_, _08392_);
  nor (_16008_, _16007_, _08622_);
  or (_16009_, _16008_, _08581_);
  and (_16010_, _16009_, _08007_);
  and (_16011_, _16010_, _16006_);
  nand (_16012_, _08006_, \oc8051_golden_model_1.ACC [2]);
  nand (_16013_, _16012_, _10007_);
  or (_16014_, _16013_, _16011_);
  and (_16015_, _16014_, _15765_);
  or (_16016_, _16015_, _07966_);
  nor (_16017_, _15871_, _07993_);
  and (_16018_, _15871_, _07993_);
  nor (_16019_, _16018_, _16017_);
  nand (_16020_, _16019_, _07966_);
  and (_16021_, _16020_, _04166_);
  and (_16022_, _16021_, _16016_);
  nor (_16023_, _08716_, _10455_);
  and (_16024_, _08716_, _10455_);
  nor (_16025_, _16024_, _16023_);
  nor (_16026_, _16025_, _04166_);
  or (_16027_, _16026_, _08691_);
  or (_16028_, _16027_, _16022_);
  nor (_16029_, _08755_, _10439_);
  and (_16030_, _08755_, _10439_);
  nor (_16031_, _16030_, _16029_);
  nand (_16032_, _16031_, _08691_);
  and (_16033_, _16032_, _10870_);
  and (_16034_, _16033_, _16028_);
  and (_16035_, _07964_, \oc8051_golden_model_1.ACC [2]);
  or (_16036_, _16035_, _03703_);
  or (_16037_, _16036_, _16034_);
  nand (_16038_, _15828_, _03703_);
  and (_16039_, _16038_, _08773_);
  and (_16040_, _16039_, _16037_);
  nor (_16041_, _15733_, _07734_);
  or (_16042_, _16041_, _08779_);
  and (_16043_, _16042_, _08772_);
  or (_16044_, _16043_, _08777_);
  or (_16045_, _16044_, _16040_);
  nand (_16046_, _08777_, _07640_);
  and (_16047_, _16046_, _03385_);
  and (_16048_, _16047_, _16045_);
  nor (_16049_, _15858_, _03385_);
  or (_16050_, _16049_, _03701_);
  or (_16051_, _16050_, _16048_);
  and (_16052_, _12792_, _05365_);
  nor (_16053_, _16052_, _15770_);
  nand (_16054_, _16053_, _03701_);
  and (_16055_, _16054_, _08795_);
  and (_16056_, _16055_, _16051_);
  or (_16057_, _15750_, \oc8051_golden_model_1.ACC [3]);
  and (_16058_, _16057_, _08803_);
  and (_16059_, _16058_, _08794_);
  or (_16060_, _16059_, _08801_);
  or (_16061_, _16060_, _16056_);
  nand (_16062_, _08801_, _07640_);
  and (_16063_, _16062_, _42908_);
  and (_16064_, _16063_, _16061_);
  or (_16065_, _16064_, _15760_);
  and (_43146_, _16065_, _41654_);
  nor (_16066_, _42908_, _07640_);
  nand (_16067_, _07964_, _07734_);
  nand (_16068_, _08006_, _07734_);
  nor (_16069_, _08069_, _08037_);
  nor (_16070_, _16069_, _08070_);
  or (_16071_, _16070_, _08080_);
  nand (_16072_, _08526_, _08739_);
  and (_16073_, _14948_, _08655_);
  nor (_16074_, _05365_, _07640_);
  and (_16075_, _12933_, _05365_);
  or (_16076_, _16075_, _16074_);
  or (_16077_, _16076_, _04703_);
  not (_16078_, _04339_);
  or (_16079_, _07979_, _16078_);
  nand (_16080_, _04446_, _03466_);
  nor (_16081_, _05898_, _08094_);
  nor (_16082_, _16081_, _16074_);
  nand (_16083_, _16082_, _07544_);
  nand (_16084_, _05898_, _04839_);
  nand (_16085_, _08105_, _05898_);
  nor (_16086_, _04234_, _07640_);
  and (_16088_, _04234_, _07640_);
  or (_16089_, _16088_, _16086_);
  or (_16090_, _16089_, _08105_);
  and (_16091_, _16090_, _08108_);
  and (_16092_, _16091_, _16085_);
  and (_16093_, _08107_, _06942_);
  or (_16094_, _16093_, _16092_);
  and (_16095_, _16094_, _08118_);
  nor (_16096_, _12828_, _08094_);
  nor (_16097_, _16096_, _16074_);
  nor (_16099_, _16097_, _04630_);
  or (_16100_, _16099_, _08120_);
  or (_16101_, _16100_, _16095_);
  nor (_16102_, _08128_, \oc8051_golden_model_1.ACC [4]);
  nor (_16103_, _16102_, _08134_);
  not (_16104_, _16103_);
  nand (_16105_, _16104_, _08120_);
  and (_16106_, _16105_, _03761_);
  and (_16107_, _16106_, _16101_);
  nor (_16108_, _06086_, _07640_);
  and (_16110_, _12832_, _06086_);
  nor (_16111_, _16110_, _16108_);
  nor (_16112_, _16111_, _03697_);
  nor (_16113_, _16082_, _04537_);
  or (_16114_, _16113_, _04839_);
  or (_16115_, _16114_, _16112_);
  or (_16116_, _16115_, _16107_);
  and (_16117_, _16116_, _16084_);
  or (_16118_, _16117_, _04645_);
  or (_16119_, _06942_, _04646_);
  and (_16121_, _16119_, _03751_);
  and (_16122_, _16121_, _16118_);
  nor (_16123_, _05900_, _03751_);
  or (_16124_, _16123_, _08098_);
  or (_16125_, _16124_, _16122_);
  nand (_16126_, _08098_, _03558_);
  and (_16127_, _16126_, _16125_);
  or (_16128_, _16127_, _03691_);
  and (_16129_, _12808_, _06086_);
  nor (_16130_, _16129_, _16108_);
  nand (_16132_, _16130_, _03691_);
  and (_16133_, _16132_, _03685_);
  and (_16134_, _16133_, _16128_);
  and (_16135_, _16110_, _12847_);
  nor (_16136_, _16135_, _16108_);
  nor (_16137_, _16136_, _03685_);
  or (_16138_, _16137_, _07024_);
  or (_16139_, _16138_, _16134_);
  nor (_16140_, _07493_, _07491_);
  nor (_16141_, _16140_, _07494_);
  or (_16143_, _16141_, _07030_);
  and (_16144_, _16143_, _16139_);
  or (_16145_, _16144_, _08182_);
  or (_16146_, _15803_, _15800_);
  nor (_16147_, _05050_, \oc8051_golden_model_1.ACC [3]);
  nand (_16148_, _05050_, \oc8051_golden_model_1.ACC [3]);
  and (_16149_, _16148_, _15796_);
  or (_16150_, _16149_, _16147_);
  nor (_16151_, _08657_, _16150_);
  and (_16152_, _08657_, _16150_);
  nor (_16154_, _16152_, _16151_);
  and (_16155_, _16154_, \oc8051_golden_model_1.PSW [7]);
  nor (_16156_, _16154_, \oc8051_golden_model_1.PSW [7]);
  nor (_16157_, _16156_, _16155_);
  and (_16158_, _16157_, _16146_);
  nor (_16159_, _16157_, _16146_);
  nor (_16160_, _16159_, _16158_);
  or (_16161_, _16160_, _08181_);
  and (_16162_, _16161_, _16145_);
  or (_16163_, _16162_, _08260_);
  or (_16165_, _15880_, _15877_);
  and (_16166_, _06937_, _07734_);
  or (_16167_, _06937_, _07734_);
  and (_16168_, _15873_, _16167_);
  or (_16169_, _16168_, _16166_);
  nor (_16170_, _16169_, _07979_);
  and (_16171_, _16169_, _07979_);
  nor (_16172_, _16171_, _16170_);
  and (_16173_, _16172_, \oc8051_golden_model_1.PSW [7]);
  nor (_16174_, _16172_, \oc8051_golden_model_1.PSW [7]);
  nor (_16176_, _16174_, _16173_);
  and (_16177_, _16176_, _16165_);
  nor (_16178_, _16176_, _16165_);
  nor (_16179_, _16178_, _16177_);
  or (_16180_, _16179_, _08261_);
  and (_16181_, _16180_, _16163_);
  or (_16182_, _16181_, _03818_);
  or (_16183_, _15896_, _15893_);
  or (_16184_, _15889_, _11671_);
  and (_16185_, _16184_, _11670_);
  nor (_16187_, _08700_, _16185_);
  and (_16188_, _08700_, _16185_);
  nor (_16189_, _16188_, _16187_);
  and (_16190_, _16189_, \oc8051_golden_model_1.PSW [7]);
  nor (_16191_, _16189_, \oc8051_golden_model_1.PSW [7]);
  nor (_16192_, _16191_, _16190_);
  and (_16193_, _16192_, _16183_);
  nor (_16194_, _16192_, _16183_);
  nor (_16195_, _16194_, _16193_);
  or (_16196_, _16195_, _03823_);
  and (_16198_, _16196_, _08288_);
  and (_16199_, _16198_, _16182_);
  or (_16200_, _15791_, _15788_);
  or (_16201_, _15784_, _11703_);
  and (_16202_, _16201_, _11702_);
  nor (_16203_, _08740_, _16202_);
  and (_16204_, _08740_, _16202_);
  nor (_16205_, _16204_, _16203_);
  and (_16206_, _16205_, \oc8051_golden_model_1.PSW [7]);
  nor (_16207_, _16205_, \oc8051_golden_model_1.PSW [7]);
  nor (_16209_, _16207_, _16206_);
  and (_16210_, _16209_, _16200_);
  nor (_16211_, _16209_, _16200_);
  nor (_16212_, _16211_, _16210_);
  and (_16213_, _16212_, _08287_);
  or (_16214_, _16213_, _03547_);
  or (_16215_, _16214_, _16199_);
  nand (_16216_, _04446_, _03547_);
  and (_16217_, _16216_, _03680_);
  and (_16218_, _16217_, _16215_);
  nor (_16220_, _12810_, _08432_);
  nor (_16221_, _16220_, _16108_);
  nor (_16222_, _16221_, _03680_);
  or (_16223_, _16222_, _07544_);
  or (_16224_, _16223_, _16218_);
  and (_16225_, _16224_, _16083_);
  or (_16226_, _16225_, _04678_);
  and (_16227_, _06942_, _05365_);
  nor (_16228_, _16227_, _16074_);
  nand (_16229_, _16228_, _04678_);
  and (_16231_, _16229_, _03415_);
  and (_16232_, _16231_, _16226_);
  nor (_16233_, _12919_, _08094_);
  nor (_16234_, _16233_, _16074_);
  nor (_16235_, _16234_, _03415_);
  or (_16236_, _16235_, _07558_);
  or (_16237_, _16236_, _16232_);
  or (_16238_, _07649_, _07565_);
  and (_16239_, _16238_, _16237_);
  or (_16240_, _16239_, _03466_);
  and (_16242_, _16240_, _16080_);
  or (_16243_, _16242_, _03839_);
  and (_16244_, _06422_, _05365_);
  nor (_16245_, _16244_, _16074_);
  nand (_16246_, _16245_, _03839_);
  and (_16247_, _16246_, _08457_);
  and (_16248_, _16247_, _16243_);
  nor (_16249_, _08457_, _04446_);
  or (_16250_, _16249_, _15616_);
  or (_16251_, _16250_, _16248_);
  or (_16253_, _15622_, _08657_);
  and (_16254_, _16253_, _15621_);
  and (_16255_, _16254_, _16251_);
  or (_16256_, _15449_, _08657_);
  and (_16257_, _16256_, _15626_);
  or (_16258_, _16257_, _16255_);
  and (_16259_, _12353_, _03485_);
  not (_16260_, _16259_);
  or (_16261_, _15450_, _08657_);
  and (_16262_, _16261_, _16260_);
  and (_16263_, _16262_, _16258_);
  or (_16264_, _07979_, _03349_);
  and (_16265_, _16264_, _08471_);
  or (_16266_, _16265_, _16263_);
  and (_16267_, _16266_, _16079_);
  or (_16268_, _16267_, _03957_);
  or (_16269_, _08700_, _03958_);
  and (_16270_, _16269_, _08479_);
  and (_16271_, _16270_, _16268_);
  and (_16272_, _08478_, _08740_);
  or (_16274_, _16272_, _03838_);
  or (_16275_, _16274_, _16271_);
  and (_16276_, _16275_, _16077_);
  or (_16277_, _16276_, _03959_);
  nor (_16278_, _16074_, _04701_);
  nor (_16279_, _16278_, _14951_);
  and (_16280_, _16279_, _16277_);
  and (_16281_, _08655_, _14951_);
  or (_16282_, _16281_, _04525_);
  or (_16283_, _16282_, _16280_);
  not (_16285_, _04525_);
  or (_16286_, _08655_, _16285_);
  and (_16287_, _16286_, _14950_);
  and (_16288_, _16287_, _16283_);
  or (_16289_, _16288_, _16073_);
  and (_16290_, _16289_, _08503_);
  and (_16291_, _08502_, _07977_);
  or (_16292_, _16291_, _03965_);
  or (_16293_, _16292_, _16290_);
  or (_16294_, _08698_, _03966_);
  and (_16296_, _16294_, _08509_);
  and (_16297_, _16296_, _16293_);
  and (_16298_, _08508_, _08738_);
  or (_16299_, _16298_, _16297_);
  and (_16300_, _16299_, _04708_);
  or (_16301_, _16245_, _08699_);
  nor (_16302_, _16301_, _04708_);
  or (_16303_, _16302_, _15658_);
  or (_16304_, _16303_, _16300_);
  nor (_16305_, _08656_, _03412_);
  or (_16307_, _16305_, _15663_);
  and (_16308_, _16307_, _16304_);
  not (_16309_, _10022_);
  nor (_16310_, _08656_, _16309_);
  or (_16311_, _16310_, _08521_);
  or (_16312_, _16311_, _16308_);
  nand (_16313_, _08521_, _07978_);
  and (_16314_, _16313_, _03953_);
  and (_16315_, _16314_, _16312_);
  nand (_16316_, _08529_, _08699_);
  and (_16318_, _16316_, _08528_);
  or (_16319_, _16318_, _16315_);
  and (_16320_, _16319_, _16072_);
  or (_16321_, _16320_, _03835_);
  nor (_16322_, _12931_, _08094_);
  nor (_16323_, _16322_, _16074_);
  nand (_16324_, _16323_, _03835_);
  and (_16325_, _16324_, _08547_);
  and (_16326_, _16325_, _16321_);
  nor (_16327_, _08562_, _08214_);
  nor (_16329_, _16327_, _08563_);
  and (_16330_, _16329_, _15379_);
  or (_16331_, _16330_, _08079_);
  or (_16332_, _16331_, _16326_);
  and (_16333_, _16332_, _16071_);
  or (_16334_, _16333_, _03963_);
  nor (_16335_, _08596_, _08319_);
  nor (_16336_, _16335_, _08597_);
  or (_16337_, _16336_, _03964_);
  and (_16338_, _16337_, _08581_);
  and (_16340_, _16338_, _16334_);
  nor (_16341_, _08623_, _08386_);
  nor (_16342_, _16341_, _08624_);
  and (_16343_, _16342_, _08580_);
  or (_16344_, _16343_, _08006_);
  or (_16345_, _16344_, _16340_);
  and (_16346_, _16345_, _16068_);
  or (_16347_, _16346_, _15145_);
  nor (_16348_, _08673_, _08657_);
  nor (_16349_, _16348_, _08674_);
  or (_16351_, _16349_, _10007_);
  and (_16352_, _16351_, _10004_);
  and (_16353_, _16352_, _16347_);
  nor (_16354_, _07995_, _07979_);
  nor (_16355_, _16354_, _07996_);
  and (_16356_, _16355_, _07966_);
  or (_16357_, _16356_, _03709_);
  or (_16358_, _16357_, _16353_);
  nor (_16359_, _08718_, _08700_);
  nor (_16360_, _16359_, _08719_);
  or (_16362_, _16360_, _04166_);
  and (_16363_, _16362_, _08692_);
  and (_16364_, _16363_, _16358_);
  nor (_16365_, _08757_, _08740_);
  nor (_16366_, _16365_, _08758_);
  and (_16367_, _16366_, _08691_);
  or (_16368_, _16367_, _07964_);
  or (_16369_, _16368_, _16364_);
  and (_16370_, _16369_, _16067_);
  or (_16371_, _16370_, _03703_);
  nand (_16373_, _16097_, _03703_);
  and (_16374_, _16373_, _08773_);
  and (_16375_, _16374_, _16371_);
  and (_16376_, _08779_, _07640_);
  nor (_16377_, _08779_, _07640_);
  nor (_16378_, _16377_, _16376_);
  not (_16379_, _16378_);
  nor (_16380_, _16379_, _08777_);
  nor (_16381_, _16380_, _10894_);
  or (_16382_, _16381_, _16375_);
  nand (_16384_, _08777_, _07634_);
  and (_16385_, _16384_, _03385_);
  and (_16386_, _16385_, _16382_);
  nor (_16387_, _16130_, _03385_);
  or (_16388_, _16387_, _03701_);
  or (_16389_, _16388_, _16386_);
  and (_16390_, _12991_, _05365_);
  nor (_16391_, _16390_, _16074_);
  nand (_16392_, _16391_, _03701_);
  and (_16393_, _16392_, _08795_);
  and (_16395_, _16393_, _16389_);
  and (_16396_, _08803_, _07640_);
  nor (_16397_, _16396_, _08804_);
  and (_16398_, _16397_, _08794_);
  or (_16399_, _16398_, _08801_);
  or (_16400_, _16399_, _16395_);
  nand (_16401_, _08801_, _07634_);
  and (_16402_, _16401_, _42908_);
  and (_16403_, _16402_, _16400_);
  or (_16404_, _16403_, _16066_);
  and (_43147_, _16404_, _41654_);
  nor (_16406_, _42908_, _07634_);
  and (_16407_, _08675_, _08654_);
  nor (_16408_, _16407_, _08676_);
  or (_16409_, _16408_, _10007_);
  and (_16410_, _08564_, _08206_);
  nor (_16411_, _16410_, _08565_);
  or (_16412_, _16411_, _08547_);
  nand (_16413_, _03858_, _03480_);
  and (_16414_, _06991_, _03480_);
  nand (_16416_, _08652_, _16414_);
  and (_16417_, _16416_, _16413_);
  nor (_16418_, _05365_, _07634_);
  and (_16419_, _13133_, _05365_);
  nor (_16420_, _16419_, _16418_);
  nand (_16421_, _16420_, _03838_);
  nand (_16422_, _04034_, _03466_);
  nor (_16423_, _05799_, _08094_);
  nor (_16424_, _16423_, _16418_);
  nand (_16425_, _16424_, _07544_);
  and (_16427_, _04446_, \oc8051_golden_model_1.ACC [4]);
  nor (_16428_, _16203_, _16427_);
  nor (_16429_, _08736_, _16428_);
  and (_16430_, _08736_, _16428_);
  nor (_16431_, _16430_, _16429_);
  and (_16432_, _16431_, \oc8051_golden_model_1.PSW [7]);
  nor (_16433_, _16431_, \oc8051_golden_model_1.PSW [7]);
  nor (_16434_, _16433_, _16432_);
  nor (_16435_, _16210_, _16206_);
  not (_16436_, _16435_);
  and (_16438_, _16436_, _16434_);
  nor (_16439_, _16436_, _16434_);
  nor (_16440_, _16439_, _16438_);
  or (_16441_, _16440_, _08288_);
  and (_16442_, _05898_, \oc8051_golden_model_1.ACC [4]);
  nor (_16443_, _16151_, _16442_);
  and (_16444_, _08654_, _16443_);
  nor (_16445_, _08654_, _16443_);
  nor (_16446_, _16445_, _16444_);
  nor (_16447_, _16446_, _08059_);
  and (_16449_, _16446_, _08059_);
  nor (_16450_, _16449_, _16447_);
  nor (_16451_, _16158_, _16155_);
  not (_16452_, _16451_);
  and (_16453_, _16452_, _16450_);
  nor (_16454_, _16452_, _16450_);
  nor (_16455_, _16454_, _16453_);
  or (_16456_, _16455_, _08181_);
  nor (_16457_, _06086_, _07634_);
  and (_16458_, _13029_, _06086_);
  and (_16461_, _16458_, _13044_);
  nor (_16462_, _16461_, _16457_);
  nor (_16463_, _16462_, _03685_);
  nand (_16464_, _05799_, _04839_);
  nand (_16465_, _08105_, _05799_);
  nor (_16466_, _04234_, _07634_);
  and (_16467_, _04234_, _07634_);
  or (_16468_, _16467_, _16466_);
  or (_16469_, _16468_, _08105_);
  and (_16470_, _16469_, _08108_);
  and (_16472_, _16470_, _16465_);
  and (_16473_, _08107_, _06941_);
  or (_16474_, _16473_, _16472_);
  and (_16475_, _16474_, _08118_);
  nor (_16476_, _13025_, _08094_);
  nor (_16477_, _16476_, _16418_);
  nor (_16478_, _16477_, _04630_);
  or (_16479_, _16478_, _08120_);
  or (_16480_, _16479_, _16475_);
  and (_16481_, _11757_, _08136_);
  nor (_16483_, _11757_, _08136_);
  nor (_16484_, _16483_, _16481_);
  nand (_16485_, _16484_, _08120_);
  and (_16486_, _16485_, _03761_);
  and (_16487_, _16486_, _16480_);
  nor (_16488_, _16458_, _16457_);
  nor (_16489_, _16488_, _03697_);
  nor (_16490_, _16424_, _04537_);
  or (_16491_, _16490_, _04839_);
  or (_16492_, _16491_, _16489_);
  or (_16494_, _16492_, _16487_);
  and (_16495_, _16494_, _16464_);
  or (_16496_, _16495_, _04645_);
  or (_16497_, _06941_, _04646_);
  and (_16498_, _16497_, _03751_);
  and (_16499_, _16498_, _16496_);
  nor (_16500_, _05801_, _03751_);
  or (_16501_, _16500_, _08098_);
  or (_16502_, _16501_, _16499_);
  nand (_16503_, _08098_, _03491_);
  and (_16505_, _16503_, _16502_);
  or (_16506_, _16505_, _03691_);
  and (_16507_, _13007_, _06086_);
  nor (_16508_, _16507_, _16457_);
  nand (_16509_, _16508_, _03691_);
  and (_16510_, _16509_, _03685_);
  and (_16511_, _16510_, _16506_);
  or (_16512_, _16511_, _16463_);
  and (_16513_, _16512_, _07030_);
  nor (_16514_, _07496_, _07494_);
  nor (_16516_, _16514_, _07497_);
  and (_16517_, _16516_, _07024_);
  or (_16518_, _16517_, _08182_);
  or (_16519_, _16518_, _16513_);
  and (_16520_, _16519_, _16456_);
  or (_16521_, _16520_, _08260_);
  and (_16522_, _06881_, \oc8051_golden_model_1.ACC [4]);
  nor (_16523_, _16170_, _16522_);
  nor (_16524_, _16523_, _07976_);
  and (_16525_, _16523_, _07976_);
  nor (_16527_, _16525_, _16524_);
  nor (_16528_, _16527_, _08059_);
  and (_16529_, _16527_, _08059_);
  nor (_16530_, _16529_, _16528_);
  nor (_16531_, _16177_, _16173_);
  not (_16532_, _16531_);
  and (_16533_, _16532_, _16530_);
  nor (_16534_, _16532_, _16530_);
  nor (_16535_, _16534_, _16533_);
  or (_16536_, _16535_, _08261_);
  and (_16538_, _16536_, _03823_);
  and (_16539_, _16538_, _16521_);
  and (_16540_, _05900_, \oc8051_golden_model_1.ACC [4]);
  nor (_16541_, _16187_, _16540_);
  nor (_16542_, _10451_, _16541_);
  and (_16543_, _10451_, _16541_);
  nor (_16544_, _16543_, _16542_);
  and (_16545_, _16544_, \oc8051_golden_model_1.PSW [7]);
  nor (_16546_, _16544_, \oc8051_golden_model_1.PSW [7]);
  nor (_16547_, _16546_, _16545_);
  nor (_16549_, _16193_, _16190_);
  not (_16550_, _16549_);
  and (_16551_, _16550_, _16547_);
  nor (_16552_, _16550_, _16547_);
  nor (_16553_, _16552_, _16551_);
  and (_16554_, _16553_, _03818_);
  or (_16555_, _16554_, _08287_);
  or (_16556_, _16555_, _16539_);
  and (_16557_, _16556_, _16441_);
  or (_16558_, _16557_, _03547_);
  nand (_16560_, _04034_, _03547_);
  and (_16561_, _16560_, _03680_);
  and (_16562_, _16561_, _16558_);
  nor (_16563_, _13009_, _08432_);
  nor (_16564_, _16563_, _16457_);
  nor (_16565_, _16564_, _03680_);
  or (_16566_, _16565_, _07544_);
  or (_16567_, _16566_, _16562_);
  and (_16568_, _16567_, _16425_);
  or (_16569_, _16568_, _04678_);
  and (_16571_, _06941_, _05365_);
  nor (_16572_, _16571_, _16418_);
  nand (_16573_, _16572_, _04678_);
  and (_16574_, _16573_, _03415_);
  and (_16575_, _16574_, _16569_);
  nor (_16576_, _13118_, _08094_);
  nor (_16577_, _16576_, _16418_);
  nor (_16578_, _16577_, _03415_);
  or (_16579_, _16578_, _07558_);
  or (_16580_, _16579_, _16575_);
  or (_16582_, _07619_, _07565_);
  and (_16583_, _16582_, _16580_);
  or (_16584_, _16583_, _03466_);
  and (_16585_, _16584_, _16422_);
  or (_16586_, _16585_, _03839_);
  and (_16587_, _06371_, _05365_);
  nor (_16588_, _16587_, _16418_);
  nand (_16589_, _16588_, _03839_);
  and (_16590_, _16589_, _08457_);
  and (_16591_, _16590_, _16586_);
  nor (_16593_, _08457_, _04034_);
  or (_16594_, _16593_, _08464_);
  or (_16595_, _16594_, _16591_);
  or (_16596_, _08469_, _08653_);
  and (_16597_, _16596_, _16260_);
  and (_16598_, _16597_, _16595_);
  and (_16599_, _16259_, _07975_);
  or (_16600_, _16599_, _16598_);
  and (_16601_, _16600_, _16078_);
  and (_16602_, _07975_, _04339_);
  or (_16604_, _16602_, _03957_);
  or (_16605_, _16604_, _16601_);
  or (_16606_, _10451_, _03958_);
  and (_16607_, _16606_, _08479_);
  and (_16608_, _16607_, _16605_);
  and (_16609_, _08478_, _08736_);
  or (_16610_, _16609_, _03838_);
  or (_16611_, _16610_, _16608_);
  and (_16612_, _16611_, _16421_);
  or (_16613_, _16612_, _03959_);
  or (_16615_, _16418_, _04701_);
  and (_16616_, _16615_, _15080_);
  and (_16617_, _16616_, _16613_);
  or (_16618_, _14948_, _08651_);
  and (_16619_, _16618_, _10611_);
  or (_16620_, _16619_, _16617_);
  or (_16621_, _14950_, _08651_);
  and (_16622_, _16621_, _08503_);
  and (_16623_, _16622_, _16620_);
  and (_16624_, _08502_, _07973_);
  or (_16626_, _16624_, _03965_);
  or (_16627_, _16626_, _16623_);
  or (_16628_, _08696_, _03966_);
  and (_16629_, _16628_, _16627_);
  or (_16630_, _16629_, _08508_);
  or (_16631_, _08509_, _08734_);
  and (_16632_, _16631_, _04708_);
  and (_16633_, _16632_, _16630_);
  or (_16634_, _16588_, _08697_);
  nor (_16635_, _16634_, _04708_);
  or (_16637_, _16635_, _16414_);
  or (_16638_, _16637_, _16633_);
  and (_16639_, _16638_, _16417_);
  nor (_16640_, _08652_, _16413_);
  or (_16641_, _16640_, _08521_);
  or (_16642_, _16641_, _16639_);
  nand (_16643_, _08521_, _07974_);
  and (_16644_, _16643_, _03953_);
  and (_16645_, _16644_, _16642_);
  nand (_16646_, _08529_, _08697_);
  and (_16648_, _16646_, _08528_);
  or (_16649_, _16648_, _16645_);
  nand (_16650_, _08526_, _08735_);
  and (_16651_, _16650_, _06532_);
  and (_16652_, _16651_, _16649_);
  nor (_16653_, _13131_, _08094_);
  nor (_16654_, _16653_, _16418_);
  nor (_16655_, _16654_, _06532_);
  or (_16656_, _16655_, _15379_);
  or (_16657_, _16656_, _16652_);
  and (_16659_, _16657_, _16412_);
  or (_16660_, _16659_, _08079_);
  and (_16661_, _08071_, _08029_);
  nor (_16662_, _16661_, _08072_);
  or (_16663_, _16662_, _08080_);
  and (_16664_, _16663_, _03964_);
  and (_16665_, _16664_, _16660_);
  and (_16666_, _08598_, _08313_);
  nor (_16667_, _16666_, _08599_);
  and (_16668_, _16667_, _03963_);
  or (_16670_, _16668_, _08580_);
  or (_16671_, _16670_, _16665_);
  and (_16672_, _08625_, _08380_);
  nor (_16673_, _16672_, _08626_);
  or (_16674_, _16673_, _08581_);
  and (_16675_, _16674_, _08007_);
  and (_16676_, _16675_, _16671_);
  nand (_16677_, _08006_, \oc8051_golden_model_1.ACC [4]);
  nand (_16678_, _16677_, _10007_);
  or (_16679_, _16678_, _16676_);
  and (_16681_, _16679_, _16409_);
  or (_16682_, _16681_, _07966_);
  and (_16683_, _07997_, _07976_);
  nor (_16684_, _16683_, _07998_);
  or (_16685_, _16684_, _10004_);
  and (_16686_, _16685_, _04166_);
  and (_16687_, _16686_, _16682_);
  nor (_16688_, _08720_, _10451_);
  and (_16689_, _08720_, _10451_);
  or (_16690_, _16689_, _16688_);
  or (_16692_, _16690_, _08691_);
  and (_16693_, _16692_, _09990_);
  or (_16694_, _16693_, _16687_);
  and (_16695_, _08759_, _08737_);
  nor (_16696_, _16695_, _08760_);
  or (_16697_, _16696_, _08692_);
  and (_16698_, _16697_, _10870_);
  and (_16699_, _16698_, _16694_);
  and (_16700_, _07964_, \oc8051_golden_model_1.ACC [4]);
  or (_16701_, _16700_, _03703_);
  or (_16703_, _16701_, _16699_);
  nand (_16704_, _16477_, _03703_);
  and (_16705_, _16704_, _08773_);
  and (_16706_, _16705_, _16703_);
  nor (_16707_, _16376_, _07634_);
  or (_16708_, _16707_, _08780_);
  and (_16709_, _16708_, _08772_);
  or (_16710_, _16709_, _08777_);
  or (_16711_, _16710_, _16706_);
  nand (_16712_, _08777_, _07586_);
  and (_16714_, _16712_, _03385_);
  and (_16715_, _16714_, _16711_);
  nor (_16716_, _16508_, _03385_);
  or (_16717_, _16716_, _03701_);
  or (_16718_, _16717_, _16715_);
  and (_16719_, _13193_, _05365_);
  nor (_16720_, _16719_, _16418_);
  nand (_16721_, _16720_, _03701_);
  and (_16722_, _16721_, _08795_);
  and (_16723_, _16722_, _16718_);
  nor (_16725_, _08804_, \oc8051_golden_model_1.ACC [5]);
  nor (_16726_, _16725_, _08805_);
  nor (_16727_, _16726_, _08801_);
  nor (_16728_, _16727_, _10917_);
  or (_16729_, _16728_, _16723_);
  nand (_16730_, _08801_, _07586_);
  and (_16731_, _16730_, _42908_);
  and (_16732_, _16731_, _16729_);
  or (_16733_, _16732_, _16406_);
  and (_43150_, _16733_, _41654_);
  nor (_16735_, _42908_, _07586_);
  nand (_16736_, _07964_, _07634_);
  nand (_16737_, _08649_, _08083_);
  not (_16738_, _04124_);
  and (_16739_, _04957_, _03476_);
  nor (_16740_, _16739_, _08085_);
  and (_16741_, _16740_, _16738_);
  not (_16742_, _16741_);
  and (_16743_, _16742_, _08648_);
  nor (_16744_, _05365_, _07586_);
  and (_16746_, _13341_, _05365_);
  nor (_16747_, _16746_, _16744_);
  nand (_16748_, _16747_, _03838_);
  or (_16749_, _07972_, _16078_);
  nand (_16750_, _03740_, _03466_);
  nor (_16751_, _06013_, _08094_);
  nor (_16752_, _16751_, _16744_);
  nand (_16753_, _16752_, _07544_);
  or (_16754_, _06941_, _07634_);
  and (_16755_, _06941_, _07634_);
  or (_16757_, _16523_, _16755_);
  and (_16758_, _16757_, _16754_);
  nor (_16759_, _16758_, _07972_);
  and (_16760_, _16758_, _07972_);
  nor (_16761_, _16760_, _16759_);
  nor (_16762_, _16533_, _16528_);
  and (_16763_, _16762_, \oc8051_golden_model_1.PSW [7]);
  nor (_16764_, _16763_, _16761_);
  and (_16765_, _16763_, _16761_);
  nor (_16766_, _16765_, _16764_);
  and (_16768_, _16766_, _08260_);
  nand (_16769_, _06013_, _04839_);
  nand (_16770_, _08105_, _06013_);
  nor (_16771_, _04234_, _07586_);
  and (_16772_, _04234_, _07586_);
  or (_16773_, _16772_, _16771_);
  or (_16774_, _16773_, _08105_);
  and (_16775_, _16774_, _08108_);
  and (_16776_, _16775_, _16770_);
  and (_16777_, _08107_, _06933_);
  or (_16779_, _16777_, _16776_);
  and (_16780_, _16779_, _08118_);
  nor (_16781_, _13234_, _08094_);
  nor (_16782_, _16781_, _16744_);
  nor (_16783_, _16782_, _04630_);
  or (_16784_, _16783_, _08120_);
  or (_16785_, _16784_, _16780_);
  not (_16786_, _08138_);
  nor (_16787_, _16483_, _16786_);
  and (_16788_, _11756_, _08139_);
  nor (_16790_, _16788_, _16787_);
  nand (_16791_, _16790_, _08120_);
  and (_16792_, _16791_, _03761_);
  and (_16793_, _16792_, _16785_);
  nor (_16794_, _06086_, _07586_);
  and (_16795_, _13238_, _06086_);
  nor (_16796_, _16795_, _16794_);
  nor (_16797_, _16796_, _03697_);
  nor (_16798_, _16752_, _04537_);
  or (_16799_, _16798_, _04839_);
  or (_16801_, _16799_, _16797_);
  or (_16802_, _16801_, _16793_);
  and (_16803_, _16802_, _16769_);
  or (_16804_, _16803_, _04645_);
  or (_16805_, _06933_, _04646_);
  and (_16806_, _16805_, _03751_);
  and (_16807_, _16806_, _16804_);
  nor (_16808_, _06015_, _03751_);
  or (_16809_, _16808_, _08098_);
  or (_16810_, _16809_, _16807_);
  nand (_16812_, _08098_, _07740_);
  and (_16813_, _16812_, _16810_);
  or (_16814_, _16813_, _03691_);
  and (_16815_, _13218_, _06086_);
  nor (_16816_, _16815_, _16794_);
  nand (_16817_, _16816_, _03691_);
  and (_16818_, _16817_, _03685_);
  and (_16819_, _16818_, _16814_);
  and (_16820_, _16795_, _13253_);
  nor (_16821_, _16820_, _16794_);
  nor (_16823_, _16821_, _03685_);
  or (_16824_, _16823_, _07024_);
  or (_16825_, _16824_, _16819_);
  nor (_16826_, _07499_, _07497_);
  nor (_16827_, _16826_, _07500_);
  or (_16828_, _16827_, _07030_);
  and (_16829_, _16828_, _16825_);
  or (_16830_, _16829_, _08182_);
  nand (_16831_, _05799_, \oc8051_golden_model_1.ACC [5]);
  nor (_16832_, _05799_, \oc8051_golden_model_1.ACC [5]);
  or (_16834_, _16443_, _16832_);
  and (_16835_, _16834_, _16831_);
  nor (_16836_, _16835_, _08650_);
  and (_16837_, _16835_, _08650_);
  nor (_16838_, _16837_, _16836_);
  nor (_16839_, _16453_, _16447_);
  and (_16840_, _16839_, \oc8051_golden_model_1.PSW [7]);
  nor (_16841_, _16840_, _16838_);
  and (_16842_, _16840_, _16838_);
  nor (_16843_, _16842_, _16841_);
  or (_16845_, _16843_, _08181_);
  and (_16846_, _16845_, _08261_);
  and (_16847_, _16846_, _16830_);
  or (_16848_, _16847_, _03818_);
  or (_16849_, _16848_, _16768_);
  or (_16850_, _16541_, _11683_);
  and (_16851_, _16850_, _11682_);
  nor (_16852_, _08695_, _16851_);
  and (_16853_, _08695_, _16851_);
  nor (_16854_, _16853_, _16852_);
  nor (_16856_, _16551_, _16545_);
  and (_16857_, _16856_, \oc8051_golden_model_1.PSW [7]);
  or (_16858_, _16857_, _16854_);
  nand (_16859_, _16857_, _16854_);
  and (_16860_, _16859_, _16858_);
  or (_16861_, _16860_, _03823_);
  and (_16862_, _16861_, _08288_);
  and (_16863_, _16862_, _16849_);
  or (_16864_, _16428_, _11714_);
  and (_16865_, _16864_, _11713_);
  nor (_16867_, _16865_, _08733_);
  and (_16868_, _16865_, _08733_);
  nor (_16869_, _16868_, _16867_);
  nor (_16870_, _16438_, _16432_);
  and (_16871_, _16870_, \oc8051_golden_model_1.PSW [7]);
  or (_16872_, _16871_, _16869_);
  nand (_16873_, _16871_, _16869_);
  and (_16874_, _16873_, _16872_);
  and (_16875_, _16874_, _08287_);
  or (_16876_, _16875_, _03547_);
  or (_16878_, _16876_, _16863_);
  nand (_16879_, _03740_, _03547_);
  and (_16880_, _16879_, _03680_);
  and (_16881_, _16880_, _16878_);
  nor (_16882_, _13220_, _08432_);
  nor (_16883_, _16882_, _16794_);
  nor (_16884_, _16883_, _03680_);
  or (_16885_, _16884_, _07544_);
  or (_16886_, _16885_, _16881_);
  and (_16887_, _16886_, _16753_);
  or (_16889_, _16887_, _04678_);
  and (_16890_, _06933_, _05365_);
  nor (_16891_, _16890_, _16744_);
  nand (_16892_, _16891_, _04678_);
  and (_16893_, _16892_, _03415_);
  and (_16894_, _16893_, _16889_);
  nor (_16895_, _13326_, _08094_);
  nor (_16896_, _16895_, _16744_);
  nor (_16897_, _16896_, _03415_);
  or (_16898_, _16897_, _07558_);
  or (_16900_, _16898_, _16894_);
  not (_16901_, _07587_);
  and (_16902_, _07591_, _16901_);
  or (_16903_, _16902_, _07565_);
  and (_16904_, _16903_, _16900_);
  or (_16905_, _16904_, _03466_);
  and (_16906_, _16905_, _16750_);
  or (_16907_, _16906_, _03839_);
  and (_16908_, _13333_, _05365_);
  nor (_16909_, _16908_, _16744_);
  nand (_16911_, _16909_, _03839_);
  and (_16912_, _16911_, _08457_);
  and (_16913_, _16912_, _16907_);
  nor (_16914_, _08457_, _03740_);
  or (_16915_, _16914_, _15616_);
  or (_16916_, _16915_, _16913_);
  not (_16917_, _15775_);
  and (_16918_, _15621_, _16917_);
  or (_16919_, _15622_, _08650_);
  and (_16920_, _16919_, _16918_);
  and (_16922_, _16920_, _16916_);
  not (_16923_, _08650_);
  nor (_16924_, _16918_, _16923_);
  or (_16925_, _16924_, _15774_);
  or (_16926_, _16925_, _16922_);
  or (_16927_, _08650_, _15939_);
  and (_16928_, _16927_, _16260_);
  and (_16929_, _16928_, _16926_);
  or (_16930_, _07972_, _03349_);
  and (_16931_, _16930_, _08471_);
  or (_16933_, _16931_, _16929_);
  and (_16934_, _16933_, _16749_);
  or (_16935_, _16934_, _03957_);
  or (_16936_, _08695_, _03958_);
  and (_16937_, _16936_, _08479_);
  and (_16938_, _16937_, _16935_);
  and (_16939_, _08478_, _08733_);
  or (_16940_, _16939_, _03838_);
  or (_16941_, _16940_, _16938_);
  and (_16942_, _16941_, _16748_);
  or (_16944_, _16942_, _03959_);
  nor (_16945_, _16744_, _04701_);
  nor (_16946_, _16945_, _04095_);
  and (_16947_, _16946_, _16944_);
  and (_16948_, _08648_, _04095_);
  or (_16949_, _16948_, _16947_);
  and (_16950_, _16949_, _16741_);
  or (_16951_, _16950_, _16743_);
  and (_16952_, _16951_, _08503_);
  and (_16953_, _08502_, _07970_);
  or (_16955_, _16953_, _03965_);
  or (_16956_, _16955_, _16952_);
  or (_16957_, _08693_, _03966_);
  and (_16958_, _16957_, _08509_);
  and (_16959_, _16958_, _16956_);
  and (_16960_, _08508_, _08731_);
  or (_16961_, _16960_, _16959_);
  and (_16962_, _16961_, _04708_);
  or (_16963_, _16909_, _08694_);
  nor (_16964_, _16963_, _04708_);
  or (_16966_, _16964_, _08083_);
  or (_16967_, _16966_, _16962_);
  and (_16968_, _16967_, _16737_);
  or (_16969_, _16968_, _08521_);
  nand (_16970_, _08521_, _07971_);
  and (_16971_, _16970_, _03953_);
  and (_16972_, _16971_, _16969_);
  nor (_16973_, _08694_, _03953_);
  or (_16974_, _16973_, _08526_);
  or (_16975_, _16974_, _16972_);
  nand (_16977_, _08526_, _08732_);
  and (_16978_, _16977_, _16975_);
  or (_16979_, _16978_, _03835_);
  nor (_16980_, _13340_, _08094_);
  nor (_16981_, _16980_, _16744_);
  nand (_16982_, _16981_, _03835_);
  and (_16983_, _16982_, _08547_);
  and (_16984_, _16983_, _16979_);
  nor (_16985_, _08566_, _08253_);
  nor (_16986_, _16985_, _08567_);
  and (_16988_, _16986_, _15379_);
  or (_16989_, _16988_, _08079_);
  or (_16990_, _16989_, _16984_);
  nor (_16991_, _08073_, _08021_);
  nor (_16992_, _16991_, _08074_);
  or (_16993_, _16992_, _08080_);
  and (_16994_, _16993_, _03964_);
  and (_16995_, _16994_, _16990_);
  nor (_16996_, _08600_, _08353_);
  nor (_16997_, _16996_, _08601_);
  and (_16999_, _16997_, _03963_);
  or (_17000_, _16999_, _16995_);
  and (_17001_, _17000_, _08581_);
  nor (_17002_, _08627_, _08420_);
  nor (_17003_, _17002_, _08628_);
  and (_17004_, _17003_, _08580_);
  or (_17005_, _17004_, _08006_);
  or (_17006_, _17005_, _17001_);
  nand (_17007_, _08006_, _07634_);
  and (_17008_, _17007_, _10007_);
  and (_17010_, _17008_, _17006_);
  nor (_17011_, _08677_, _08650_);
  nor (_17012_, _17011_, _08678_);
  and (_17013_, _17012_, _15145_);
  or (_17014_, _17013_, _07966_);
  or (_17015_, _17014_, _17010_);
  nor (_17016_, _07999_, _07972_);
  nor (_17017_, _17016_, _08000_);
  or (_17018_, _17017_, _10004_);
  and (_17019_, _17018_, _17015_);
  or (_17021_, _17019_, _03709_);
  nor (_17022_, _08722_, _08695_);
  nor (_17023_, _17022_, _08723_);
  or (_17024_, _17023_, _04166_);
  and (_17025_, _17024_, _08692_);
  and (_17026_, _17025_, _17021_);
  nor (_17027_, _08761_, _08733_);
  nor (_17028_, _17027_, _08762_);
  and (_17029_, _17028_, _08691_);
  or (_17030_, _17029_, _07964_);
  or (_17032_, _17030_, _17026_);
  and (_17033_, _17032_, _16736_);
  or (_17034_, _17033_, _03703_);
  nand (_17035_, _16782_, _03703_);
  and (_17036_, _17035_, _08773_);
  and (_17037_, _17036_, _17034_);
  nor (_17038_, _08780_, _07586_);
  or (_17039_, _17038_, _08781_);
  and (_17040_, _17039_, _08772_);
  or (_17041_, _17040_, _08777_);
  or (_17043_, _17041_, _17037_);
  nand (_17044_, _08777_, _06142_);
  and (_17045_, _17044_, _03385_);
  and (_17046_, _17045_, _17043_);
  nor (_17047_, _16816_, _03385_);
  or (_17048_, _17047_, _03701_);
  or (_17049_, _17048_, _17046_);
  nor (_17050_, _13399_, _08094_);
  nor (_17051_, _17050_, _16744_);
  nand (_17052_, _17051_, _03701_);
  and (_17054_, _17052_, _08795_);
  and (_17055_, _17054_, _17049_);
  nor (_17056_, _08805_, \oc8051_golden_model_1.ACC [6]);
  nor (_17057_, _17056_, _08806_);
  nor (_17058_, _17057_, _08801_);
  nor (_17059_, _17058_, _10917_);
  or (_17060_, _17059_, _17055_);
  nand (_17061_, _08801_, _06142_);
  and (_17062_, _17061_, _42908_);
  and (_17063_, _17062_, _17060_);
  or (_17065_, _17063_, _16735_);
  and (_43151_, _17065_, _41654_);
  not (_17066_, _04170_);
  not (_17067_, \oc8051_golden_model_1.SBUF [0]);
  nor (_17068_, _05396_, _17067_);
  nor (_17069_, _05652_, _08839_);
  nor (_17070_, _17069_, _17068_);
  and (_17071_, _17070_, _17066_);
  and (_17072_, _05396_, \oc8051_golden_model_1.ACC [0]);
  nor (_17073_, _17072_, _17068_);
  nor (_17075_, _17073_, _03751_);
  nor (_17076_, _17073_, _04616_);
  nor (_17077_, _04615_, _17067_);
  or (_17078_, _17077_, _17076_);
  and (_17079_, _17078_, _04630_);
  nor (_17080_, _17070_, _04630_);
  or (_17081_, _17080_, _17079_);
  and (_17082_, _17081_, _04537_);
  and (_17083_, _05396_, _04608_);
  nor (_17084_, _17083_, _17068_);
  nor (_17086_, _17084_, _04537_);
  nor (_17087_, _17086_, _17082_);
  nor (_17088_, _17087_, _03750_);
  or (_17089_, _17088_, _07544_);
  nor (_17090_, _17089_, _17075_);
  and (_17091_, _17084_, _07544_);
  nor (_17092_, _17091_, _17090_);
  nor (_17093_, _17092_, _04678_);
  and (_17094_, _06935_, _05396_);
  nor (_17095_, _17068_, _04679_);
  not (_17097_, _17095_);
  nor (_17098_, _17097_, _17094_);
  nor (_17099_, _17098_, _17093_);
  and (_17100_, _17099_, _03415_);
  nor (_17101_, _12119_, _08839_);
  nor (_17102_, _17101_, _17068_);
  nor (_17103_, _17102_, _03415_);
  or (_17104_, _17103_, _17100_);
  and (_17105_, _17104_, _04694_);
  and (_17106_, _05396_, _06428_);
  nor (_17108_, _17106_, _17068_);
  nor (_17109_, _17108_, _04694_);
  or (_17110_, _17109_, _17105_);
  and (_17111_, _17110_, _04703_);
  and (_17112_, _12133_, _05396_);
  nor (_17113_, _17112_, _17068_);
  nor (_17114_, _17113_, _04703_);
  or (_17115_, _17114_, _17111_);
  and (_17116_, _17115_, _04701_);
  nor (_17117_, _10458_, _08839_);
  nor (_17119_, _17117_, _17068_);
  and (_17120_, _17072_, _05652_);
  or (_17121_, _17120_, _04701_);
  nor (_17122_, _17121_, _17119_);
  nor (_17123_, _17122_, _17116_);
  nor (_17124_, _17123_, _03866_);
  and (_17125_, _12013_, _05396_);
  or (_17126_, _17125_, _17068_);
  and (_17127_, _17126_, _03866_);
  or (_17128_, _17127_, _17124_);
  and (_17130_, _17128_, _04706_);
  nor (_17131_, _17120_, _17068_);
  nor (_17132_, _17131_, _04706_);
  or (_17133_, _17132_, _17130_);
  and (_17134_, _17133_, _06532_);
  nor (_17135_, _12132_, _08839_);
  nor (_17136_, _17135_, _17068_);
  nor (_17137_, _17136_, _06532_);
  or (_17138_, _17137_, _17134_);
  and (_17139_, _17138_, _06537_);
  nor (_17141_, _17119_, _06537_);
  nor (_17142_, _17141_, _17066_);
  not (_17143_, _17142_);
  nor (_17144_, _17143_, _17139_);
  nor (_17145_, _17144_, _17071_);
  or (_17146_, _17145_, _42912_);
  or (_17147_, _42908_, \oc8051_golden_model_1.SBUF [0]);
  and (_17148_, _17147_, _41654_);
  and (_43152_, _17148_, _17146_);
  and (_17149_, _06934_, _05396_);
  and (_17151_, _08839_, \oc8051_golden_model_1.SBUF [1]);
  or (_17152_, _17151_, _04679_);
  or (_17153_, _17152_, _17149_);
  and (_17154_, _05396_, _04813_);
  or (_17155_, _17154_, _17151_);
  or (_17156_, _17155_, _06994_);
  or (_17157_, _05396_, \oc8051_golden_model_1.SBUF [1]);
  and (_17158_, _12225_, _05396_);
  not (_17159_, _17158_);
  and (_17160_, _17159_, _17157_);
  or (_17162_, _17160_, _04630_);
  and (_17163_, _05396_, \oc8051_golden_model_1.ACC [1]);
  or (_17164_, _17163_, _17151_);
  and (_17165_, _17164_, _04615_);
  and (_17166_, _04616_, \oc8051_golden_model_1.SBUF [1]);
  or (_17167_, _17166_, _03757_);
  or (_17168_, _17167_, _17165_);
  and (_17169_, _17168_, _04537_);
  and (_17170_, _17169_, _17162_);
  and (_17171_, _17155_, _03755_);
  or (_17172_, _17171_, _17170_);
  and (_17173_, _17172_, _03751_);
  and (_17174_, _17164_, _03750_);
  or (_17175_, _17174_, _07544_);
  or (_17176_, _17175_, _17173_);
  and (_17177_, _17176_, _17156_);
  or (_17178_, _17177_, _04678_);
  and (_17179_, _17178_, _03415_);
  and (_17180_, _17179_, _17153_);
  nand (_17181_, _12313_, _05396_);
  and (_17184_, _17157_, _07559_);
  and (_17185_, _17184_, _17181_);
  or (_17186_, _17185_, _17180_);
  and (_17187_, _17186_, _03840_);
  or (_17188_, _12207_, _08839_);
  and (_17189_, _17157_, _03838_);
  and (_17190_, _17189_, _17188_);
  nand (_17191_, _05396_, _04515_);
  and (_17192_, _17191_, _03839_);
  and (_17193_, _17192_, _17157_);
  or (_17194_, _17193_, _03959_);
  or (_17195_, _17194_, _17190_);
  or (_17196_, _17195_, _17187_);
  nor (_17197_, _08710_, _08839_);
  or (_17198_, _17197_, _17151_);
  nand (_17199_, _08709_, _05396_);
  and (_17200_, _17199_, _17198_);
  or (_17201_, _17200_, _04701_);
  and (_17202_, _17201_, _04708_);
  and (_17203_, _17202_, _17196_);
  or (_17206_, _12206_, _08839_);
  and (_17207_, _17157_, _03866_);
  and (_17208_, _17207_, _17206_);
  or (_17209_, _17208_, _03967_);
  or (_17210_, _17209_, _17203_);
  nor (_17211_, _17151_, _04706_);
  nand (_17212_, _17211_, _17199_);
  and (_17213_, _17212_, _06532_);
  and (_17214_, _17213_, _17210_);
  or (_17215_, _17191_, _05603_);
  and (_17217_, _17215_, _03835_);
  and (_17218_, _17217_, _17157_);
  or (_17219_, _17218_, _03954_);
  or (_17220_, _17219_, _17214_);
  or (_17221_, _17198_, _06537_);
  and (_17222_, _17221_, _17220_);
  or (_17223_, _17222_, _03703_);
  or (_17224_, _17160_, _03704_);
  and (_17225_, _17224_, _03702_);
  and (_17226_, _17225_, _17223_);
  or (_17228_, _17158_, _17151_);
  and (_17229_, _17228_, _03701_);
  or (_17230_, _17229_, _17226_);
  or (_17231_, _17230_, _42912_);
  or (_17232_, _42908_, \oc8051_golden_model_1.SBUF [1]);
  and (_17233_, _17232_, _41654_);
  and (_43155_, _17233_, _17231_);
  not (_17234_, \oc8051_golden_model_1.SBUF [2]);
  nor (_17235_, _05396_, _17234_);
  and (_17236_, _05396_, \oc8051_golden_model_1.ACC [2]);
  nor (_17238_, _17236_, _17235_);
  nor (_17239_, _17238_, _03751_);
  nor (_17240_, _17238_, _04616_);
  nor (_17241_, _04615_, _17234_);
  or (_17242_, _17241_, _17240_);
  and (_17243_, _17242_, _04630_);
  nor (_17244_, _12427_, _08839_);
  nor (_17245_, _17244_, _17235_);
  nor (_17246_, _17245_, _04630_);
  or (_17247_, _17246_, _17243_);
  and (_17249_, _17247_, _04537_);
  nor (_17250_, _08839_, _05236_);
  nor (_17251_, _17250_, _17235_);
  nor (_17252_, _17251_, _04537_);
  nor (_17253_, _17252_, _17249_);
  nor (_17254_, _17253_, _03750_);
  or (_17255_, _17254_, _07544_);
  nor (_17256_, _17255_, _17239_);
  and (_17257_, _17251_, _07544_);
  nor (_17258_, _17257_, _17256_);
  nor (_17260_, _17258_, _04678_);
  and (_17261_, _06938_, _05396_);
  nor (_17262_, _17235_, _04679_);
  not (_17263_, _17262_);
  nor (_17264_, _17263_, _17261_);
  nor (_17265_, _17264_, _07559_);
  not (_17266_, _17265_);
  nor (_17267_, _17266_, _17260_);
  nor (_17268_, _12523_, _08839_);
  nor (_17269_, _17268_, _17235_);
  nor (_17271_, _17269_, _03415_);
  or (_17272_, _17271_, _08854_);
  or (_17273_, _17272_, _17267_);
  and (_17274_, _12537_, _05396_);
  or (_17275_, _17235_, _04703_);
  nor (_17276_, _17275_, _17274_);
  and (_17277_, _05396_, _06457_);
  nor (_17278_, _17277_, _17235_);
  and (_17279_, _17278_, _03839_);
  or (_17280_, _17279_, _03959_);
  nor (_17282_, _17280_, _17276_);
  and (_17283_, _17282_, _17273_);
  and (_17284_, _08707_, _05396_);
  nor (_17285_, _17284_, _17235_);
  nor (_17286_, _17285_, _04701_);
  nor (_17287_, _17286_, _17283_);
  nor (_17288_, _17287_, _03866_);
  nor (_17289_, _17235_, _05700_);
  not (_17290_, _17289_);
  nor (_17291_, _17278_, _04708_);
  and (_17293_, _17291_, _17290_);
  nor (_17294_, _17293_, _17288_);
  nor (_17295_, _17294_, _03967_);
  nor (_17296_, _17238_, _04706_);
  and (_17297_, _17296_, _17290_);
  or (_17298_, _17297_, _17295_);
  and (_17299_, _17298_, _06532_);
  nor (_17300_, _12536_, _08839_);
  nor (_17301_, _17300_, _17235_);
  nor (_17302_, _17301_, _06532_);
  or (_17304_, _17302_, _17299_);
  and (_17305_, _17304_, _06537_);
  nor (_17306_, _08706_, _08839_);
  nor (_17307_, _17306_, _17235_);
  nor (_17308_, _17307_, _06537_);
  or (_17309_, _17308_, _03703_);
  nor (_17310_, _17309_, _17305_);
  and (_17311_, _17245_, _03703_);
  or (_17312_, _17311_, _03701_);
  nor (_17313_, _17312_, _17310_);
  and (_17315_, _12596_, _05396_);
  nor (_17316_, _17315_, _17235_);
  nor (_17317_, _17316_, _03702_);
  or (_17318_, _17317_, _17313_);
  or (_17319_, _17318_, _42912_);
  or (_17320_, _42908_, \oc8051_golden_model_1.SBUF [2]);
  and (_17321_, _17320_, _41654_);
  and (_43156_, _17321_, _17319_);
  not (_17322_, \oc8051_golden_model_1.SBUF [3]);
  nor (_17323_, _05396_, _17322_);
  and (_17325_, _06937_, _05396_);
  or (_17326_, _17325_, _17323_);
  and (_17327_, _17326_, _04678_);
  and (_17328_, _05396_, \oc8051_golden_model_1.ACC [3]);
  nor (_17329_, _17328_, _17323_);
  nor (_17330_, _17329_, _04616_);
  nor (_17331_, _04615_, _17322_);
  or (_17332_, _17331_, _17330_);
  and (_17333_, _17332_, _04630_);
  nor (_17334_, _12610_, _08839_);
  nor (_17336_, _17334_, _17323_);
  nor (_17337_, _17336_, _04630_);
  or (_17338_, _17337_, _17333_);
  and (_17339_, _17338_, _04537_);
  nor (_17340_, _08839_, _05050_);
  nor (_17341_, _17340_, _17323_);
  nor (_17342_, _17341_, _04537_);
  nor (_17343_, _17342_, _17339_);
  nor (_17344_, _17343_, _03750_);
  nor (_17345_, _17329_, _03751_);
  nor (_17347_, _17345_, _07544_);
  not (_17348_, _17347_);
  nor (_17349_, _17348_, _17344_);
  and (_17350_, _17341_, _07544_);
  or (_17351_, _17350_, _04678_);
  nor (_17352_, _17351_, _17349_);
  or (_17353_, _17352_, _17327_);
  and (_17354_, _17353_, _03415_);
  nor (_17355_, _12724_, _08839_);
  nor (_17356_, _17355_, _17323_);
  nor (_17358_, _17356_, _03415_);
  or (_17359_, _17358_, _08854_);
  or (_17360_, _17359_, _17354_);
  and (_17361_, _12738_, _05396_);
  or (_17362_, _17323_, _04703_);
  or (_17363_, _17362_, _17361_);
  and (_17364_, _05396_, _06415_);
  nor (_17365_, _17364_, _17323_);
  and (_17366_, _17365_, _03839_);
  nor (_17367_, _17366_, _03959_);
  and (_17369_, _17367_, _17363_);
  and (_17370_, _17369_, _17360_);
  and (_17371_, _10455_, _05396_);
  nor (_17372_, _17371_, _17323_);
  nor (_17373_, _17372_, _04701_);
  nor (_17374_, _17373_, _17370_);
  nor (_17375_, _17374_, _03866_);
  nor (_17376_, _17323_, _05554_);
  not (_17377_, _17376_);
  nor (_17378_, _17365_, _04708_);
  and (_17380_, _17378_, _17377_);
  nor (_17381_, _17380_, _17375_);
  nor (_17382_, _17381_, _03967_);
  nor (_17383_, _17329_, _04706_);
  and (_17384_, _17383_, _17377_);
  or (_17385_, _17384_, _17382_);
  and (_17386_, _17385_, _06532_);
  nor (_17387_, _12737_, _08839_);
  nor (_17388_, _17387_, _17323_);
  nor (_17389_, _17388_, _06532_);
  or (_17391_, _17389_, _17386_);
  and (_17392_, _17391_, _06537_);
  nor (_17393_, _08701_, _08839_);
  nor (_17394_, _17393_, _17323_);
  nor (_17395_, _17394_, _06537_);
  or (_17396_, _17395_, _03703_);
  nor (_17397_, _17396_, _17392_);
  and (_17398_, _17336_, _03703_);
  or (_17399_, _17398_, _03701_);
  nor (_17400_, _17399_, _17397_);
  and (_17402_, _12792_, _05396_);
  nor (_17403_, _17402_, _17323_);
  nor (_17404_, _17403_, _03702_);
  or (_17405_, _17404_, _17400_);
  or (_17406_, _17405_, _42912_);
  or (_17407_, _42908_, \oc8051_golden_model_1.SBUF [3]);
  and (_17408_, _17407_, _41654_);
  and (_43157_, _17408_, _17406_);
  not (_17409_, \oc8051_golden_model_1.SBUF [4]);
  nor (_17410_, _05396_, _17409_);
  and (_17412_, _06422_, _05396_);
  nor (_17413_, _17412_, _17410_);
  and (_17414_, _17413_, _03839_);
  and (_17415_, _05396_, \oc8051_golden_model_1.ACC [4]);
  nor (_17416_, _17415_, _17410_);
  nor (_17417_, _17416_, _03751_);
  nor (_17418_, _17416_, _04616_);
  nor (_17419_, _04615_, _17409_);
  or (_17420_, _17419_, _17418_);
  and (_17421_, _17420_, _04630_);
  nor (_17423_, _12828_, _08839_);
  nor (_17424_, _17423_, _17410_);
  nor (_17425_, _17424_, _04630_);
  or (_17426_, _17425_, _17421_);
  and (_17427_, _17426_, _04537_);
  nor (_17428_, _05898_, _08839_);
  nor (_17429_, _17428_, _17410_);
  nor (_17430_, _17429_, _04537_);
  nor (_17431_, _17430_, _17427_);
  nor (_17432_, _17431_, _03750_);
  or (_17434_, _17432_, _07544_);
  nor (_17435_, _17434_, _17417_);
  and (_17436_, _17429_, _07544_);
  nor (_17437_, _17436_, _17435_);
  nor (_17438_, _17437_, _04678_);
  and (_17439_, _06942_, _05396_);
  nor (_17440_, _17410_, _04679_);
  not (_17441_, _17440_);
  nor (_17442_, _17441_, _17439_);
  or (_17443_, _17442_, _07559_);
  nor (_17445_, _17443_, _17438_);
  nor (_17446_, _12919_, _08839_);
  nor (_17447_, _17446_, _17410_);
  nor (_17448_, _17447_, _03415_);
  or (_17449_, _17448_, _03839_);
  nor (_17450_, _17449_, _17445_);
  nor (_17451_, _17450_, _17414_);
  or (_17452_, _17451_, _03838_);
  and (_17453_, _12933_, _05396_);
  or (_17454_, _17410_, _04703_);
  nor (_17456_, _17454_, _17453_);
  nor (_17457_, _17456_, _03959_);
  and (_17458_, _17457_, _17452_);
  and (_17459_, _08700_, _05396_);
  nor (_17460_, _17459_, _17410_);
  nor (_17461_, _17460_, _04701_);
  nor (_17462_, _17461_, _17458_);
  nor (_17463_, _17462_, _03866_);
  nor (_17464_, _17410_, _08303_);
  not (_17465_, _17464_);
  nor (_17467_, _17413_, _04708_);
  and (_17468_, _17467_, _17465_);
  nor (_17469_, _17468_, _17463_);
  nor (_17470_, _17469_, _03967_);
  nor (_17471_, _17416_, _04706_);
  and (_17472_, _17471_, _17465_);
  or (_17473_, _17472_, _17470_);
  and (_17474_, _17473_, _06532_);
  nor (_17475_, _12931_, _08839_);
  nor (_17476_, _17475_, _17410_);
  nor (_17478_, _17476_, _06532_);
  or (_17479_, _17478_, _17474_);
  and (_17480_, _17479_, _06537_);
  nor (_17481_, _08699_, _08839_);
  nor (_17482_, _17481_, _17410_);
  nor (_17483_, _17482_, _06537_);
  or (_17484_, _17483_, _03703_);
  nor (_17485_, _17484_, _17480_);
  and (_17486_, _17424_, _03703_);
  or (_17487_, _17486_, _03701_);
  nor (_17489_, _17487_, _17485_);
  and (_17490_, _12991_, _05396_);
  nor (_17491_, _17490_, _17410_);
  nor (_17492_, _17491_, _03702_);
  or (_17493_, _17492_, _17489_);
  or (_17494_, _17493_, _42912_);
  or (_17495_, _42908_, \oc8051_golden_model_1.SBUF [4]);
  and (_17496_, _17495_, _41654_);
  and (_43158_, _17496_, _17494_);
  and (_17497_, _08839_, \oc8051_golden_model_1.SBUF [5]);
  nor (_17499_, _13025_, _08839_);
  or (_17500_, _17499_, _17497_);
  or (_17501_, _17500_, _04630_);
  and (_17502_, _05396_, \oc8051_golden_model_1.ACC [5]);
  or (_17503_, _17502_, _17497_);
  and (_17504_, _17503_, _04615_);
  and (_17505_, _04616_, \oc8051_golden_model_1.SBUF [5]);
  or (_17506_, _17505_, _03757_);
  or (_17507_, _17506_, _17504_);
  and (_17508_, _17507_, _04537_);
  and (_17510_, _17508_, _17501_);
  nor (_17511_, _05799_, _08839_);
  or (_17512_, _17511_, _17497_);
  and (_17513_, _17512_, _03755_);
  or (_17514_, _17513_, _17510_);
  and (_17515_, _17514_, _03751_);
  and (_17516_, _17503_, _03750_);
  or (_17517_, _17516_, _07544_);
  or (_17518_, _17517_, _17515_);
  or (_17519_, _17512_, _06994_);
  and (_17521_, _17519_, _17518_);
  or (_17522_, _17521_, _04678_);
  and (_17523_, _06941_, _05396_);
  or (_17524_, _17497_, _04679_);
  or (_17525_, _17524_, _17523_);
  and (_17526_, _17525_, _03415_);
  and (_17527_, _17526_, _17522_);
  nor (_17528_, _13118_, _08839_);
  or (_17529_, _17528_, _17497_);
  and (_17530_, _17529_, _07559_);
  or (_17532_, _17530_, _08854_);
  or (_17533_, _17532_, _17527_);
  and (_17534_, _13133_, _05396_);
  or (_17535_, _17497_, _04703_);
  or (_17536_, _17535_, _17534_);
  and (_17537_, _06371_, _05396_);
  or (_17538_, _17537_, _17497_);
  or (_17539_, _17538_, _04694_);
  and (_17540_, _17539_, _04701_);
  and (_17541_, _17540_, _17536_);
  and (_17543_, _17541_, _17533_);
  and (_17544_, _10451_, _05396_);
  or (_17545_, _17544_, _17497_);
  and (_17546_, _17545_, _03959_);
  or (_17547_, _17546_, _17543_);
  and (_17548_, _17547_, _04708_);
  or (_17549_, _17497_, _08302_);
  and (_17550_, _17538_, _03866_);
  and (_17551_, _17550_, _17549_);
  or (_17552_, _17551_, _17548_);
  and (_17554_, _17552_, _04706_);
  and (_17555_, _17503_, _03967_);
  and (_17556_, _17555_, _17549_);
  or (_17557_, _17556_, _03835_);
  or (_17558_, _17557_, _17554_);
  nor (_17559_, _13131_, _08839_);
  or (_17560_, _17497_, _06532_);
  or (_17561_, _17560_, _17559_);
  and (_17562_, _17561_, _06537_);
  and (_17563_, _17562_, _17558_);
  nor (_17565_, _08697_, _08839_);
  or (_17566_, _17565_, _17497_);
  and (_17567_, _17566_, _03954_);
  or (_17568_, _17567_, _17563_);
  and (_17569_, _17568_, _03704_);
  and (_17570_, _17500_, _03703_);
  or (_17571_, _17570_, _03701_);
  or (_17572_, _17571_, _17569_);
  and (_17573_, _13193_, _05396_);
  or (_17574_, _17573_, _17497_);
  or (_17576_, _17574_, _03702_);
  and (_17577_, _17576_, _17572_);
  or (_17578_, _17577_, _42912_);
  or (_17579_, _42908_, \oc8051_golden_model_1.SBUF [5]);
  and (_17580_, _17579_, _41654_);
  and (_43159_, _17580_, _17578_);
  not (_17581_, \oc8051_golden_model_1.SBUF [6]);
  nor (_17582_, _05396_, _17581_);
  and (_17583_, _13333_, _05396_);
  nor (_17584_, _17583_, _17582_);
  and (_17586_, _17584_, _03839_);
  and (_17587_, _05396_, \oc8051_golden_model_1.ACC [6]);
  nor (_17588_, _17587_, _17582_);
  nor (_17589_, _17588_, _03751_);
  nor (_17590_, _17588_, _04616_);
  nor (_17591_, _04615_, _17581_);
  or (_17592_, _17591_, _17590_);
  and (_17593_, _17592_, _04630_);
  nor (_17594_, _13234_, _08839_);
  nor (_17595_, _17594_, _17582_);
  nor (_17597_, _17595_, _04630_);
  or (_17598_, _17597_, _17593_);
  and (_17599_, _17598_, _04537_);
  nor (_17600_, _06013_, _08839_);
  nor (_17601_, _17600_, _17582_);
  nor (_17602_, _17601_, _04537_);
  nor (_17603_, _17602_, _17599_);
  nor (_17604_, _17603_, _03750_);
  or (_17605_, _17604_, _07544_);
  nor (_17606_, _17605_, _17589_);
  and (_17608_, _17601_, _07544_);
  nor (_17609_, _17608_, _17606_);
  nor (_17610_, _17609_, _04678_);
  and (_17611_, _06933_, _05396_);
  nor (_17612_, _17582_, _04679_);
  not (_17613_, _17612_);
  nor (_17614_, _17613_, _17611_);
  or (_17615_, _17614_, _07559_);
  nor (_17616_, _17615_, _17610_);
  nor (_17617_, _13326_, _08839_);
  nor (_17619_, _17617_, _17582_);
  nor (_17620_, _17619_, _03415_);
  or (_17621_, _17620_, _03839_);
  nor (_17622_, _17621_, _17616_);
  nor (_17623_, _17622_, _17586_);
  or (_17624_, _17623_, _03838_);
  and (_17625_, _13341_, _05396_);
  or (_17626_, _17582_, _04703_);
  nor (_17627_, _17626_, _17625_);
  nor (_17628_, _17627_, _03959_);
  and (_17630_, _17628_, _17624_);
  and (_17631_, _08695_, _05396_);
  nor (_17632_, _17631_, _17582_);
  nor (_17633_, _17632_, _04701_);
  nor (_17634_, _17633_, _17630_);
  nor (_17635_, _17634_, _03866_);
  nor (_17636_, _17582_, _08289_);
  not (_17637_, _17636_);
  nor (_17638_, _17584_, _04708_);
  and (_17639_, _17638_, _17637_);
  nor (_17641_, _17639_, _17635_);
  nor (_17642_, _17641_, _03967_);
  nor (_17643_, _17588_, _04706_);
  and (_17644_, _17643_, _17637_);
  or (_17645_, _17644_, _17642_);
  and (_17646_, _17645_, _06532_);
  nor (_17647_, _13340_, _08839_);
  nor (_17648_, _17647_, _17582_);
  nor (_17649_, _17648_, _06532_);
  or (_17650_, _17649_, _17646_);
  and (_17652_, _17650_, _06537_);
  nor (_17653_, _08694_, _08839_);
  nor (_17654_, _17653_, _17582_);
  nor (_17655_, _17654_, _06537_);
  or (_17656_, _17655_, _03703_);
  nor (_17657_, _17656_, _17652_);
  and (_17658_, _17595_, _03703_);
  or (_17659_, _17658_, _03701_);
  nor (_17660_, _17659_, _17657_);
  nor (_17661_, _13399_, _08839_);
  nor (_17663_, _17661_, _17582_);
  nor (_17664_, _17663_, _03702_);
  or (_17665_, _17664_, _17660_);
  or (_17666_, _17665_, _42912_);
  or (_17667_, _42908_, \oc8051_golden_model_1.SBUF [6]);
  and (_17668_, _17667_, _41654_);
  and (_43160_, _17668_, _17666_);
  not (_17669_, \oc8051_golden_model_1.SCON [0]);
  nor (_17670_, _05406_, _17669_);
  nor (_17671_, _05652_, _08924_);
  nor (_17673_, _17671_, _17670_);
  nor (_17674_, _17673_, _03702_);
  and (_17675_, _05406_, _06428_);
  nor (_17676_, _17675_, _17670_);
  and (_17677_, _17676_, _03839_);
  and (_17678_, _05406_, _04608_);
  nor (_17679_, _17678_, _17670_);
  and (_17680_, _17679_, _07544_);
  and (_17681_, _05406_, \oc8051_golden_model_1.ACC [0]);
  nor (_17682_, _17681_, _17670_);
  nor (_17684_, _17682_, _04616_);
  nor (_17685_, _04615_, _17669_);
  or (_17686_, _17685_, _17684_);
  and (_17687_, _17686_, _04630_);
  nor (_17688_, _17673_, _04630_);
  or (_17689_, _17688_, _17687_);
  and (_17690_, _17689_, _03697_);
  nor (_17691_, _06099_, _17669_);
  and (_17692_, _12032_, _06099_);
  nor (_17693_, _17692_, _17691_);
  nor (_17695_, _17693_, _03697_);
  nor (_17696_, _17695_, _17690_);
  nor (_17697_, _17696_, _03755_);
  nor (_17698_, _17679_, _04537_);
  or (_17699_, _17698_, _17697_);
  and (_17700_, _17699_, _03751_);
  nor (_17701_, _17682_, _03751_);
  or (_17702_, _17701_, _17700_);
  and (_17703_, _17702_, _03692_);
  and (_17704_, _17670_, _03691_);
  or (_17706_, _17704_, _17703_);
  and (_17707_, _17706_, _03685_);
  nor (_17708_, _17673_, _03685_);
  or (_17709_, _17708_, _17707_);
  and (_17710_, _17709_, _03680_);
  nor (_17711_, _17691_, _14175_);
  or (_17712_, _17711_, _03680_);
  nor (_17713_, _17712_, _17693_);
  nor (_17714_, _17713_, _07544_);
  not (_17715_, _17714_);
  nor (_17717_, _17715_, _17710_);
  nor (_17718_, _17717_, _17680_);
  nor (_17719_, _17718_, _04678_);
  and (_17720_, _06935_, _05406_);
  nor (_17721_, _17670_, _04679_);
  not (_17722_, _17721_);
  nor (_17723_, _17722_, _17720_);
  or (_17724_, _17723_, _07559_);
  nor (_17725_, _17724_, _17719_);
  nor (_17726_, _12119_, _08924_);
  nor (_17728_, _17726_, _17670_);
  nor (_17729_, _17728_, _03415_);
  or (_17730_, _17729_, _03839_);
  nor (_17731_, _17730_, _17725_);
  nor (_17732_, _17731_, _17677_);
  or (_17733_, _17732_, _03838_);
  and (_17734_, _12133_, _05406_);
  or (_17735_, _17670_, _04703_);
  nor (_17736_, _17735_, _17734_);
  nor (_17737_, _17736_, _03959_);
  and (_17739_, _17737_, _17733_);
  nor (_17740_, _10458_, _08924_);
  nor (_17741_, _17740_, _17670_);
  not (_17742_, _17741_);
  and (_17743_, _08712_, _05406_);
  nor (_17744_, _17743_, _04701_);
  and (_17745_, _17744_, _17742_);
  nor (_17746_, _17745_, _17739_);
  nor (_17747_, _17746_, _03866_);
  and (_17748_, _12013_, _05406_);
  or (_17750_, _17748_, _17670_);
  and (_17751_, _17750_, _03866_);
  or (_17752_, _17751_, _17747_);
  and (_17753_, _17752_, _04706_);
  nor (_17754_, _17743_, _17670_);
  nor (_17755_, _17754_, _04706_);
  or (_17756_, _17755_, _17753_);
  and (_17757_, _17756_, _06532_);
  nor (_17758_, _12132_, _08924_);
  nor (_17759_, _17758_, _17670_);
  nor (_17761_, _17759_, _06532_);
  or (_17762_, _17761_, _17757_);
  and (_17763_, _17762_, _06537_);
  nor (_17764_, _17741_, _06537_);
  or (_17765_, _17764_, _03703_);
  or (_17766_, _17765_, _17763_);
  nand (_17767_, _17673_, _03703_);
  and (_17768_, _17767_, _17766_);
  nor (_17769_, _17768_, _03384_);
  nor (_17770_, _17670_, _03385_);
  nor (_17772_, _17770_, _17769_);
  and (_17773_, _17772_, _03702_);
  nor (_17774_, _17773_, _17674_);
  nand (_17775_, _17774_, _42908_);
  or (_17776_, _42908_, \oc8051_golden_model_1.SCON [0]);
  and (_17777_, _17776_, _41654_);
  and (_43161_, _17777_, _17775_);
  not (_17778_, \oc8051_golden_model_1.SCON [1]);
  nor (_17779_, _05406_, _17778_);
  and (_17780_, _06934_, _05406_);
  or (_17782_, _17780_, _17779_);
  and (_17783_, _17782_, _04678_);
  and (_17784_, _05406_, \oc8051_golden_model_1.ACC [1]);
  nor (_17785_, _17784_, _17779_);
  nor (_17786_, _17785_, _04616_);
  nor (_17787_, _04615_, _17778_);
  or (_17788_, _17787_, _17786_);
  and (_17789_, _17788_, _04630_);
  nor (_17790_, _05406_, \oc8051_golden_model_1.SCON [1]);
  and (_17791_, _12225_, _05406_);
  nor (_17793_, _17791_, _17790_);
  and (_17794_, _17793_, _03757_);
  or (_17795_, _17794_, _17789_);
  and (_17796_, _17795_, _03697_);
  nor (_17797_, _06099_, _17778_);
  and (_17798_, _12212_, _06099_);
  nor (_17799_, _17798_, _17797_);
  nor (_17800_, _17799_, _03697_);
  or (_17801_, _17800_, _17796_);
  and (_17802_, _17801_, _04537_);
  and (_17804_, _05406_, _04813_);
  nor (_17805_, _17804_, _17779_);
  nor (_17806_, _17805_, _04537_);
  or (_17807_, _17806_, _17802_);
  and (_17808_, _17807_, _03751_);
  nor (_17809_, _17785_, _03751_);
  or (_17810_, _17809_, _17808_);
  and (_17811_, _17810_, _03692_);
  and (_17812_, _12200_, _06099_);
  nor (_17813_, _17812_, _17797_);
  nor (_17815_, _17813_, _03692_);
  or (_17816_, _17815_, _03684_);
  or (_17817_, _17816_, _17811_);
  and (_17818_, _17798_, _12211_);
  or (_17819_, _17797_, _03685_);
  or (_17820_, _17819_, _17818_);
  and (_17821_, _17820_, _17817_);
  and (_17822_, _17821_, _03680_);
  nor (_17823_, _12256_, _08945_);
  nor (_17824_, _17797_, _17823_);
  nor (_17826_, _17824_, _03680_);
  or (_17827_, _17826_, _07544_);
  nor (_17828_, _17827_, _17822_);
  and (_17829_, _17805_, _07544_);
  or (_17830_, _17829_, _04678_);
  nor (_17831_, _17830_, _17828_);
  or (_17832_, _17831_, _17783_);
  and (_17833_, _17832_, _03415_);
  nor (_17834_, _12313_, _08924_);
  nor (_17835_, _17834_, _17779_);
  nor (_17837_, _17835_, _03415_);
  nor (_17838_, _17837_, _17833_);
  nor (_17839_, _17838_, _08854_);
  nor (_17840_, _12207_, _08924_);
  or (_17841_, _17840_, _04703_);
  and (_17842_, _05406_, _04515_);
  or (_17843_, _17842_, _04694_);
  and (_17844_, _17843_, _17841_);
  nor (_17845_, _17844_, _17790_);
  or (_17846_, _17845_, _03959_);
  nor (_17848_, _17846_, _17839_);
  nor (_17849_, _08710_, _08924_);
  nor (_17850_, _17849_, _17779_);
  and (_17851_, _08709_, _05406_);
  nor (_17852_, _17851_, _17850_);
  nor (_17853_, _17852_, _04701_);
  nor (_17854_, _17853_, _03866_);
  not (_17855_, _17854_);
  nor (_17856_, _17855_, _17848_);
  and (_17857_, _12206_, _05406_);
  or (_17859_, _17857_, _17779_);
  and (_17860_, _17859_, _03866_);
  or (_17861_, _17860_, _17856_);
  and (_17862_, _17861_, _04706_);
  nor (_17863_, _17851_, _17779_);
  nor (_17864_, _17863_, _04706_);
  or (_17865_, _17864_, _17862_);
  and (_17866_, _17865_, _06532_);
  and (_17867_, _17842_, _05602_);
  or (_17868_, _17867_, _06532_);
  nor (_17870_, _17868_, _17790_);
  or (_17871_, _17870_, _17866_);
  and (_17872_, _17871_, _06537_);
  nor (_17873_, _17850_, _06537_);
  or (_17874_, _17873_, _17872_);
  and (_17875_, _17874_, _03704_);
  and (_17876_, _17793_, _03703_);
  or (_17877_, _17876_, _17875_);
  and (_17878_, _17877_, _03385_);
  nor (_17879_, _17813_, _03385_);
  or (_17881_, _17879_, _17878_);
  and (_17882_, _17881_, _03702_);
  nor (_17883_, _17791_, _17779_);
  nor (_17884_, _17883_, _03702_);
  or (_17885_, _17884_, _17882_);
  or (_17886_, _17885_, _42912_);
  or (_17887_, _42908_, \oc8051_golden_model_1.SCON [1]);
  and (_17888_, _17887_, _41654_);
  and (_43162_, _17888_, _17886_);
  not (_17889_, \oc8051_golden_model_1.SCON [2]);
  nor (_17891_, _05406_, _17889_);
  and (_17892_, _05406_, _06457_);
  nor (_17893_, _17892_, _17891_);
  and (_17894_, _17893_, _03839_);
  nor (_17895_, _08924_, _05236_);
  nor (_17896_, _17895_, _17891_);
  and (_17897_, _17896_, _07544_);
  and (_17898_, _05406_, \oc8051_golden_model_1.ACC [2]);
  nor (_17899_, _17898_, _17891_);
  nor (_17900_, _17899_, _04616_);
  nor (_17902_, _04615_, _17889_);
  or (_17903_, _17902_, _17900_);
  and (_17904_, _17903_, _04630_);
  nor (_17905_, _12427_, _08924_);
  nor (_17906_, _17905_, _17891_);
  nor (_17907_, _17906_, _04630_);
  or (_17908_, _17907_, _17904_);
  and (_17909_, _17908_, _03697_);
  nor (_17910_, _06099_, _17889_);
  and (_17911_, _12419_, _06099_);
  nor (_17913_, _17911_, _17910_);
  nor (_17914_, _17913_, _03697_);
  or (_17915_, _17914_, _17909_);
  and (_17916_, _17915_, _04537_);
  nor (_17917_, _17896_, _04537_);
  or (_17918_, _17917_, _17916_);
  and (_17919_, _17918_, _03751_);
  nor (_17920_, _17899_, _03751_);
  or (_17921_, _17920_, _17919_);
  and (_17922_, _17921_, _03692_);
  and (_17924_, _12422_, _06099_);
  nor (_17925_, _17924_, _17910_);
  nor (_17926_, _17925_, _03692_);
  or (_17927_, _17926_, _17922_);
  and (_17928_, _17927_, _03685_);
  and (_17929_, _17911_, _12418_);
  or (_17930_, _17929_, _17910_);
  and (_17931_, _17930_, _03684_);
  or (_17932_, _17931_, _17928_);
  and (_17933_, _17932_, _03680_);
  nor (_17935_, _12465_, _08945_);
  nor (_17936_, _17935_, _17910_);
  nor (_17937_, _17936_, _03680_);
  nor (_17938_, _17937_, _07544_);
  not (_17939_, _17938_);
  nor (_17940_, _17939_, _17933_);
  nor (_17941_, _17940_, _17897_);
  nor (_17942_, _17941_, _04678_);
  and (_17943_, _06938_, _05406_);
  nor (_17944_, _17891_, _04679_);
  not (_17946_, _17944_);
  nor (_17947_, _17946_, _17943_);
  or (_17948_, _17947_, _07559_);
  nor (_17949_, _17948_, _17942_);
  nor (_17950_, _12523_, _08924_);
  nor (_17951_, _17891_, _17950_);
  nor (_17952_, _17951_, _03415_);
  or (_17953_, _17952_, _03839_);
  nor (_17954_, _17953_, _17949_);
  nor (_17955_, _17954_, _17894_);
  or (_17957_, _17955_, _03838_);
  and (_17958_, _12537_, _05406_);
  or (_17959_, _17891_, _04703_);
  nor (_17960_, _17959_, _17958_);
  nor (_17961_, _17960_, _03959_);
  and (_17962_, _17961_, _17957_);
  and (_17963_, _08707_, _05406_);
  nor (_17964_, _17963_, _17891_);
  nor (_17965_, _17964_, _04701_);
  nor (_17966_, _17965_, _17962_);
  nor (_17968_, _17966_, _03866_);
  nor (_17969_, _17891_, _05700_);
  not (_17970_, _17969_);
  nor (_17971_, _17893_, _04708_);
  and (_17972_, _17971_, _17970_);
  nor (_17973_, _17972_, _17968_);
  nor (_17974_, _17973_, _03967_);
  nor (_17975_, _17899_, _04706_);
  and (_17976_, _17975_, _17970_);
  or (_17977_, _17976_, _17974_);
  and (_17979_, _17977_, _06532_);
  nor (_17980_, _12536_, _08924_);
  nor (_17981_, _17980_, _17891_);
  nor (_17982_, _17981_, _06532_);
  or (_17983_, _17982_, _17979_);
  and (_17984_, _17983_, _06537_);
  nor (_17985_, _08706_, _08924_);
  nor (_17986_, _17985_, _17891_);
  nor (_17987_, _17986_, _06537_);
  or (_17988_, _17987_, _17984_);
  and (_17990_, _17988_, _03704_);
  nor (_17991_, _17906_, _03704_);
  or (_17992_, _17991_, _17990_);
  and (_17993_, _17992_, _03385_);
  nor (_17994_, _17925_, _03385_);
  or (_17995_, _17994_, _17993_);
  and (_17996_, _17995_, _03702_);
  and (_17997_, _12596_, _05406_);
  nor (_17998_, _17997_, _17891_);
  nor (_17999_, _17998_, _03702_);
  or (_18001_, _17999_, _17996_);
  or (_18002_, _18001_, _42912_);
  or (_18003_, _42908_, \oc8051_golden_model_1.SCON [2]);
  and (_18004_, _18003_, _41654_);
  and (_43163_, _18004_, _18002_);
  and (_18005_, _08924_, \oc8051_golden_model_1.SCON [3]);
  nor (_18006_, _08924_, _05050_);
  or (_18007_, _18006_, _18005_);
  or (_18008_, _18007_, _06994_);
  nor (_18009_, _12610_, _08924_);
  or (_18011_, _18009_, _18005_);
  or (_18012_, _18011_, _04630_);
  and (_18013_, _05406_, \oc8051_golden_model_1.ACC [3]);
  or (_18014_, _18013_, _18005_);
  and (_18015_, _18014_, _04615_);
  and (_18016_, _04616_, \oc8051_golden_model_1.SCON [3]);
  or (_18017_, _18016_, _03757_);
  or (_18018_, _18017_, _18015_);
  and (_18019_, _18018_, _03697_);
  and (_18020_, _18019_, _18012_);
  and (_18022_, _08945_, \oc8051_golden_model_1.SCON [3]);
  and (_18023_, _12619_, _06099_);
  or (_18024_, _18023_, _18022_);
  and (_18025_, _18024_, _03696_);
  or (_18026_, _18025_, _03755_);
  or (_18027_, _18026_, _18020_);
  or (_18028_, _18007_, _04537_);
  and (_18029_, _18028_, _18027_);
  or (_18030_, _18029_, _03750_);
  or (_18031_, _18014_, _03751_);
  and (_18033_, _18031_, _03692_);
  and (_18034_, _18033_, _18030_);
  and (_18035_, _12622_, _06099_);
  or (_18036_, _18035_, _18022_);
  and (_18037_, _18036_, _03691_);
  or (_18038_, _18037_, _03684_);
  or (_18039_, _18038_, _18034_);
  or (_18040_, _18022_, _12618_);
  and (_18041_, _18040_, _18024_);
  or (_18042_, _18041_, _03685_);
  and (_18044_, _18042_, _03680_);
  and (_18045_, _18044_, _18039_);
  nor (_18046_, _12665_, _08945_);
  or (_18047_, _18046_, _18022_);
  and (_18048_, _18047_, _03679_);
  or (_18049_, _18048_, _07544_);
  or (_18050_, _18049_, _18045_);
  and (_18051_, _18050_, _18008_);
  or (_18052_, _18051_, _04678_);
  and (_18053_, _06937_, _05406_);
  or (_18055_, _18005_, _04679_);
  or (_18056_, _18055_, _18053_);
  and (_18057_, _18056_, _03415_);
  and (_18058_, _18057_, _18052_);
  nor (_18059_, _12724_, _08924_);
  or (_18060_, _18005_, _18059_);
  and (_18061_, _18060_, _07559_);
  or (_18062_, _18061_, _18058_);
  or (_18063_, _18062_, _08854_);
  and (_18064_, _12738_, _05406_);
  or (_18066_, _18005_, _04703_);
  or (_18067_, _18066_, _18064_);
  and (_18068_, _05406_, _06415_);
  or (_18069_, _18068_, _18005_);
  or (_18070_, _18069_, _04694_);
  and (_18071_, _18070_, _04701_);
  and (_18072_, _18071_, _18067_);
  and (_18073_, _18072_, _18063_);
  and (_18074_, _10455_, _05406_);
  or (_18075_, _18074_, _18005_);
  and (_18077_, _18075_, _03959_);
  or (_18078_, _18077_, _18073_);
  and (_18079_, _18078_, _04708_);
  or (_18080_, _18005_, _05554_);
  and (_18081_, _18069_, _03866_);
  and (_18082_, _18081_, _18080_);
  or (_18083_, _18082_, _18079_);
  and (_18084_, _18083_, _04706_);
  and (_18085_, _18014_, _03967_);
  and (_18086_, _18085_, _18080_);
  or (_18088_, _18086_, _03835_);
  or (_18089_, _18088_, _18084_);
  nor (_18090_, _12737_, _08924_);
  or (_18091_, _18005_, _06532_);
  or (_18092_, _18091_, _18090_);
  and (_18093_, _18092_, _06537_);
  and (_18094_, _18093_, _18089_);
  nor (_18095_, _08701_, _08924_);
  or (_18096_, _18095_, _18005_);
  and (_18097_, _18096_, _03954_);
  or (_18099_, _18097_, _03703_);
  or (_18100_, _18099_, _18094_);
  or (_18101_, _18011_, _03704_);
  and (_18102_, _18101_, _03385_);
  and (_18103_, _18102_, _18100_);
  and (_18104_, _18036_, _03384_);
  or (_18105_, _18104_, _03701_);
  or (_18106_, _18105_, _18103_);
  and (_18107_, _12792_, _05406_);
  or (_18108_, _18107_, _18005_);
  or (_18110_, _18108_, _03702_);
  and (_18111_, _18110_, _18106_);
  or (_18112_, _18111_, _42912_);
  or (_18113_, _42908_, \oc8051_golden_model_1.SCON [3]);
  and (_18114_, _18113_, _41654_);
  and (_43164_, _18114_, _18112_);
  and (_18115_, _08924_, \oc8051_golden_model_1.SCON [4]);
  nor (_18116_, _05898_, _08924_);
  or (_18117_, _18116_, _18115_);
  or (_18118_, _18117_, _06994_);
  and (_18120_, _08945_, \oc8051_golden_model_1.SCON [4]);
  and (_18121_, _12808_, _06099_);
  or (_18122_, _18121_, _18120_);
  and (_18123_, _18122_, _03691_);
  nor (_18124_, _12828_, _08924_);
  or (_18125_, _18124_, _18115_);
  or (_18126_, _18125_, _04630_);
  and (_18127_, _05406_, \oc8051_golden_model_1.ACC [4]);
  or (_18128_, _18127_, _18115_);
  and (_18129_, _18128_, _04615_);
  and (_18131_, _04616_, \oc8051_golden_model_1.SCON [4]);
  or (_18132_, _18131_, _03757_);
  or (_18133_, _18132_, _18129_);
  and (_18134_, _18133_, _03697_);
  and (_18135_, _18134_, _18126_);
  and (_18136_, _12832_, _06099_);
  or (_18137_, _18136_, _18120_);
  and (_18138_, _18137_, _03696_);
  or (_18139_, _18138_, _03755_);
  or (_18140_, _18139_, _18135_);
  or (_18142_, _18117_, _04537_);
  and (_18143_, _18142_, _18140_);
  or (_18144_, _18143_, _03750_);
  or (_18145_, _18128_, _03751_);
  and (_18146_, _18145_, _03692_);
  and (_18147_, _18146_, _18144_);
  or (_18148_, _18147_, _18123_);
  and (_18149_, _18148_, _03685_);
  and (_18150_, _12848_, _06099_);
  or (_18151_, _18150_, _18120_);
  and (_18153_, _18151_, _03684_);
  or (_18154_, _18153_, _18149_);
  and (_18155_, _18154_, _03680_);
  nor (_18156_, _12810_, _08945_);
  or (_18157_, _18156_, _18120_);
  and (_18158_, _18157_, _03679_);
  or (_18159_, _18158_, _07544_);
  or (_18160_, _18159_, _18155_);
  and (_18161_, _18160_, _18118_);
  or (_18162_, _18161_, _04678_);
  and (_18164_, _06942_, _05406_);
  or (_18165_, _18115_, _04679_);
  or (_18166_, _18165_, _18164_);
  and (_18167_, _18166_, _03415_);
  and (_18168_, _18167_, _18162_);
  nor (_18169_, _12919_, _08924_);
  or (_18170_, _18169_, _18115_);
  and (_18171_, _18170_, _07559_);
  or (_18172_, _18171_, _08854_);
  or (_18173_, _18172_, _18168_);
  and (_18175_, _12933_, _05406_);
  or (_18176_, _18115_, _04703_);
  or (_18177_, _18176_, _18175_);
  and (_18178_, _06422_, _05406_);
  or (_18179_, _18178_, _18115_);
  or (_18180_, _18179_, _04694_);
  and (_18181_, _18180_, _04701_);
  and (_18182_, _18181_, _18177_);
  and (_18183_, _18182_, _18173_);
  and (_18184_, _08700_, _05406_);
  or (_18186_, _18184_, _18115_);
  and (_18187_, _18186_, _03959_);
  or (_18188_, _18187_, _18183_);
  and (_18189_, _18188_, _04708_);
  or (_18190_, _18115_, _08303_);
  and (_18191_, _18179_, _03866_);
  and (_18192_, _18191_, _18190_);
  or (_18193_, _18192_, _18189_);
  and (_18194_, _18193_, _04706_);
  and (_18195_, _18128_, _03967_);
  and (_18197_, _18195_, _18190_);
  or (_18198_, _18197_, _03835_);
  or (_18199_, _18198_, _18194_);
  nor (_18200_, _12931_, _08924_);
  or (_18201_, _18115_, _06532_);
  or (_18202_, _18201_, _18200_);
  and (_18203_, _18202_, _06537_);
  and (_18204_, _18203_, _18199_);
  nor (_18205_, _08699_, _08924_);
  or (_18206_, _18205_, _18115_);
  and (_18208_, _18206_, _03954_);
  or (_18209_, _18208_, _03703_);
  or (_18210_, _18209_, _18204_);
  or (_18211_, _18125_, _03704_);
  and (_18212_, _18211_, _03385_);
  and (_18213_, _18212_, _18210_);
  and (_18214_, _18122_, _03384_);
  or (_18215_, _18214_, _03701_);
  or (_18216_, _18215_, _18213_);
  and (_18217_, _12991_, _05406_);
  or (_18219_, _18217_, _18115_);
  or (_18220_, _18219_, _03702_);
  and (_18221_, _18220_, _18216_);
  or (_18222_, _18221_, _42912_);
  or (_18223_, _42908_, \oc8051_golden_model_1.SCON [4]);
  and (_18224_, _18223_, _41654_);
  and (_43165_, _18224_, _18222_);
  and (_18225_, _08924_, \oc8051_golden_model_1.SCON [5]);
  nor (_18226_, _13025_, _08924_);
  or (_18227_, _18226_, _18225_);
  or (_18229_, _18227_, _04630_);
  and (_18230_, _05406_, \oc8051_golden_model_1.ACC [5]);
  or (_18231_, _18230_, _18225_);
  and (_18232_, _18231_, _04615_);
  and (_18233_, _04616_, \oc8051_golden_model_1.SCON [5]);
  or (_18234_, _18233_, _03757_);
  or (_18235_, _18234_, _18232_);
  and (_18236_, _18235_, _03697_);
  and (_18237_, _18236_, _18229_);
  and (_18238_, _08945_, \oc8051_golden_model_1.SCON [5]);
  and (_18240_, _13029_, _06099_);
  or (_18241_, _18240_, _18238_);
  and (_18242_, _18241_, _03696_);
  or (_18243_, _18242_, _03755_);
  or (_18244_, _18243_, _18237_);
  nor (_18245_, _05799_, _08924_);
  or (_18246_, _18245_, _18225_);
  or (_18247_, _18246_, _04537_);
  and (_18248_, _18247_, _18244_);
  or (_18249_, _18248_, _03750_);
  or (_18251_, _18231_, _03751_);
  and (_18252_, _18251_, _03692_);
  and (_18253_, _18252_, _18249_);
  and (_18254_, _13007_, _06099_);
  or (_18255_, _18254_, _18238_);
  and (_18256_, _18255_, _03691_);
  or (_18257_, _18256_, _03684_);
  or (_18258_, _18257_, _18253_);
  or (_18259_, _18238_, _13044_);
  and (_18260_, _18259_, _18241_);
  or (_18262_, _18260_, _03685_);
  and (_18263_, _18262_, _03680_);
  and (_18264_, _18263_, _18258_);
  nor (_18265_, _13009_, _08945_);
  or (_18266_, _18265_, _18238_);
  and (_18267_, _18266_, _03679_);
  or (_18268_, _18267_, _07544_);
  or (_18269_, _18268_, _18264_);
  or (_18270_, _18246_, _06994_);
  and (_18271_, _18270_, _18269_);
  or (_18273_, _18271_, _04678_);
  and (_18274_, _06941_, _05406_);
  or (_18275_, _18225_, _04679_);
  or (_18276_, _18275_, _18274_);
  and (_18277_, _18276_, _03415_);
  and (_18278_, _18277_, _18273_);
  nor (_18279_, _13118_, _08924_);
  or (_18280_, _18279_, _18225_);
  and (_18281_, _18280_, _07559_);
  or (_18282_, _18281_, _08854_);
  or (_18284_, _18282_, _18278_);
  and (_18285_, _13133_, _05406_);
  or (_18286_, _18225_, _04703_);
  or (_18287_, _18286_, _18285_);
  and (_18288_, _06371_, _05406_);
  or (_18289_, _18288_, _18225_);
  or (_18290_, _18289_, _04694_);
  and (_18291_, _18290_, _04701_);
  and (_18292_, _18291_, _18287_);
  and (_18293_, _18292_, _18284_);
  and (_18295_, _10451_, _05406_);
  or (_18296_, _18295_, _18225_);
  and (_18297_, _18296_, _03959_);
  or (_18298_, _18297_, _18293_);
  and (_18299_, _18298_, _04708_);
  or (_18300_, _18225_, _08302_);
  and (_18301_, _18289_, _03866_);
  and (_18302_, _18301_, _18300_);
  or (_18303_, _18302_, _18299_);
  and (_18304_, _18303_, _04706_);
  and (_18306_, _18231_, _03967_);
  and (_18307_, _18306_, _18300_);
  or (_18308_, _18307_, _03835_);
  or (_18309_, _18308_, _18304_);
  nor (_18310_, _13131_, _08924_);
  or (_18311_, _18225_, _06532_);
  or (_18312_, _18311_, _18310_);
  and (_18313_, _18312_, _06537_);
  and (_18314_, _18313_, _18309_);
  nor (_18315_, _08697_, _08924_);
  or (_18317_, _18315_, _18225_);
  and (_18318_, _18317_, _03954_);
  or (_18319_, _18318_, _03703_);
  or (_18320_, _18319_, _18314_);
  or (_18321_, _18227_, _03704_);
  and (_18322_, _18321_, _03385_);
  and (_18323_, _18322_, _18320_);
  and (_18324_, _18255_, _03384_);
  or (_18325_, _18324_, _03701_);
  or (_18326_, _18325_, _18323_);
  and (_18328_, _13193_, _05406_);
  or (_18329_, _18328_, _18225_);
  or (_18330_, _18329_, _03702_);
  and (_18331_, _18330_, _18326_);
  or (_18332_, _18331_, _42912_);
  or (_18333_, _42908_, \oc8051_golden_model_1.SCON [5]);
  and (_18334_, _18333_, _41654_);
  and (_43166_, _18334_, _18332_);
  and (_18335_, _08924_, \oc8051_golden_model_1.SCON [6]);
  nor (_18336_, _06013_, _08924_);
  or (_18338_, _18336_, _18335_);
  or (_18339_, _18338_, _06994_);
  and (_18340_, _08945_, \oc8051_golden_model_1.SCON [6]);
  and (_18341_, _13218_, _06099_);
  or (_18342_, _18341_, _18340_);
  and (_18343_, _18342_, _03691_);
  nor (_18344_, _13234_, _08924_);
  or (_18345_, _18344_, _18335_);
  or (_18346_, _18345_, _04630_);
  and (_18347_, _05406_, \oc8051_golden_model_1.ACC [6]);
  or (_18349_, _18347_, _18335_);
  and (_18350_, _18349_, _04615_);
  and (_18351_, _04616_, \oc8051_golden_model_1.SCON [6]);
  or (_18352_, _18351_, _03757_);
  or (_18353_, _18352_, _18350_);
  and (_18354_, _18353_, _03697_);
  and (_18355_, _18354_, _18346_);
  and (_18356_, _13238_, _06099_);
  or (_18357_, _18356_, _18340_);
  and (_18358_, _18357_, _03696_);
  or (_18360_, _18358_, _03755_);
  or (_18361_, _18360_, _18355_);
  or (_18362_, _18338_, _04537_);
  and (_18363_, _18362_, _18361_);
  or (_18364_, _18363_, _03750_);
  or (_18365_, _18349_, _03751_);
  and (_18366_, _18365_, _03692_);
  and (_18367_, _18366_, _18364_);
  or (_18368_, _18367_, _18343_);
  and (_18369_, _18368_, _03685_);
  and (_18371_, _13254_, _06099_);
  or (_18372_, _18371_, _18340_);
  and (_18373_, _18372_, _03684_);
  or (_18374_, _18373_, _18369_);
  and (_18375_, _18374_, _03680_);
  nor (_18376_, _13220_, _08945_);
  or (_18377_, _18376_, _18340_);
  and (_18378_, _18377_, _03679_);
  or (_18379_, _18378_, _07544_);
  or (_18380_, _18379_, _18375_);
  and (_18382_, _18380_, _18339_);
  or (_18383_, _18382_, _04678_);
  and (_18384_, _06933_, _05406_);
  or (_18385_, _18335_, _04679_);
  or (_18386_, _18385_, _18384_);
  and (_18387_, _18386_, _03415_);
  and (_18388_, _18387_, _18383_);
  nor (_18389_, _13326_, _08924_);
  or (_18390_, _18389_, _18335_);
  and (_18391_, _18390_, _07559_);
  or (_18393_, _18391_, _08854_);
  or (_18394_, _18393_, _18388_);
  and (_18395_, _13341_, _05406_);
  or (_18396_, _18335_, _04703_);
  or (_18397_, _18396_, _18395_);
  and (_18398_, _13333_, _05406_);
  or (_18399_, _18398_, _18335_);
  or (_18400_, _18399_, _04694_);
  and (_18401_, _18400_, _04701_);
  and (_18402_, _18401_, _18397_);
  and (_18404_, _18402_, _18394_);
  and (_18405_, _08695_, _05406_);
  or (_18406_, _18405_, _18335_);
  and (_18407_, _18406_, _03959_);
  or (_18408_, _18407_, _18404_);
  and (_18409_, _18408_, _04708_);
  or (_18410_, _18335_, _08289_);
  and (_18411_, _18399_, _03866_);
  and (_18412_, _18411_, _18410_);
  or (_18413_, _18412_, _18409_);
  and (_18415_, _18413_, _04706_);
  and (_18416_, _18349_, _03967_);
  and (_18417_, _18416_, _18410_);
  or (_18418_, _18417_, _03835_);
  or (_18419_, _18418_, _18415_);
  nor (_18420_, _13340_, _08924_);
  or (_18421_, _18335_, _06532_);
  or (_18422_, _18421_, _18420_);
  and (_18423_, _18422_, _06537_);
  and (_18424_, _18423_, _18419_);
  nor (_18426_, _08694_, _08924_);
  or (_18427_, _18426_, _18335_);
  and (_18428_, _18427_, _03954_);
  or (_18429_, _18428_, _03703_);
  or (_18430_, _18429_, _18424_);
  or (_18431_, _18345_, _03704_);
  and (_18432_, _18431_, _03385_);
  and (_18433_, _18432_, _18430_);
  and (_18434_, _18342_, _03384_);
  or (_18435_, _18434_, _03701_);
  or (_18437_, _18435_, _18433_);
  nor (_18438_, _13399_, _08924_);
  or (_18439_, _18438_, _18335_);
  or (_18440_, _18439_, _03702_);
  and (_18441_, _18440_, _18437_);
  or (_18442_, _18441_, _42912_);
  or (_18443_, _42908_, \oc8051_golden_model_1.SCON [6]);
  and (_18444_, _18443_, _41654_);
  and (_43167_, _18444_, _18442_);
  not (_18445_, \oc8051_golden_model_1.PCON [0]);
  nor (_18447_, _05391_, _18445_);
  nor (_18448_, _05652_, _09032_);
  nor (_18449_, _18448_, _18447_);
  and (_18450_, _18449_, _17066_);
  and (_18451_, _05391_, \oc8051_golden_model_1.ACC [0]);
  nor (_18452_, _18451_, _18447_);
  nor (_18453_, _18452_, _03751_);
  nor (_18454_, _18452_, _04616_);
  nor (_18455_, _04615_, _18445_);
  or (_18456_, _18455_, _18454_);
  and (_18458_, _18456_, _04630_);
  nor (_18459_, _18449_, _04630_);
  or (_18460_, _18459_, _18458_);
  and (_18461_, _18460_, _04537_);
  and (_18462_, _05391_, _04608_);
  nor (_18463_, _18462_, _18447_);
  nor (_18464_, _18463_, _04537_);
  nor (_18465_, _18464_, _18461_);
  nor (_18466_, _18465_, _03750_);
  or (_18467_, _18466_, _07544_);
  nor (_18469_, _18467_, _18453_);
  and (_18470_, _18463_, _07544_);
  nor (_18471_, _18470_, _18469_);
  nor (_18472_, _18471_, _04678_);
  and (_18473_, _06935_, _05391_);
  nor (_18474_, _18447_, _04679_);
  not (_18475_, _18474_);
  nor (_18476_, _18475_, _18473_);
  nor (_18477_, _18476_, _18472_);
  and (_18478_, _18477_, _03415_);
  nor (_18480_, _12119_, _09032_);
  nor (_18481_, _18480_, _18447_);
  nor (_18482_, _18481_, _03415_);
  or (_18483_, _18482_, _18478_);
  and (_18484_, _18483_, _04694_);
  and (_18485_, _05391_, _06428_);
  nor (_18486_, _18485_, _18447_);
  nor (_18487_, _18486_, _04694_);
  or (_18488_, _18487_, _03838_);
  nor (_18489_, _18488_, _18484_);
  and (_18491_, _12133_, _05391_);
  or (_18492_, _18447_, _04703_);
  nor (_18493_, _18492_, _18491_);
  or (_18494_, _18493_, _03959_);
  nor (_18495_, _18494_, _18489_);
  nor (_18496_, _10458_, _09032_);
  nor (_18497_, _18496_, _18447_);
  not (_18498_, _18497_);
  and (_18499_, _08712_, _05391_);
  nor (_18500_, _18499_, _04701_);
  and (_18502_, _18500_, _18498_);
  nor (_18503_, _18502_, _18495_);
  nor (_18504_, _18503_, _03866_);
  and (_18505_, _12013_, _05391_);
  or (_18506_, _18505_, _18447_);
  and (_18507_, _18506_, _03866_);
  or (_18508_, _18507_, _18504_);
  and (_18509_, _18508_, _04706_);
  nor (_18510_, _18499_, _18447_);
  nor (_18511_, _18510_, _04706_);
  or (_18513_, _18511_, _18509_);
  and (_18514_, _18513_, _06532_);
  nor (_18515_, _12132_, _09032_);
  nor (_18516_, _18515_, _18447_);
  nor (_18517_, _18516_, _06532_);
  or (_18518_, _18517_, _18514_);
  and (_18519_, _18518_, _06537_);
  nor (_18520_, _18497_, _06537_);
  nor (_18521_, _18520_, _17066_);
  not (_18522_, _18521_);
  nor (_18524_, _18522_, _18519_);
  nor (_18525_, _18524_, _18450_);
  or (_18526_, _18525_, _42912_);
  or (_18527_, _42908_, \oc8051_golden_model_1.PCON [0]);
  and (_18528_, _18527_, _41654_);
  and (_43170_, _18528_, _18526_);
  and (_18529_, _06934_, _05391_);
  not (_18530_, \oc8051_golden_model_1.PCON [1]);
  nor (_18531_, _05391_, _18530_);
  nor (_18532_, _18531_, _04679_);
  not (_18534_, _18532_);
  nor (_18535_, _18534_, _18529_);
  not (_18536_, _18535_);
  and (_18537_, _05391_, \oc8051_golden_model_1.ACC [1]);
  nor (_18538_, _18537_, _18531_);
  nor (_18539_, _18538_, _03751_);
  nor (_18540_, _18538_, _04616_);
  nor (_18541_, _04615_, _18530_);
  or (_18542_, _18541_, _18540_);
  and (_18543_, _18542_, _04630_);
  nor (_18545_, _05391_, \oc8051_golden_model_1.PCON [1]);
  and (_18546_, _12225_, _05391_);
  nor (_18547_, _18546_, _18545_);
  and (_18548_, _18547_, _03757_);
  or (_18549_, _18548_, _18543_);
  and (_18550_, _18549_, _04537_);
  and (_18551_, _05391_, _04813_);
  nor (_18552_, _18551_, _18531_);
  nor (_18553_, _18552_, _04537_);
  nor (_18554_, _18553_, _18550_);
  nor (_18556_, _18554_, _03750_);
  or (_18557_, _18556_, _07544_);
  nor (_18558_, _18557_, _18539_);
  and (_18559_, _18552_, _07544_);
  nor (_18560_, _18559_, _18558_);
  nor (_18561_, _18560_, _04678_);
  nor (_18562_, _18561_, _07559_);
  and (_18563_, _18562_, _18536_);
  and (_18564_, _12313_, _05391_);
  or (_18565_, _18564_, _03415_);
  nor (_18567_, _18565_, _18545_);
  nor (_18568_, _18567_, _18563_);
  nor (_18569_, _18568_, _08854_);
  nor (_18570_, _12207_, _09032_);
  or (_18571_, _18570_, _04703_);
  and (_18572_, _05391_, _04515_);
  or (_18573_, _18572_, _04694_);
  and (_18574_, _18573_, _18571_);
  nor (_18575_, _18574_, _18545_);
  or (_18576_, _18575_, _03959_);
  nor (_18578_, _18576_, _18569_);
  nor (_18579_, _08710_, _09032_);
  nor (_18580_, _18579_, _18531_);
  and (_18581_, _08709_, _05391_);
  nor (_18582_, _18581_, _18580_);
  nor (_18583_, _18582_, _04701_);
  nor (_18584_, _18583_, _03866_);
  not (_18585_, _18584_);
  nor (_18586_, _18585_, _18578_);
  and (_18587_, _12206_, _05391_);
  or (_18589_, _18587_, _18531_);
  and (_18590_, _18589_, _03866_);
  or (_18591_, _18590_, _18586_);
  and (_18592_, _18591_, _04706_);
  nor (_18593_, _18581_, _18531_);
  nor (_18594_, _18593_, _04706_);
  or (_18595_, _18594_, _18592_);
  and (_18596_, _18595_, _06532_);
  and (_18597_, _18572_, _05602_);
  or (_18598_, _18597_, _06532_);
  nor (_18600_, _18598_, _18545_);
  or (_18601_, _18600_, _18596_);
  and (_18602_, _18601_, _06537_);
  nor (_18603_, _18580_, _06537_);
  or (_18604_, _18603_, _18602_);
  and (_18605_, _18604_, _03704_);
  and (_18606_, _18547_, _03703_);
  or (_18607_, _18606_, _18605_);
  and (_18608_, _18607_, _03702_);
  nor (_18609_, _18546_, _18531_);
  nor (_18611_, _18609_, _03702_);
  nor (_18612_, _18611_, _18608_);
  nand (_18613_, _18612_, _42908_);
  or (_18614_, _42908_, \oc8051_golden_model_1.PCON [1]);
  and (_18615_, _18614_, _41654_);
  and (_43171_, _18615_, _18613_);
  not (_18616_, \oc8051_golden_model_1.PCON [2]);
  nor (_18617_, _05391_, _18616_);
  and (_18618_, _05391_, \oc8051_golden_model_1.ACC [2]);
  nor (_18619_, _18618_, _18617_);
  nor (_18621_, _18619_, _03751_);
  nor (_18622_, _18619_, _04616_);
  nor (_18623_, _04615_, _18616_);
  or (_18624_, _18623_, _18622_);
  and (_18625_, _18624_, _04630_);
  nor (_18626_, _12427_, _09032_);
  nor (_18627_, _18626_, _18617_);
  nor (_18628_, _18627_, _04630_);
  or (_18629_, _18628_, _18625_);
  and (_18630_, _18629_, _04537_);
  nor (_18632_, _09032_, _05236_);
  nor (_18633_, _18632_, _18617_);
  nor (_18634_, _18633_, _04537_);
  nor (_18635_, _18634_, _18630_);
  nor (_18636_, _18635_, _03750_);
  or (_18637_, _18636_, _07544_);
  nor (_18638_, _18637_, _18621_);
  and (_18639_, _18633_, _07544_);
  nor (_18640_, _18639_, _18638_);
  nor (_18641_, _18640_, _04678_);
  and (_18643_, _06938_, _05391_);
  nor (_18644_, _18617_, _04679_);
  not (_18645_, _18644_);
  nor (_18646_, _18645_, _18643_);
  nor (_18647_, _18646_, _07559_);
  not (_18648_, _18647_);
  nor (_18649_, _18648_, _18641_);
  nor (_18650_, _12523_, _09032_);
  nor (_18651_, _18650_, _18617_);
  nor (_18652_, _18651_, _03415_);
  or (_18654_, _18652_, _08854_);
  or (_18655_, _18654_, _18649_);
  and (_18656_, _12537_, _05391_);
  or (_18657_, _18617_, _04703_);
  nor (_18658_, _18657_, _18656_);
  and (_18659_, _05391_, _06457_);
  nor (_18660_, _18659_, _18617_);
  and (_18661_, _18660_, _03839_);
  or (_18662_, _18661_, _03959_);
  nor (_18663_, _18662_, _18658_);
  and (_18665_, _18663_, _18655_);
  and (_18666_, _08707_, _05391_);
  nor (_18667_, _18666_, _18617_);
  nor (_18668_, _18667_, _04701_);
  nor (_18669_, _18668_, _18665_);
  nor (_18670_, _18669_, _03866_);
  nor (_18671_, _18617_, _05700_);
  not (_18672_, _18671_);
  nor (_18673_, _18660_, _04708_);
  and (_18674_, _18673_, _18672_);
  nor (_18676_, _18674_, _18670_);
  nor (_18677_, _18676_, _03967_);
  nor (_18678_, _18619_, _04706_);
  and (_18679_, _18678_, _18672_);
  or (_18680_, _18679_, _18677_);
  and (_18681_, _18680_, _06532_);
  nor (_18682_, _12536_, _09032_);
  nor (_18683_, _18682_, _18617_);
  nor (_18684_, _18683_, _06532_);
  or (_18685_, _18684_, _18681_);
  and (_18687_, _18685_, _06537_);
  nor (_18688_, _08706_, _09032_);
  nor (_18689_, _18688_, _18617_);
  nor (_18690_, _18689_, _06537_);
  or (_18691_, _18690_, _03703_);
  nor (_18692_, _18691_, _18687_);
  and (_18693_, _18627_, _03703_);
  or (_18694_, _18693_, _03701_);
  nor (_18695_, _18694_, _18692_);
  and (_18696_, _12596_, _05391_);
  nor (_18698_, _18696_, _18617_);
  nor (_18699_, _18698_, _03702_);
  or (_18700_, _18699_, _18695_);
  or (_18701_, _18700_, _42912_);
  or (_18702_, _42908_, \oc8051_golden_model_1.PCON [2]);
  and (_18703_, _18702_, _41654_);
  and (_43172_, _18703_, _18701_);
  and (_18704_, _09032_, \oc8051_golden_model_1.PCON [3]);
  nor (_18705_, _12610_, _09032_);
  or (_18706_, _18705_, _18704_);
  or (_18708_, _18706_, _04630_);
  and (_18709_, _05391_, \oc8051_golden_model_1.ACC [3]);
  or (_18710_, _18709_, _18704_);
  and (_18711_, _18710_, _04615_);
  and (_18712_, _04616_, \oc8051_golden_model_1.PCON [3]);
  or (_18713_, _18712_, _03757_);
  or (_18714_, _18713_, _18711_);
  and (_18715_, _18714_, _04537_);
  and (_18716_, _18715_, _18708_);
  nor (_18717_, _09032_, _05050_);
  or (_18719_, _18717_, _18704_);
  and (_18720_, _18719_, _03755_);
  or (_18721_, _18720_, _18716_);
  and (_18722_, _18721_, _03751_);
  and (_18723_, _18710_, _03750_);
  or (_18724_, _18723_, _07544_);
  or (_18725_, _18724_, _18722_);
  or (_18726_, _18719_, _06994_);
  and (_18727_, _18726_, _18725_);
  or (_18728_, _18727_, _04678_);
  and (_18730_, _06937_, _05391_);
  or (_18731_, _18704_, _04679_);
  or (_18732_, _18731_, _18730_);
  and (_18733_, _18732_, _03415_);
  and (_18734_, _18733_, _18728_);
  nor (_18735_, _12724_, _09032_);
  or (_18736_, _18735_, _18704_);
  and (_18737_, _18736_, _07559_);
  or (_18738_, _18737_, _08854_);
  or (_18739_, _18738_, _18734_);
  and (_18741_, _12738_, _05391_);
  or (_18742_, _18704_, _04703_);
  or (_18743_, _18742_, _18741_);
  and (_18744_, _05391_, _06415_);
  or (_18745_, _18744_, _18704_);
  or (_18746_, _18745_, _04694_);
  and (_18747_, _18746_, _04701_);
  and (_18748_, _18747_, _18743_);
  and (_18749_, _18748_, _18739_);
  and (_18750_, _10455_, _05391_);
  or (_18752_, _18750_, _18704_);
  and (_18753_, _18752_, _03959_);
  or (_18754_, _18753_, _18749_);
  and (_18755_, _18754_, _04708_);
  or (_18756_, _18704_, _05554_);
  and (_18757_, _18745_, _03866_);
  and (_18758_, _18757_, _18756_);
  or (_18759_, _18758_, _18755_);
  and (_18760_, _18759_, _04706_);
  and (_18761_, _18710_, _03967_);
  and (_18763_, _18761_, _18756_);
  or (_18764_, _18763_, _03835_);
  or (_18765_, _18764_, _18760_);
  nor (_18766_, _12737_, _09032_);
  or (_18767_, _18704_, _06532_);
  or (_18768_, _18767_, _18766_);
  and (_18769_, _18768_, _06537_);
  and (_18770_, _18769_, _18765_);
  nor (_18771_, _08701_, _09032_);
  or (_18772_, _18771_, _18704_);
  and (_18774_, _18772_, _03954_);
  or (_18775_, _18774_, _03703_);
  or (_18776_, _18775_, _18770_);
  or (_18777_, _18706_, _03704_);
  and (_18778_, _18777_, _03702_);
  and (_18779_, _18778_, _18776_);
  and (_18780_, _12792_, _05391_);
  or (_18781_, _18780_, _18704_);
  and (_18782_, _18781_, _03701_);
  or (_18783_, _18782_, _18779_);
  or (_18785_, _18783_, _42912_);
  or (_18786_, _42908_, \oc8051_golden_model_1.PCON [3]);
  and (_18787_, _18786_, _41654_);
  and (_43175_, _18787_, _18785_);
  not (_18788_, \oc8051_golden_model_1.PCON [4]);
  nor (_18789_, _05391_, _18788_);
  and (_18790_, _06422_, _05391_);
  nor (_18791_, _18790_, _18789_);
  and (_18792_, _18791_, _03839_);
  nor (_18793_, _05898_, _09032_);
  nor (_18795_, _18793_, _18789_);
  and (_18796_, _18795_, _07544_);
  and (_18797_, _05391_, \oc8051_golden_model_1.ACC [4]);
  nor (_18798_, _18797_, _18789_);
  nor (_18799_, _18798_, _04616_);
  nor (_18800_, _04615_, _18788_);
  or (_18801_, _18800_, _18799_);
  and (_18802_, _18801_, _04630_);
  nor (_18803_, _12828_, _09032_);
  nor (_18804_, _18803_, _18789_);
  nor (_18806_, _18804_, _04630_);
  or (_18807_, _18806_, _18802_);
  and (_18808_, _18807_, _04537_);
  nor (_18809_, _18795_, _04537_);
  nor (_18810_, _18809_, _18808_);
  nor (_18811_, _18810_, _03750_);
  nor (_18812_, _18798_, _03751_);
  nor (_18813_, _18812_, _07544_);
  not (_18814_, _18813_);
  nor (_18815_, _18814_, _18811_);
  nor (_18817_, _18815_, _18796_);
  nor (_18818_, _18817_, _04678_);
  and (_18819_, _06942_, _05391_);
  nor (_18820_, _18789_, _04679_);
  not (_18821_, _18820_);
  nor (_18822_, _18821_, _18819_);
  or (_18823_, _18822_, _07559_);
  nor (_18824_, _18823_, _18818_);
  nor (_18825_, _12919_, _09032_);
  nor (_18826_, _18825_, _18789_);
  nor (_18828_, _18826_, _03415_);
  or (_18829_, _18828_, _03839_);
  nor (_18830_, _18829_, _18824_);
  nor (_18831_, _18830_, _18792_);
  or (_18832_, _18831_, _03838_);
  and (_18833_, _12933_, _05391_);
  or (_18834_, _18833_, _18789_);
  or (_18835_, _18834_, _04703_);
  and (_18836_, _18835_, _04701_);
  and (_18837_, _18836_, _18832_);
  and (_18839_, _08700_, _05391_);
  nor (_18840_, _18839_, _18789_);
  nor (_18841_, _18840_, _04701_);
  nor (_18842_, _18841_, _18837_);
  nor (_18843_, _18842_, _03866_);
  nor (_18844_, _18789_, _08303_);
  not (_18845_, _18844_);
  nor (_18846_, _18791_, _04708_);
  and (_18847_, _18846_, _18845_);
  nor (_18848_, _18847_, _18843_);
  nor (_18850_, _18848_, _03967_);
  nor (_18851_, _18798_, _04706_);
  and (_18852_, _18851_, _18845_);
  or (_18853_, _18852_, _18850_);
  and (_18854_, _18853_, _06532_);
  nor (_18855_, _12931_, _09032_);
  nor (_18856_, _18855_, _18789_);
  nor (_18857_, _18856_, _06532_);
  or (_18858_, _18857_, _18854_);
  and (_18859_, _18858_, _06537_);
  nor (_18861_, _08699_, _09032_);
  nor (_18862_, _18861_, _18789_);
  nor (_18863_, _18862_, _06537_);
  or (_18864_, _18863_, _03703_);
  nor (_18865_, _18864_, _18859_);
  and (_18866_, _18804_, _03703_);
  or (_18867_, _18866_, _03701_);
  nor (_18868_, _18867_, _18865_);
  and (_18869_, _12991_, _05391_);
  nor (_18870_, _18869_, _18789_);
  nor (_18872_, _18870_, _03702_);
  or (_18873_, _18872_, _18868_);
  or (_18874_, _18873_, _42912_);
  or (_18875_, _42908_, \oc8051_golden_model_1.PCON [4]);
  and (_18876_, _18875_, _41654_);
  and (_43176_, _18876_, _18874_);
  and (_18877_, _09032_, \oc8051_golden_model_1.PCON [5]);
  nor (_18878_, _13025_, _09032_);
  or (_18879_, _18878_, _18877_);
  or (_18880_, _18879_, _04630_);
  and (_18882_, _05391_, \oc8051_golden_model_1.ACC [5]);
  or (_18883_, _18882_, _18877_);
  and (_18884_, _18883_, _04615_);
  and (_18885_, _04616_, \oc8051_golden_model_1.PCON [5]);
  or (_18886_, _18885_, _03757_);
  or (_18887_, _18886_, _18884_);
  and (_18888_, _18887_, _04537_);
  and (_18889_, _18888_, _18880_);
  nor (_18890_, _05799_, _09032_);
  or (_18891_, _18890_, _18877_);
  and (_18893_, _18891_, _03755_);
  or (_18894_, _18893_, _18889_);
  and (_18895_, _18894_, _03751_);
  and (_18896_, _18883_, _03750_);
  or (_18897_, _18896_, _07544_);
  or (_18898_, _18897_, _18895_);
  or (_18899_, _18891_, _06994_);
  and (_18900_, _18899_, _18898_);
  or (_18901_, _18900_, _04678_);
  and (_18902_, _06941_, _05391_);
  or (_18904_, _18877_, _04679_);
  or (_18905_, _18904_, _18902_);
  and (_18906_, _18905_, _03415_);
  and (_18907_, _18906_, _18901_);
  nor (_18908_, _13118_, _09032_);
  or (_18909_, _18908_, _18877_);
  and (_18910_, _18909_, _07559_);
  or (_18911_, _18910_, _08854_);
  or (_18912_, _18911_, _18907_);
  and (_18913_, _13133_, _05391_);
  or (_18915_, _18877_, _04703_);
  or (_18916_, _18915_, _18913_);
  and (_18917_, _06371_, _05391_);
  or (_18918_, _18917_, _18877_);
  or (_18919_, _18918_, _04694_);
  and (_18920_, _18919_, _04701_);
  and (_18921_, _18920_, _18916_);
  and (_18922_, _18921_, _18912_);
  and (_18923_, _10451_, _05391_);
  or (_18924_, _18923_, _18877_);
  and (_18926_, _18924_, _03959_);
  or (_18927_, _18926_, _18922_);
  and (_18928_, _18927_, _04708_);
  or (_18929_, _18877_, _08302_);
  and (_18930_, _18918_, _03866_);
  and (_18931_, _18930_, _18929_);
  or (_18932_, _18931_, _18928_);
  and (_18933_, _18932_, _04706_);
  and (_18934_, _18883_, _03967_);
  and (_18935_, _18934_, _18929_);
  or (_18937_, _18935_, _03835_);
  or (_18938_, _18937_, _18933_);
  nor (_18939_, _13131_, _09032_);
  or (_18940_, _18877_, _06532_);
  or (_18941_, _18940_, _18939_);
  and (_18942_, _18941_, _06537_);
  and (_18943_, _18942_, _18938_);
  nor (_18944_, _08697_, _09032_);
  or (_18945_, _18944_, _18877_);
  and (_18946_, _18945_, _03954_);
  or (_18948_, _18946_, _18943_);
  and (_18949_, _18948_, _03704_);
  and (_18950_, _18879_, _03703_);
  or (_18951_, _18950_, _03701_);
  or (_18952_, _18951_, _18949_);
  and (_18953_, _13193_, _05391_);
  or (_18954_, _18953_, _18877_);
  or (_18955_, _18954_, _03702_);
  and (_18956_, _18955_, _18952_);
  or (_18957_, _18956_, _42912_);
  or (_18959_, _42908_, \oc8051_golden_model_1.PCON [5]);
  and (_18960_, _18959_, _41654_);
  and (_43177_, _18960_, _18957_);
  not (_18961_, \oc8051_golden_model_1.PCON [6]);
  nor (_18962_, _05391_, _18961_);
  and (_18963_, _13333_, _05391_);
  nor (_18964_, _18963_, _18962_);
  and (_18965_, _18964_, _03839_);
  nor (_18966_, _06013_, _09032_);
  nor (_18967_, _18966_, _18962_);
  and (_18969_, _18967_, _07544_);
  and (_18970_, _05391_, \oc8051_golden_model_1.ACC [6]);
  nor (_18971_, _18970_, _18962_);
  nor (_18972_, _18971_, _04616_);
  nor (_18973_, _04615_, _18961_);
  or (_18974_, _18973_, _18972_);
  and (_18975_, _18974_, _04630_);
  nor (_18976_, _13234_, _09032_);
  nor (_18977_, _18976_, _18962_);
  nor (_18978_, _18977_, _04630_);
  or (_18980_, _18978_, _18975_);
  and (_18981_, _18980_, _04537_);
  nor (_18982_, _18967_, _04537_);
  nor (_18983_, _18982_, _18981_);
  nor (_18984_, _18983_, _03750_);
  nor (_18985_, _18971_, _03751_);
  nor (_18986_, _18985_, _07544_);
  not (_18987_, _18986_);
  nor (_18988_, _18987_, _18984_);
  nor (_18989_, _18988_, _18969_);
  nor (_18991_, _18989_, _04678_);
  and (_18992_, _06933_, _05391_);
  nor (_18993_, _18962_, _04679_);
  not (_18994_, _18993_);
  nor (_18995_, _18994_, _18992_);
  or (_18996_, _18995_, _07559_);
  nor (_18997_, _18996_, _18991_);
  nor (_18998_, _13326_, _09032_);
  nor (_18999_, _18998_, _18962_);
  nor (_19000_, _18999_, _03415_);
  or (_19002_, _19000_, _03839_);
  nor (_19003_, _19002_, _18997_);
  nor (_19004_, _19003_, _18965_);
  or (_19005_, _19004_, _03838_);
  and (_19006_, _13341_, _05391_);
  or (_19007_, _18962_, _04703_);
  nor (_19008_, _19007_, _19006_);
  nor (_19009_, _19008_, _03959_);
  and (_19010_, _19009_, _19005_);
  and (_19011_, _08695_, _05391_);
  nor (_19013_, _19011_, _18962_);
  nor (_19014_, _19013_, _04701_);
  nor (_19015_, _19014_, _19010_);
  nor (_19016_, _19015_, _03866_);
  nor (_19017_, _18962_, _08289_);
  not (_19018_, _19017_);
  nor (_19019_, _18964_, _04708_);
  and (_19020_, _19019_, _19018_);
  nor (_19021_, _19020_, _19016_);
  nor (_19022_, _19021_, _03967_);
  nor (_19024_, _18971_, _04706_);
  and (_19025_, _19024_, _19018_);
  nor (_19026_, _19025_, _03835_);
  not (_19027_, _19026_);
  nor (_19028_, _19027_, _19022_);
  nor (_19029_, _13340_, _09032_);
  or (_19030_, _18962_, _06532_);
  nor (_19031_, _19030_, _19029_);
  or (_19032_, _19031_, _03954_);
  nor (_19033_, _19032_, _19028_);
  nor (_19035_, _08694_, _09032_);
  nor (_19036_, _19035_, _18962_);
  nor (_19037_, _19036_, _06537_);
  or (_19038_, _19037_, _03703_);
  nor (_19039_, _19038_, _19033_);
  and (_19040_, _18977_, _03703_);
  or (_19041_, _19040_, _03701_);
  nor (_19042_, _19041_, _19039_);
  nor (_19043_, _13399_, _09032_);
  nor (_19044_, _19043_, _18962_);
  nor (_19046_, _19044_, _03702_);
  or (_19047_, _19046_, _19042_);
  or (_19048_, _19047_, _42912_);
  or (_19049_, _42908_, \oc8051_golden_model_1.PCON [6]);
  and (_19050_, _19049_, _41654_);
  and (_43178_, _19050_, _19048_);
  not (_19051_, \oc8051_golden_model_1.TCON [0]);
  nor (_19052_, _05438_, _19051_);
  nor (_19053_, _05652_, _09090_);
  nor (_19054_, _19053_, _19052_);
  nor (_19056_, _19054_, _03702_);
  and (_19057_, _05438_, _06428_);
  nor (_19058_, _19057_, _19052_);
  and (_19059_, _19058_, _03839_);
  and (_19060_, _05438_, _04608_);
  nor (_19061_, _19060_, _19052_);
  and (_19062_, _19061_, _07544_);
  and (_19063_, _05438_, \oc8051_golden_model_1.ACC [0]);
  nor (_19064_, _19063_, _19052_);
  nor (_19065_, _19064_, _04616_);
  nor (_19067_, _04615_, _19051_);
  or (_19068_, _19067_, _19065_);
  and (_19069_, _19068_, _04630_);
  nor (_19070_, _19054_, _04630_);
  or (_19071_, _19070_, _19069_);
  and (_19072_, _19071_, _03697_);
  nor (_19073_, _06081_, _19051_);
  and (_19074_, _12032_, _06081_);
  nor (_19075_, _19074_, _19073_);
  nor (_19076_, _19075_, _03697_);
  nor (_19078_, _19076_, _19072_);
  nor (_19079_, _19078_, _03755_);
  nor (_19080_, _19061_, _04537_);
  or (_19081_, _19080_, _19079_);
  and (_19082_, _19081_, _03751_);
  nor (_19083_, _19064_, _03751_);
  or (_19084_, _19083_, _19082_);
  and (_19085_, _19084_, _03692_);
  and (_19086_, _19052_, _03691_);
  or (_19087_, _19086_, _19085_);
  and (_19089_, _19087_, _03685_);
  nor (_19090_, _19054_, _03685_);
  or (_19091_, _19090_, _19089_);
  and (_19092_, _19091_, _03680_);
  nor (_19093_, _19073_, _14175_);
  or (_19094_, _19093_, _03680_);
  or (_19095_, _19094_, _19075_);
  and (_19096_, _19095_, _06994_);
  not (_19097_, _19096_);
  nor (_19098_, _19097_, _19092_);
  nor (_19100_, _19098_, _19062_);
  nor (_19101_, _19100_, _04678_);
  and (_19102_, _06935_, _05438_);
  nor (_19103_, _19052_, _04679_);
  not (_19104_, _19103_);
  nor (_19105_, _19104_, _19102_);
  or (_19106_, _19105_, _07559_);
  nor (_19107_, _19106_, _19101_);
  nor (_19108_, _12119_, _09090_);
  nor (_19109_, _19108_, _19052_);
  nor (_19111_, _19109_, _03415_);
  or (_19112_, _19111_, _03839_);
  nor (_19113_, _19112_, _19107_);
  nor (_19114_, _19113_, _19059_);
  or (_19115_, _19114_, _03838_);
  and (_19116_, _12133_, _05438_);
  or (_19117_, _19052_, _04703_);
  nor (_19118_, _19117_, _19116_);
  nor (_19119_, _19118_, _03959_);
  and (_19120_, _19119_, _19115_);
  nor (_19122_, _10458_, _09090_);
  nor (_19123_, _19122_, _19052_);
  and (_19124_, _19063_, _05652_);
  or (_19125_, _19124_, _04701_);
  nor (_19126_, _19125_, _19123_);
  nor (_19127_, _19126_, _19120_);
  nor (_19128_, _19127_, _03866_);
  and (_19129_, _12013_, _05438_);
  or (_19130_, _19129_, _19052_);
  and (_19131_, _19130_, _03866_);
  or (_19133_, _19131_, _19128_);
  and (_19134_, _19133_, _04706_);
  nor (_19135_, _19124_, _19052_);
  nor (_19136_, _19135_, _04706_);
  or (_19137_, _19136_, _19134_);
  and (_19138_, _19137_, _06532_);
  nor (_19139_, _12132_, _09090_);
  nor (_19140_, _19139_, _19052_);
  nor (_19141_, _19140_, _06532_);
  or (_19142_, _19141_, _19138_);
  and (_19144_, _19142_, _06537_);
  nor (_19145_, _19123_, _06537_);
  or (_19146_, _19145_, _03703_);
  or (_19147_, _19146_, _19144_);
  nand (_19148_, _19054_, _03703_);
  and (_19149_, _19148_, _19147_);
  nor (_19150_, _19149_, _03384_);
  nor (_19151_, _19052_, _03385_);
  nor (_19152_, _19151_, _19150_);
  and (_19153_, _19152_, _03702_);
  nor (_19155_, _19153_, _19056_);
  nand (_19156_, _19155_, _42908_);
  or (_19157_, _42908_, \oc8051_golden_model_1.TCON [0]);
  and (_19158_, _19157_, _41654_);
  and (_43179_, _19158_, _19156_);
  and (_19159_, _09090_, \oc8051_golden_model_1.TCON [1]);
  nor (_19160_, _08710_, _09090_);
  or (_19161_, _19160_, _19159_);
  or (_19162_, _19161_, _06537_);
  and (_19163_, _05438_, _04813_);
  or (_19165_, _19163_, _19159_);
  or (_19166_, _19165_, _04537_);
  or (_19167_, _05438_, \oc8051_golden_model_1.TCON [1]);
  and (_19168_, _12225_, _05438_);
  not (_19169_, _19168_);
  and (_19170_, _19169_, _19167_);
  or (_19171_, _19170_, _04630_);
  and (_19172_, _05438_, \oc8051_golden_model_1.ACC [1]);
  or (_19173_, _19172_, _19159_);
  and (_19174_, _19173_, _04615_);
  and (_19176_, _04616_, \oc8051_golden_model_1.TCON [1]);
  or (_19177_, _19176_, _03757_);
  or (_19178_, _19177_, _19174_);
  and (_19179_, _19178_, _03697_);
  and (_19180_, _19179_, _19171_);
  and (_19181_, _09103_, \oc8051_golden_model_1.TCON [1]);
  and (_19182_, _12212_, _06081_);
  or (_19183_, _19182_, _19181_);
  and (_19184_, _19183_, _03696_);
  or (_19185_, _19184_, _03755_);
  or (_19187_, _19185_, _19180_);
  and (_19188_, _19187_, _19166_);
  or (_19189_, _19188_, _03750_);
  or (_19190_, _19173_, _03751_);
  and (_19191_, _19190_, _03692_);
  and (_19192_, _19191_, _19189_);
  and (_19193_, _12200_, _06081_);
  or (_19194_, _19193_, _19181_);
  and (_19195_, _19194_, _03691_);
  or (_19196_, _19195_, _03684_);
  or (_19198_, _19196_, _19192_);
  and (_19199_, _19182_, _12211_);
  or (_19200_, _19181_, _03685_);
  or (_19201_, _19200_, _19199_);
  and (_19202_, _19201_, _19198_);
  and (_19203_, _19202_, _03680_);
  nor (_19204_, _12256_, _09103_);
  or (_19205_, _19181_, _19204_);
  and (_19206_, _19205_, _03679_);
  or (_19207_, _19206_, _07544_);
  or (_19209_, _19207_, _19203_);
  or (_19210_, _19165_, _06994_);
  and (_19211_, _19210_, _19209_);
  or (_19212_, _19211_, _04678_);
  and (_19213_, _06934_, _05438_);
  or (_19214_, _19159_, _04679_);
  or (_19215_, _19214_, _19213_);
  and (_19216_, _19215_, _03415_);
  and (_19217_, _19216_, _19212_);
  nor (_19218_, _12313_, _09090_);
  or (_19220_, _19218_, _19159_);
  and (_19221_, _19220_, _07559_);
  or (_19222_, _19221_, _19217_);
  and (_19223_, _19222_, _03840_);
  or (_19224_, _12207_, _09090_);
  and (_19225_, _19224_, _03838_);
  nand (_19226_, _05438_, _04515_);
  and (_19227_, _19226_, _03839_);
  or (_19228_, _19227_, _19225_);
  and (_19229_, _19228_, _19167_);
  or (_19231_, _19229_, _03959_);
  or (_19232_, _19231_, _19223_);
  and (_19233_, _08711_, _05438_);
  or (_19234_, _19233_, _19159_);
  or (_19235_, _19234_, _04701_);
  and (_19236_, _19235_, _04708_);
  and (_19237_, _19236_, _19232_);
  or (_19238_, _12206_, _09090_);
  and (_19239_, _19167_, _03866_);
  and (_19240_, _19239_, _19238_);
  or (_19242_, _19240_, _03967_);
  or (_19243_, _19242_, _19237_);
  and (_19244_, _19172_, _05603_);
  or (_19245_, _19159_, _04706_);
  or (_19246_, _19245_, _19244_);
  and (_19247_, _19246_, _06532_);
  and (_19248_, _19247_, _19243_);
  or (_19249_, _19226_, _05603_);
  and (_19250_, _19167_, _03835_);
  and (_19251_, _19250_, _19249_);
  or (_19253_, _19251_, _03954_);
  or (_19254_, _19253_, _19248_);
  and (_19255_, _19254_, _19162_);
  or (_19256_, _19255_, _03703_);
  or (_19257_, _19170_, _03704_);
  and (_19258_, _19257_, _03385_);
  and (_19259_, _19258_, _19256_);
  and (_19260_, _19194_, _03384_);
  or (_19261_, _19260_, _03701_);
  or (_19262_, _19261_, _19259_);
  or (_19264_, _19168_, _19159_);
  or (_19265_, _19264_, _03702_);
  and (_19266_, _19265_, _19262_);
  and (_19267_, _19266_, _42908_);
  nor (_19268_, \oc8051_golden_model_1.TCON [1], rst);
  nor (_19269_, _19268_, _00000_);
  or (_43180_, _19269_, _19267_);
  not (_19270_, \oc8051_golden_model_1.TCON [2]);
  nor (_19271_, _05438_, _19270_);
  and (_19272_, _05438_, _06457_);
  nor (_19274_, _19272_, _19271_);
  and (_19275_, _19274_, _03839_);
  nor (_19276_, _09090_, _05236_);
  nor (_19277_, _19276_, _19271_);
  and (_19278_, _19277_, _07544_);
  and (_19279_, _05438_, \oc8051_golden_model_1.ACC [2]);
  nor (_19280_, _19279_, _19271_);
  nor (_19281_, _19280_, _04616_);
  nor (_19282_, _04615_, _19270_);
  or (_19283_, _19282_, _19281_);
  and (_19285_, _19283_, _04630_);
  nor (_19286_, _12427_, _09090_);
  nor (_19287_, _19286_, _19271_);
  nor (_19288_, _19287_, _04630_);
  or (_19289_, _19288_, _19285_);
  and (_19290_, _19289_, _03697_);
  nor (_19291_, _06081_, _19270_);
  and (_19292_, _12419_, _06081_);
  nor (_19293_, _19292_, _19291_);
  nor (_19294_, _19293_, _03697_);
  or (_19296_, _19294_, _19290_);
  and (_19297_, _19296_, _04537_);
  nor (_19298_, _19277_, _04537_);
  or (_19299_, _19298_, _19297_);
  and (_19300_, _19299_, _03751_);
  nor (_19301_, _19280_, _03751_);
  or (_19302_, _19301_, _19300_);
  and (_19303_, _19302_, _03692_);
  and (_19304_, _12422_, _06081_);
  nor (_19305_, _19304_, _19291_);
  nor (_19307_, _19305_, _03692_);
  or (_19308_, _19307_, _19303_);
  and (_19309_, _19308_, _03685_);
  and (_19310_, _19292_, _12418_);
  or (_19311_, _19310_, _19291_);
  and (_19312_, _19311_, _03684_);
  or (_19313_, _19312_, _19309_);
  and (_19314_, _19313_, _03680_);
  nor (_19315_, _12465_, _09103_);
  nor (_19316_, _19315_, _19291_);
  nor (_19318_, _19316_, _03680_);
  nor (_19319_, _19318_, _07544_);
  not (_19320_, _19319_);
  nor (_19321_, _19320_, _19314_);
  nor (_19322_, _19321_, _19278_);
  nor (_19323_, _19322_, _04678_);
  and (_19324_, _06938_, _05438_);
  nor (_19325_, _19271_, _04679_);
  not (_19326_, _19325_);
  nor (_19327_, _19326_, _19324_);
  or (_19329_, _19327_, _07559_);
  nor (_19330_, _19329_, _19323_);
  nor (_19331_, _12523_, _09090_);
  nor (_19332_, _19271_, _19331_);
  nor (_19333_, _19332_, _03415_);
  or (_19334_, _19333_, _03839_);
  nor (_19335_, _19334_, _19330_);
  nor (_19336_, _19335_, _19275_);
  or (_19337_, _19336_, _03838_);
  and (_19338_, _12537_, _05438_);
  or (_19340_, _19338_, _19271_);
  or (_19341_, _19340_, _04703_);
  and (_19342_, _19341_, _04701_);
  and (_19343_, _19342_, _19337_);
  and (_19344_, _08707_, _05438_);
  nor (_19345_, _19344_, _19271_);
  nor (_19346_, _19345_, _04701_);
  nor (_19347_, _19346_, _19343_);
  nor (_19348_, _19347_, _03866_);
  nor (_19349_, _19271_, _05700_);
  not (_19351_, _19349_);
  nor (_19352_, _19274_, _04708_);
  and (_19353_, _19352_, _19351_);
  nor (_19354_, _19353_, _19348_);
  nor (_19355_, _19354_, _03967_);
  nor (_19356_, _19280_, _04706_);
  and (_19357_, _19356_, _19351_);
  or (_19358_, _19357_, _19355_);
  and (_19359_, _19358_, _06532_);
  nor (_19360_, _12536_, _09090_);
  nor (_19362_, _19360_, _19271_);
  nor (_19363_, _19362_, _06532_);
  or (_19364_, _19363_, _19359_);
  and (_19365_, _19364_, _06537_);
  nor (_19366_, _08706_, _09090_);
  nor (_19367_, _19366_, _19271_);
  nor (_19368_, _19367_, _06537_);
  or (_19369_, _19368_, _19365_);
  and (_19370_, _19369_, _03704_);
  nor (_19371_, _19287_, _03704_);
  or (_19373_, _19371_, _19370_);
  and (_19374_, _19373_, _03385_);
  nor (_19375_, _19305_, _03385_);
  or (_19376_, _19375_, _19374_);
  and (_19377_, _19376_, _03702_);
  and (_19378_, _12596_, _05438_);
  nor (_19379_, _19378_, _19271_);
  nor (_19380_, _19379_, _03702_);
  or (_19381_, _19380_, _19377_);
  or (_19382_, _19381_, _42912_);
  or (_19384_, _42908_, \oc8051_golden_model_1.TCON [2]);
  and (_19385_, _19384_, _41654_);
  and (_43181_, _19385_, _19382_);
  and (_19386_, _09090_, \oc8051_golden_model_1.TCON [3]);
  nor (_19387_, _09090_, _05050_);
  or (_19388_, _19387_, _19386_);
  or (_19389_, _19388_, _06994_);
  nor (_19390_, _12610_, _09090_);
  or (_19391_, _19390_, _19386_);
  or (_19392_, _19391_, _04630_);
  and (_19394_, _05438_, \oc8051_golden_model_1.ACC [3]);
  or (_19395_, _19394_, _19386_);
  and (_19396_, _19395_, _04615_);
  and (_19397_, _04616_, \oc8051_golden_model_1.TCON [3]);
  or (_19398_, _19397_, _03757_);
  or (_19399_, _19398_, _19396_);
  and (_19400_, _19399_, _03697_);
  and (_19401_, _19400_, _19392_);
  and (_19402_, _09103_, \oc8051_golden_model_1.TCON [3]);
  and (_19403_, _12619_, _06081_);
  or (_19405_, _19403_, _19402_);
  and (_19406_, _19405_, _03696_);
  or (_19407_, _19406_, _03755_);
  or (_19408_, _19407_, _19401_);
  or (_19409_, _19388_, _04537_);
  and (_19410_, _19409_, _19408_);
  or (_19411_, _19410_, _03750_);
  or (_19412_, _19395_, _03751_);
  and (_19413_, _19412_, _03692_);
  and (_19414_, _19413_, _19411_);
  and (_19416_, _12622_, _06081_);
  or (_19417_, _19416_, _19402_);
  and (_19418_, _19417_, _03691_);
  or (_19419_, _19418_, _03684_);
  or (_19420_, _19419_, _19414_);
  or (_19421_, _19402_, _12618_);
  and (_19422_, _19421_, _19405_);
  or (_19423_, _19422_, _03685_);
  and (_19424_, _19423_, _03680_);
  and (_19425_, _19424_, _19420_);
  nor (_19427_, _12665_, _09103_);
  or (_19428_, _19427_, _19402_);
  and (_19429_, _19428_, _03679_);
  or (_19430_, _19429_, _07544_);
  or (_19431_, _19430_, _19425_);
  and (_19432_, _19431_, _19389_);
  or (_19433_, _19432_, _04678_);
  and (_19434_, _06937_, _05438_);
  or (_19435_, _19386_, _04679_);
  or (_19436_, _19435_, _19434_);
  and (_19438_, _19436_, _03415_);
  and (_19439_, _19438_, _19433_);
  nor (_19440_, _12724_, _09090_);
  or (_19441_, _19386_, _19440_);
  and (_19442_, _19441_, _07559_);
  or (_19443_, _19442_, _19439_);
  or (_19444_, _19443_, _08854_);
  and (_19445_, _12738_, _05438_);
  or (_19446_, _19386_, _04703_);
  or (_19447_, _19446_, _19445_);
  and (_19449_, _05438_, _06415_);
  or (_19450_, _19449_, _19386_);
  or (_19451_, _19450_, _04694_);
  and (_19452_, _19451_, _04701_);
  and (_19453_, _19452_, _19447_);
  and (_19454_, _19453_, _19444_);
  and (_19455_, _10455_, _05438_);
  or (_19456_, _19455_, _19386_);
  and (_19457_, _19456_, _03959_);
  or (_19458_, _19457_, _19454_);
  and (_19460_, _19458_, _04708_);
  or (_19461_, _19386_, _05554_);
  and (_19462_, _19450_, _03866_);
  and (_19463_, _19462_, _19461_);
  or (_19464_, _19463_, _19460_);
  and (_19465_, _19464_, _04706_);
  and (_19466_, _19395_, _03967_);
  and (_19467_, _19466_, _19461_);
  or (_19468_, _19467_, _03835_);
  or (_19469_, _19468_, _19465_);
  nor (_19471_, _12737_, _09090_);
  or (_19472_, _19386_, _06532_);
  or (_19473_, _19472_, _19471_);
  and (_19474_, _19473_, _06537_);
  and (_19475_, _19474_, _19469_);
  nor (_19476_, _08701_, _09090_);
  or (_19477_, _19476_, _19386_);
  and (_19478_, _19477_, _03954_);
  or (_19479_, _19478_, _03703_);
  or (_19480_, _19479_, _19475_);
  or (_19482_, _19391_, _03704_);
  and (_19483_, _19482_, _03385_);
  and (_19484_, _19483_, _19480_);
  and (_19485_, _19417_, _03384_);
  or (_19486_, _19485_, _03701_);
  or (_19487_, _19486_, _19484_);
  and (_19488_, _12792_, _05438_);
  or (_19489_, _19488_, _19386_);
  or (_19490_, _19489_, _03702_);
  and (_19491_, _19490_, _19487_);
  or (_19493_, _19491_, _42912_);
  or (_19494_, _42908_, \oc8051_golden_model_1.TCON [3]);
  and (_19495_, _19494_, _41654_);
  and (_43182_, _19495_, _19493_);
  and (_19496_, _09090_, \oc8051_golden_model_1.TCON [4]);
  nor (_19497_, _05898_, _09090_);
  or (_19498_, _19497_, _19496_);
  or (_19499_, _19498_, _06994_);
  and (_19500_, _09103_, \oc8051_golden_model_1.TCON [4]);
  and (_19501_, _12808_, _06081_);
  or (_19503_, _19501_, _19500_);
  and (_19504_, _19503_, _03691_);
  nor (_19505_, _12828_, _09090_);
  or (_19506_, _19505_, _19496_);
  or (_19507_, _19506_, _04630_);
  and (_19508_, _05438_, \oc8051_golden_model_1.ACC [4]);
  or (_19509_, _19508_, _19496_);
  and (_19510_, _19509_, _04615_);
  and (_19511_, _04616_, \oc8051_golden_model_1.TCON [4]);
  or (_19512_, _19511_, _03757_);
  or (_19514_, _19512_, _19510_);
  and (_19515_, _19514_, _03697_);
  and (_19516_, _19515_, _19507_);
  and (_19517_, _12832_, _06081_);
  or (_19518_, _19517_, _19500_);
  and (_19519_, _19518_, _03696_);
  or (_19520_, _19519_, _03755_);
  or (_19521_, _19520_, _19516_);
  or (_19522_, _19498_, _04537_);
  and (_19523_, _19522_, _19521_);
  or (_19525_, _19523_, _03750_);
  or (_19526_, _19509_, _03751_);
  and (_19527_, _19526_, _03692_);
  and (_19528_, _19527_, _19525_);
  or (_19529_, _19528_, _19504_);
  and (_19530_, _19529_, _03685_);
  or (_19531_, _19500_, _12847_);
  and (_19532_, _19531_, _03684_);
  and (_19533_, _19532_, _19518_);
  or (_19534_, _19533_, _19530_);
  and (_19536_, _19534_, _03680_);
  nor (_19537_, _12810_, _09103_);
  or (_19538_, _19537_, _19500_);
  and (_19539_, _19538_, _03679_);
  or (_19540_, _19539_, _07544_);
  or (_19541_, _19540_, _19536_);
  and (_19542_, _19541_, _19499_);
  or (_19543_, _19542_, _04678_);
  and (_19544_, _06942_, _05438_);
  or (_19545_, _19496_, _04679_);
  or (_19547_, _19545_, _19544_);
  and (_19548_, _19547_, _03415_);
  and (_19549_, _19548_, _19543_);
  nor (_19550_, _12919_, _09090_);
  or (_19551_, _19550_, _19496_);
  and (_19552_, _19551_, _07559_);
  or (_19553_, _19552_, _08854_);
  or (_19554_, _19553_, _19549_);
  and (_19555_, _12933_, _05438_);
  or (_19556_, _19496_, _04703_);
  or (_19558_, _19556_, _19555_);
  and (_19559_, _06422_, _05438_);
  or (_19560_, _19559_, _19496_);
  or (_19561_, _19560_, _04694_);
  and (_19562_, _19561_, _04701_);
  and (_19563_, _19562_, _19558_);
  and (_19564_, _19563_, _19554_);
  and (_19565_, _08700_, _05438_);
  or (_19566_, _19565_, _19496_);
  and (_19567_, _19566_, _03959_);
  or (_19569_, _19567_, _19564_);
  and (_19570_, _19569_, _04708_);
  or (_19571_, _19496_, _08303_);
  and (_19572_, _19560_, _03866_);
  and (_19573_, _19572_, _19571_);
  or (_19574_, _19573_, _19570_);
  and (_19575_, _19574_, _04706_);
  and (_19576_, _19509_, _03967_);
  and (_19577_, _19576_, _19571_);
  or (_19578_, _19577_, _03835_);
  or (_19580_, _19578_, _19575_);
  nor (_19581_, _12931_, _09090_);
  or (_19582_, _19496_, _06532_);
  or (_19583_, _19582_, _19581_);
  and (_19584_, _19583_, _06537_);
  and (_19585_, _19584_, _19580_);
  nor (_19586_, _08699_, _09090_);
  or (_19587_, _19586_, _19496_);
  and (_19588_, _19587_, _03954_);
  or (_19589_, _19588_, _03703_);
  or (_19591_, _19589_, _19585_);
  or (_19592_, _19506_, _03704_);
  and (_19593_, _19592_, _03385_);
  and (_19594_, _19593_, _19591_);
  and (_19595_, _19503_, _03384_);
  or (_19596_, _19595_, _03701_);
  or (_19597_, _19596_, _19594_);
  and (_19598_, _12991_, _05438_);
  or (_19599_, _19598_, _19496_);
  or (_19600_, _19599_, _03702_);
  and (_19602_, _19600_, _19597_);
  or (_19603_, _19602_, _42912_);
  or (_19604_, _42908_, \oc8051_golden_model_1.TCON [4]);
  and (_19605_, _19604_, _41654_);
  and (_43183_, _19605_, _19603_);
  and (_19606_, _09090_, \oc8051_golden_model_1.TCON [5]);
  nor (_19607_, _13025_, _09090_);
  or (_19608_, _19607_, _19606_);
  or (_19609_, _19608_, _04630_);
  and (_19610_, _05438_, \oc8051_golden_model_1.ACC [5]);
  or (_19612_, _19610_, _19606_);
  and (_19613_, _19612_, _04615_);
  and (_19614_, _04616_, \oc8051_golden_model_1.TCON [5]);
  or (_19615_, _19614_, _03757_);
  or (_19616_, _19615_, _19613_);
  and (_19617_, _19616_, _03697_);
  and (_19618_, _19617_, _19609_);
  and (_19619_, _09103_, \oc8051_golden_model_1.TCON [5]);
  and (_19620_, _13029_, _06081_);
  or (_19621_, _19620_, _19619_);
  and (_19623_, _19621_, _03696_);
  or (_19624_, _19623_, _03755_);
  or (_19625_, _19624_, _19618_);
  nor (_19626_, _05799_, _09090_);
  or (_19627_, _19626_, _19606_);
  or (_19628_, _19627_, _04537_);
  and (_19629_, _19628_, _19625_);
  or (_19630_, _19629_, _03750_);
  or (_19631_, _19612_, _03751_);
  and (_19632_, _19631_, _03692_);
  and (_19634_, _19632_, _19630_);
  and (_19635_, _13007_, _06081_);
  or (_19636_, _19635_, _19619_);
  and (_19637_, _19636_, _03691_);
  or (_19638_, _19637_, _03684_);
  or (_19639_, _19638_, _19634_);
  or (_19640_, _19619_, _13044_);
  and (_19641_, _19640_, _19621_);
  or (_19642_, _19641_, _03685_);
  and (_19643_, _19642_, _03680_);
  and (_19645_, _19643_, _19639_);
  nor (_19646_, _13009_, _09103_);
  or (_19647_, _19646_, _19619_);
  and (_19648_, _19647_, _03679_);
  or (_19649_, _19648_, _07544_);
  or (_19650_, _19649_, _19645_);
  or (_19651_, _19627_, _06994_);
  and (_19652_, _19651_, _19650_);
  or (_19653_, _19652_, _04678_);
  and (_19654_, _06941_, _05438_);
  or (_19656_, _19606_, _04679_);
  or (_19657_, _19656_, _19654_);
  and (_19658_, _19657_, _03415_);
  and (_19659_, _19658_, _19653_);
  nor (_19660_, _13118_, _09090_);
  or (_19661_, _19660_, _19606_);
  and (_19662_, _19661_, _07559_);
  or (_19663_, _19662_, _08854_);
  or (_19664_, _19663_, _19659_);
  and (_19665_, _13133_, _05438_);
  or (_19667_, _19606_, _04703_);
  or (_19668_, _19667_, _19665_);
  and (_19669_, _06371_, _05438_);
  or (_19670_, _19669_, _19606_);
  or (_19671_, _19670_, _04694_);
  and (_19672_, _19671_, _04701_);
  and (_19673_, _19672_, _19668_);
  and (_19674_, _19673_, _19664_);
  and (_19675_, _10451_, _05438_);
  or (_19676_, _19675_, _19606_);
  and (_19678_, _19676_, _03959_);
  or (_19679_, _19678_, _19674_);
  and (_19680_, _19679_, _04708_);
  or (_19681_, _19606_, _08302_);
  and (_19682_, _19670_, _03866_);
  and (_19683_, _19682_, _19681_);
  or (_19684_, _19683_, _19680_);
  and (_19685_, _19684_, _04706_);
  and (_19686_, _19612_, _03967_);
  and (_19687_, _19686_, _19681_);
  or (_19689_, _19687_, _03835_);
  or (_19690_, _19689_, _19685_);
  nor (_19691_, _13131_, _09090_);
  or (_19692_, _19606_, _06532_);
  or (_19693_, _19692_, _19691_);
  and (_19694_, _19693_, _06537_);
  and (_19695_, _19694_, _19690_);
  nor (_19696_, _08697_, _09090_);
  or (_19697_, _19696_, _19606_);
  and (_19698_, _19697_, _03954_);
  or (_19700_, _19698_, _03703_);
  or (_19701_, _19700_, _19695_);
  or (_19702_, _19608_, _03704_);
  and (_19703_, _19702_, _03385_);
  and (_19704_, _19703_, _19701_);
  and (_19705_, _19636_, _03384_);
  or (_19706_, _19705_, _03701_);
  or (_19707_, _19706_, _19704_);
  and (_19708_, _13193_, _05438_);
  or (_19709_, _19708_, _19606_);
  or (_19711_, _19709_, _03702_);
  and (_19712_, _19711_, _19707_);
  or (_19713_, _19712_, _42912_);
  or (_19714_, _42908_, \oc8051_golden_model_1.TCON [5]);
  and (_19715_, _19714_, _41654_);
  and (_43184_, _19715_, _19713_);
  and (_19716_, _09090_, \oc8051_golden_model_1.TCON [6]);
  nor (_19717_, _06013_, _09090_);
  or (_19718_, _19717_, _19716_);
  or (_19719_, _19718_, _06994_);
  and (_19721_, _09103_, \oc8051_golden_model_1.TCON [6]);
  and (_19722_, _13218_, _06081_);
  or (_19723_, _19722_, _19721_);
  and (_19724_, _19723_, _03691_);
  nor (_19725_, _13234_, _09090_);
  or (_19726_, _19725_, _19716_);
  or (_19727_, _19726_, _04630_);
  and (_19728_, _05438_, \oc8051_golden_model_1.ACC [6]);
  or (_19729_, _19728_, _19716_);
  and (_19730_, _19729_, _04615_);
  and (_19732_, _04616_, \oc8051_golden_model_1.TCON [6]);
  or (_19733_, _19732_, _03757_);
  or (_19734_, _19733_, _19730_);
  and (_19735_, _19734_, _03697_);
  and (_19736_, _19735_, _19727_);
  and (_19737_, _13238_, _06081_);
  or (_19738_, _19737_, _19721_);
  and (_19739_, _19738_, _03696_);
  or (_19740_, _19739_, _03755_);
  or (_19741_, _19740_, _19736_);
  or (_19743_, _19718_, _04537_);
  and (_19744_, _19743_, _19741_);
  or (_19745_, _19744_, _03750_);
  or (_19746_, _19729_, _03751_);
  and (_19747_, _19746_, _03692_);
  and (_19748_, _19747_, _19745_);
  or (_19749_, _19748_, _19724_);
  and (_19750_, _19749_, _03685_);
  and (_19751_, _13254_, _06081_);
  or (_19752_, _19751_, _19721_);
  and (_19754_, _19752_, _03684_);
  or (_19755_, _19754_, _19750_);
  and (_19756_, _19755_, _03680_);
  nor (_19757_, _13220_, _09103_);
  or (_19758_, _19757_, _19721_);
  and (_19759_, _19758_, _03679_);
  or (_19760_, _19759_, _07544_);
  or (_19761_, _19760_, _19756_);
  and (_19762_, _19761_, _19719_);
  or (_19763_, _19762_, _04678_);
  and (_19765_, _06933_, _05438_);
  or (_19766_, _19716_, _04679_);
  or (_19767_, _19766_, _19765_);
  and (_19768_, _19767_, _03415_);
  and (_19769_, _19768_, _19763_);
  nor (_19770_, _13326_, _09090_);
  or (_19771_, _19770_, _19716_);
  and (_19772_, _19771_, _07559_);
  or (_19773_, _19772_, _08854_);
  or (_19774_, _19773_, _19769_);
  and (_19776_, _13341_, _05438_);
  or (_19777_, _19716_, _04703_);
  or (_19778_, _19777_, _19776_);
  and (_19779_, _13333_, _05438_);
  or (_19780_, _19779_, _19716_);
  or (_19781_, _19780_, _04694_);
  and (_19782_, _19781_, _04701_);
  and (_19783_, _19782_, _19778_);
  and (_19784_, _19783_, _19774_);
  and (_19785_, _08695_, _05438_);
  or (_19787_, _19785_, _19716_);
  and (_19788_, _19787_, _03959_);
  or (_19789_, _19788_, _19784_);
  and (_19790_, _19789_, _04708_);
  or (_19791_, _19716_, _08289_);
  and (_19792_, _19780_, _03866_);
  and (_19793_, _19792_, _19791_);
  or (_19794_, _19793_, _19790_);
  and (_19795_, _19794_, _04706_);
  and (_19796_, _19729_, _03967_);
  and (_19798_, _19796_, _19791_);
  or (_19799_, _19798_, _03835_);
  or (_19800_, _19799_, _19795_);
  nor (_19801_, _13340_, _09090_);
  or (_19802_, _19716_, _06532_);
  or (_19803_, _19802_, _19801_);
  and (_19804_, _19803_, _06537_);
  and (_19805_, _19804_, _19800_);
  nor (_19806_, _08694_, _09090_);
  or (_19807_, _19806_, _19716_);
  and (_19809_, _19807_, _03954_);
  or (_19810_, _19809_, _03703_);
  or (_19811_, _19810_, _19805_);
  or (_19812_, _19726_, _03704_);
  and (_19813_, _19812_, _03385_);
  and (_19814_, _19813_, _19811_);
  and (_19815_, _19723_, _03384_);
  or (_19816_, _19815_, _03701_);
  or (_19817_, _19816_, _19814_);
  nor (_19818_, _13399_, _09090_);
  or (_19820_, _19818_, _19716_);
  or (_19821_, _19820_, _03702_);
  and (_19822_, _19821_, _19817_);
  or (_19823_, _19822_, _42912_);
  or (_19824_, _42908_, \oc8051_golden_model_1.TCON [6]);
  and (_19825_, _19824_, _41654_);
  and (_43185_, _19825_, _19823_);
  not (_19826_, \oc8051_golden_model_1.TL0 [0]);
  nor (_19827_, _05411_, _19826_);
  nor (_19828_, _05652_, _09215_);
  nor (_19830_, _19828_, _19827_);
  and (_19831_, _19830_, _17066_);
  and (_19832_, _05411_, \oc8051_golden_model_1.ACC [0]);
  nor (_19833_, _19832_, _19827_);
  nor (_19834_, _19833_, _03751_);
  nor (_19835_, _19834_, _07544_);
  nor (_19836_, _19830_, _04630_);
  nor (_19837_, _04615_, _19826_);
  nor (_19838_, _19833_, _04616_);
  nor (_19839_, _19838_, _19837_);
  nor (_19841_, _19839_, _03757_);
  or (_19842_, _19841_, _03755_);
  nor (_19843_, _19842_, _19836_);
  or (_19844_, _19843_, _03750_);
  and (_19845_, _19844_, _19835_);
  and (_19846_, _05411_, _04608_);
  and (_19847_, _06994_, _04537_);
  or (_19848_, _19847_, _19827_);
  nor (_19849_, _19848_, _19846_);
  nor (_19850_, _19849_, _19845_);
  nor (_19852_, _19850_, _04678_);
  and (_19853_, _06935_, _05411_);
  nor (_19854_, _19827_, _04679_);
  not (_19855_, _19854_);
  nor (_19856_, _19855_, _19853_);
  nor (_19857_, _19856_, _19852_);
  and (_19858_, _19857_, _03415_);
  nor (_19859_, _12119_, _09215_);
  nor (_19860_, _19859_, _19827_);
  nor (_19861_, _19860_, _03415_);
  or (_19863_, _19861_, _19858_);
  and (_19864_, _19863_, _04694_);
  and (_19865_, _05411_, _06428_);
  nor (_19866_, _19865_, _19827_);
  nor (_19867_, _19866_, _04694_);
  or (_19868_, _19867_, _19864_);
  and (_19869_, _19868_, _04703_);
  and (_19870_, _12133_, _05411_);
  nor (_19871_, _19870_, _19827_);
  nor (_19872_, _19871_, _04703_);
  or (_19874_, _19872_, _19869_);
  and (_19875_, _19874_, _04701_);
  nor (_19876_, _10458_, _09215_);
  nor (_19877_, _19876_, _19827_);
  not (_19878_, _19877_);
  and (_19879_, _08712_, _05411_);
  nor (_19880_, _19879_, _04701_);
  and (_19881_, _19880_, _19878_);
  nor (_19882_, _19881_, _19875_);
  nor (_19883_, _19882_, _03866_);
  and (_19885_, _12013_, _05411_);
  or (_19886_, _19885_, _19827_);
  and (_19887_, _19886_, _03866_);
  or (_19888_, _19887_, _19883_);
  and (_19889_, _19888_, _04706_);
  nor (_19890_, _19879_, _19827_);
  nor (_19891_, _19890_, _04706_);
  or (_19892_, _19891_, _19889_);
  and (_19893_, _19892_, _06532_);
  nor (_19894_, _12132_, _09215_);
  nor (_19896_, _19894_, _19827_);
  nor (_19897_, _19896_, _06532_);
  or (_19898_, _19897_, _19893_);
  and (_19899_, _19898_, _06537_);
  nor (_19900_, _19877_, _06537_);
  nor (_19901_, _19900_, _17066_);
  not (_19902_, _19901_);
  nor (_19903_, _19902_, _19899_);
  nor (_19904_, _19903_, _19831_);
  or (_19905_, _19904_, _42912_);
  or (_19907_, _42908_, \oc8051_golden_model_1.TL0 [0]);
  and (_19908_, _19907_, _41654_);
  and (_43188_, _19908_, _19905_);
  and (_19909_, _06934_, _05411_);
  not (_19910_, \oc8051_golden_model_1.TL0 [1]);
  nor (_19911_, _05411_, _19910_);
  nor (_19912_, _19911_, _04679_);
  not (_19913_, _19912_);
  nor (_19914_, _19913_, _19909_);
  not (_19915_, _19914_);
  and (_19917_, _05411_, \oc8051_golden_model_1.ACC [1]);
  nor (_19918_, _19917_, _19911_);
  nor (_19919_, _19918_, _03751_);
  nor (_19920_, _19918_, _04616_);
  nor (_19921_, _04615_, _19910_);
  or (_19922_, _19921_, _19920_);
  and (_19923_, _19922_, _04630_);
  nor (_19924_, _05411_, \oc8051_golden_model_1.TL0 [1]);
  and (_19925_, _12225_, _05411_);
  nor (_19926_, _19925_, _19924_);
  and (_19928_, _19926_, _03757_);
  or (_19929_, _19928_, _19923_);
  and (_19930_, _19929_, _04537_);
  and (_19931_, _05411_, _04813_);
  nor (_19932_, _19931_, _19911_);
  nor (_19933_, _19932_, _04537_);
  nor (_19934_, _19933_, _19930_);
  nor (_19935_, _19934_, _03750_);
  or (_19936_, _19935_, _07544_);
  nor (_19937_, _19936_, _19919_);
  and (_19939_, _19932_, _07544_);
  nor (_19940_, _19939_, _19937_);
  nor (_19941_, _19940_, _04678_);
  nor (_19942_, _19941_, _07559_);
  and (_19943_, _19942_, _19915_);
  and (_19944_, _12313_, _05411_);
  or (_19945_, _19944_, _03415_);
  nor (_19946_, _19945_, _19924_);
  nor (_19947_, _19946_, _19943_);
  nor (_19948_, _19947_, _08854_);
  nor (_19950_, _12207_, _09215_);
  or (_19951_, _19950_, _04703_);
  and (_19952_, _05411_, _04515_);
  or (_19953_, _19952_, _04694_);
  and (_19954_, _19953_, _19951_);
  nor (_19955_, _19954_, _19924_);
  or (_19956_, _19955_, _03959_);
  nor (_19957_, _19956_, _19948_);
  nor (_19958_, _08710_, _09215_);
  nor (_19959_, _19958_, _19911_);
  and (_19961_, _08709_, _05411_);
  nor (_19962_, _19961_, _19959_);
  nor (_19963_, _19962_, _04701_);
  nor (_19964_, _19963_, _03866_);
  not (_19965_, _19964_);
  nor (_19966_, _19965_, _19957_);
  and (_19967_, _12206_, _05411_);
  or (_19968_, _19967_, _19911_);
  and (_19969_, _19968_, _03866_);
  or (_19970_, _19969_, _19966_);
  and (_19972_, _19970_, _04706_);
  nor (_19973_, _19961_, _19911_);
  nor (_19974_, _19973_, _04706_);
  or (_19975_, _19974_, _19972_);
  and (_19976_, _19975_, _06532_);
  nor (_19977_, _12205_, _09215_);
  or (_19978_, _19977_, _19911_);
  and (_19979_, _19978_, _03835_);
  or (_19980_, _19979_, _19976_);
  and (_19981_, _19980_, _06537_);
  nor (_19983_, _19959_, _06537_);
  or (_19984_, _19983_, _19981_);
  and (_19985_, _19984_, _03704_);
  and (_19986_, _19926_, _03703_);
  or (_19987_, _19986_, _19985_);
  and (_19988_, _19987_, _03702_);
  nor (_19989_, _19925_, _19911_);
  nor (_19990_, _19989_, _03702_);
  nor (_19991_, _19990_, _19988_);
  nand (_19992_, _19991_, _42908_);
  or (_19994_, _42908_, \oc8051_golden_model_1.TL0 [1]);
  and (_19995_, _19994_, _41654_);
  and (_43189_, _19995_, _19992_);
  not (_19996_, \oc8051_golden_model_1.TL0 [2]);
  nor (_19997_, _05411_, _19996_);
  nor (_19998_, _09215_, _05236_);
  nor (_19999_, _19998_, _19997_);
  and (_20000_, _19999_, _07544_);
  and (_20001_, _05411_, \oc8051_golden_model_1.ACC [2]);
  nor (_20002_, _20001_, _19997_);
  nor (_20004_, _20002_, _03751_);
  nor (_20005_, _20002_, _04616_);
  nor (_20006_, _04615_, _19996_);
  or (_20007_, _20006_, _20005_);
  and (_20008_, _20007_, _04630_);
  nor (_20009_, _12427_, _09215_);
  nor (_20010_, _20009_, _19997_);
  nor (_20011_, _20010_, _04630_);
  or (_20012_, _20011_, _20008_);
  and (_20013_, _20012_, _04537_);
  nor (_20015_, _19999_, _04537_);
  nor (_20016_, _20015_, _20013_);
  nor (_20017_, _20016_, _03750_);
  or (_20018_, _20017_, _07544_);
  nor (_20019_, _20018_, _20004_);
  nor (_20020_, _20019_, _20000_);
  nor (_20021_, _20020_, _04678_);
  and (_20022_, _06938_, _05411_);
  nor (_20023_, _19997_, _04679_);
  not (_20024_, _20023_);
  nor (_20026_, _20024_, _20022_);
  nor (_20027_, _20026_, _07559_);
  not (_20028_, _20027_);
  nor (_20029_, _20028_, _20021_);
  nor (_20030_, _12523_, _09215_);
  nor (_20031_, _20030_, _19997_);
  nor (_20032_, _20031_, _03415_);
  or (_20033_, _20032_, _08854_);
  or (_20034_, _20033_, _20029_);
  and (_20035_, _12537_, _05411_);
  or (_20037_, _19997_, _04703_);
  or (_20038_, _20037_, _20035_);
  and (_20039_, _05411_, _06457_);
  nor (_20040_, _20039_, _19997_);
  and (_20041_, _20040_, _03839_);
  nor (_20042_, _20041_, _03959_);
  and (_20043_, _20042_, _20038_);
  and (_20044_, _20043_, _20034_);
  and (_20045_, _08707_, _05411_);
  nor (_20046_, _20045_, _19997_);
  nor (_20048_, _20046_, _04701_);
  nor (_20049_, _20048_, _20044_);
  nor (_20050_, _20049_, _03866_);
  nor (_20051_, _19997_, _05700_);
  not (_20052_, _20051_);
  nor (_20053_, _20040_, _04708_);
  and (_20054_, _20053_, _20052_);
  nor (_20055_, _20054_, _20050_);
  nor (_20056_, _20055_, _03967_);
  nor (_20057_, _20002_, _04706_);
  and (_20059_, _20057_, _20052_);
  nor (_20060_, _20059_, _03835_);
  not (_20061_, _20060_);
  nor (_20062_, _20061_, _20056_);
  nor (_20063_, _12536_, _09215_);
  or (_20064_, _19997_, _06532_);
  nor (_20065_, _20064_, _20063_);
  or (_20066_, _20065_, _03954_);
  nor (_20067_, _20066_, _20062_);
  nor (_20068_, _08706_, _09215_);
  nor (_20070_, _20068_, _19997_);
  nor (_20071_, _20070_, _06537_);
  or (_20072_, _20071_, _03703_);
  nor (_20073_, _20072_, _20067_);
  and (_20074_, _20010_, _03703_);
  or (_20075_, _20074_, _03701_);
  nor (_20076_, _20075_, _20073_);
  and (_20077_, _12596_, _05411_);
  nor (_20078_, _20077_, _19997_);
  nor (_20079_, _20078_, _03702_);
  or (_20081_, _20079_, _20076_);
  or (_20082_, _20081_, _42912_);
  or (_20083_, _42908_, \oc8051_golden_model_1.TL0 [2]);
  and (_20084_, _20083_, _41654_);
  and (_43190_, _20084_, _20082_);
  and (_20085_, _09215_, \oc8051_golden_model_1.TL0 [3]);
  nor (_20086_, _12610_, _09215_);
  or (_20087_, _20086_, _20085_);
  or (_20088_, _20087_, _04630_);
  and (_20089_, _05411_, \oc8051_golden_model_1.ACC [3]);
  or (_20091_, _20089_, _20085_);
  and (_20092_, _20091_, _04615_);
  and (_20093_, _04616_, \oc8051_golden_model_1.TL0 [3]);
  or (_20094_, _20093_, _03757_);
  or (_20095_, _20094_, _20092_);
  and (_20096_, _20095_, _04537_);
  and (_20097_, _20096_, _20088_);
  nor (_20098_, _09215_, _05050_);
  or (_20099_, _20098_, _20085_);
  and (_20100_, _20099_, _03755_);
  or (_20102_, _20100_, _20097_);
  and (_20103_, _20102_, _03751_);
  and (_20104_, _20091_, _03750_);
  or (_20105_, _20104_, _07544_);
  or (_20106_, _20105_, _20103_);
  or (_20107_, _20099_, _06994_);
  and (_20108_, _20107_, _20106_);
  or (_20109_, _20108_, _04678_);
  and (_20110_, _06937_, _05411_);
  or (_20111_, _20085_, _04679_);
  or (_20113_, _20111_, _20110_);
  and (_20114_, _20113_, _03415_);
  and (_20115_, _20114_, _20109_);
  nor (_20116_, _12724_, _09215_);
  or (_20117_, _20116_, _20085_);
  and (_20118_, _20117_, _07559_);
  or (_20119_, _20118_, _08854_);
  or (_20120_, _20119_, _20115_);
  and (_20121_, _12738_, _05411_);
  or (_20122_, _20085_, _04703_);
  or (_20124_, _20122_, _20121_);
  and (_20125_, _05411_, _06415_);
  or (_20126_, _20125_, _20085_);
  or (_20127_, _20126_, _04694_);
  and (_20128_, _20127_, _04701_);
  and (_20129_, _20128_, _20124_);
  and (_20130_, _20129_, _20120_);
  and (_20131_, _10455_, _05411_);
  or (_20132_, _20131_, _20085_);
  and (_20133_, _20132_, _03959_);
  or (_20135_, _20133_, _20130_);
  and (_20136_, _20135_, _04708_);
  or (_20137_, _20085_, _05554_);
  and (_20138_, _20126_, _03866_);
  and (_20139_, _20138_, _20137_);
  or (_20140_, _20139_, _20136_);
  and (_20141_, _20140_, _04706_);
  and (_20142_, _20091_, _03967_);
  and (_20143_, _20142_, _20137_);
  or (_20144_, _20143_, _03835_);
  or (_20146_, _20144_, _20141_);
  nor (_20147_, _12737_, _09215_);
  or (_20148_, _20085_, _06532_);
  or (_20149_, _20148_, _20147_);
  and (_20150_, _20149_, _06537_);
  and (_20151_, _20150_, _20146_);
  nor (_20152_, _08701_, _09215_);
  or (_20153_, _20152_, _20085_);
  and (_20154_, _20153_, _03954_);
  or (_20155_, _20154_, _03703_);
  or (_20157_, _20155_, _20151_);
  or (_20158_, _20087_, _03704_);
  and (_20159_, _20158_, _03702_);
  and (_20160_, _20159_, _20157_);
  and (_20161_, _12792_, _05411_);
  or (_20162_, _20161_, _20085_);
  and (_20163_, _20162_, _03701_);
  or (_20164_, _20163_, _20160_);
  or (_20165_, _20164_, _42912_);
  or (_20166_, _42908_, \oc8051_golden_model_1.TL0 [3]);
  and (_20168_, _20166_, _41654_);
  and (_43191_, _20168_, _20165_);
  not (_20169_, \oc8051_golden_model_1.TL0 [4]);
  nor (_20170_, _05411_, _20169_);
  and (_20171_, _06422_, _05411_);
  nor (_20172_, _20171_, _20170_);
  and (_20173_, _20172_, _03839_);
  nor (_20174_, _05898_, _09215_);
  nor (_20175_, _20174_, _20170_);
  and (_20176_, _20175_, _07544_);
  and (_20178_, _05411_, \oc8051_golden_model_1.ACC [4]);
  nor (_20179_, _20178_, _20170_);
  nor (_20180_, _20179_, _03751_);
  nor (_20181_, _20179_, _04616_);
  nor (_20182_, _04615_, _20169_);
  or (_20183_, _20182_, _20181_);
  and (_20184_, _20183_, _04630_);
  nor (_20185_, _12828_, _09215_);
  nor (_20186_, _20185_, _20170_);
  nor (_20187_, _20186_, _04630_);
  or (_20189_, _20187_, _20184_);
  and (_20190_, _20189_, _04537_);
  nor (_20191_, _20175_, _04537_);
  nor (_20192_, _20191_, _20190_);
  nor (_20193_, _20192_, _03750_);
  or (_20194_, _20193_, _07544_);
  nor (_20195_, _20194_, _20180_);
  nor (_20196_, _20195_, _20176_);
  nor (_20197_, _20196_, _04678_);
  and (_20198_, _06942_, _05411_);
  nor (_20200_, _20170_, _04679_);
  not (_20201_, _20200_);
  nor (_20202_, _20201_, _20198_);
  or (_20203_, _20202_, _07559_);
  nor (_20204_, _20203_, _20197_);
  nor (_20205_, _12919_, _09215_);
  nor (_20206_, _20205_, _20170_);
  nor (_20207_, _20206_, _03415_);
  or (_20208_, _20207_, _03839_);
  nor (_20209_, _20208_, _20204_);
  nor (_20211_, _20209_, _20173_);
  or (_20212_, _20211_, _03838_);
  and (_20213_, _12933_, _05411_);
  or (_20214_, _20170_, _04703_);
  nor (_20215_, _20214_, _20213_);
  nor (_20216_, _20215_, _03959_);
  and (_20217_, _20216_, _20212_);
  and (_20218_, _08700_, _05411_);
  nor (_20219_, _20218_, _20170_);
  nor (_20220_, _20219_, _04701_);
  nor (_20222_, _20220_, _20217_);
  nor (_20223_, _20222_, _03866_);
  nor (_20224_, _20170_, _08303_);
  not (_20225_, _20224_);
  nor (_20226_, _20172_, _04708_);
  and (_20227_, _20226_, _20225_);
  nor (_20228_, _20227_, _20223_);
  nor (_20229_, _20228_, _03967_);
  nor (_20230_, _20179_, _04706_);
  and (_20231_, _20230_, _20225_);
  nor (_20233_, _20231_, _03835_);
  not (_20234_, _20233_);
  nor (_20235_, _20234_, _20229_);
  nor (_20236_, _12931_, _09215_);
  or (_20237_, _20170_, _06532_);
  nor (_20238_, _20237_, _20236_);
  or (_20239_, _20238_, _03954_);
  nor (_20240_, _20239_, _20235_);
  nor (_20241_, _08699_, _09215_);
  nor (_20242_, _20241_, _20170_);
  nor (_20244_, _20242_, _06537_);
  or (_20245_, _20244_, _03703_);
  nor (_20246_, _20245_, _20240_);
  and (_20247_, _20186_, _03703_);
  or (_20248_, _20247_, _03701_);
  nor (_20249_, _20248_, _20246_);
  and (_20250_, _12991_, _05411_);
  nor (_20251_, _20250_, _20170_);
  nor (_20252_, _20251_, _03702_);
  or (_20253_, _20252_, _20249_);
  or (_20255_, _20253_, _42912_);
  or (_20256_, _42908_, \oc8051_golden_model_1.TL0 [4]);
  and (_20257_, _20256_, _41654_);
  and (_43192_, _20257_, _20255_);
  and (_20258_, _09215_, \oc8051_golden_model_1.TL0 [5]);
  nor (_20259_, _13025_, _09215_);
  or (_20260_, _20259_, _20258_);
  or (_20261_, _20260_, _04630_);
  and (_20262_, _05411_, \oc8051_golden_model_1.ACC [5]);
  or (_20263_, _20262_, _20258_);
  and (_20265_, _20263_, _04615_);
  and (_20266_, _04616_, \oc8051_golden_model_1.TL0 [5]);
  or (_20267_, _20266_, _03757_);
  or (_20268_, _20267_, _20265_);
  and (_20269_, _20268_, _04537_);
  and (_20270_, _20269_, _20261_);
  nor (_20271_, _05799_, _09215_);
  or (_20272_, _20271_, _20258_);
  and (_20273_, _20272_, _03755_);
  or (_20274_, _20273_, _20270_);
  and (_20276_, _20274_, _03751_);
  and (_20277_, _20263_, _03750_);
  or (_20278_, _20277_, _07544_);
  or (_20279_, _20278_, _20276_);
  or (_20280_, _20272_, _06994_);
  and (_20281_, _20280_, _20279_);
  or (_20282_, _20281_, _04678_);
  and (_20283_, _06941_, _05411_);
  or (_20284_, _20258_, _04679_);
  or (_20285_, _20284_, _20283_);
  and (_20287_, _20285_, _03415_);
  and (_20288_, _20287_, _20282_);
  nor (_20289_, _13118_, _09215_);
  or (_20290_, _20289_, _20258_);
  and (_20291_, _20290_, _07559_);
  or (_20292_, _20291_, _08854_);
  or (_20293_, _20292_, _20288_);
  and (_20294_, _13133_, _05411_);
  or (_20295_, _20258_, _04703_);
  or (_20296_, _20295_, _20294_);
  and (_20298_, _06371_, _05411_);
  or (_20299_, _20298_, _20258_);
  or (_20300_, _20299_, _04694_);
  and (_20301_, _20300_, _04701_);
  and (_20302_, _20301_, _20296_);
  and (_20303_, _20302_, _20293_);
  and (_20304_, _10451_, _05411_);
  or (_20305_, _20304_, _20258_);
  and (_20306_, _20305_, _03959_);
  or (_20307_, _20306_, _20303_);
  and (_20309_, _20307_, _04708_);
  or (_20310_, _20258_, _08302_);
  and (_20311_, _20299_, _03866_);
  and (_20312_, _20311_, _20310_);
  or (_20313_, _20312_, _20309_);
  and (_20314_, _20313_, _04706_);
  and (_20315_, _20263_, _03967_);
  and (_20316_, _20315_, _20310_);
  or (_20317_, _20316_, _03835_);
  or (_20318_, _20317_, _20314_);
  nor (_20320_, _13131_, _09215_);
  or (_20321_, _20258_, _06532_);
  or (_20322_, _20321_, _20320_);
  and (_20323_, _20322_, _06537_);
  and (_20324_, _20323_, _20318_);
  nor (_20325_, _08697_, _09215_);
  or (_20326_, _20325_, _20258_);
  and (_20327_, _20326_, _03954_);
  or (_20328_, _20327_, _20324_);
  and (_20329_, _20328_, _03704_);
  and (_20331_, _20260_, _03703_);
  or (_20332_, _20331_, _03701_);
  or (_20333_, _20332_, _20329_);
  and (_20334_, _13193_, _05411_);
  or (_20335_, _20334_, _20258_);
  or (_20336_, _20335_, _03702_);
  and (_20337_, _20336_, _20333_);
  or (_20338_, _20337_, _42912_);
  or (_20339_, _42908_, \oc8051_golden_model_1.TL0 [5]);
  and (_20340_, _20339_, _41654_);
  and (_43195_, _20340_, _20338_);
  not (_20342_, \oc8051_golden_model_1.TL0 [6]);
  nor (_20343_, _05411_, _20342_);
  and (_20344_, _13333_, _05411_);
  nor (_20345_, _20344_, _20343_);
  and (_20346_, _20345_, _03839_);
  and (_20347_, _05411_, \oc8051_golden_model_1.ACC [6]);
  nor (_20348_, _20347_, _20343_);
  nor (_20349_, _20348_, _03751_);
  nor (_20350_, _20348_, _04616_);
  nor (_20352_, _04615_, _20342_);
  or (_20353_, _20352_, _20350_);
  and (_20354_, _20353_, _04630_);
  nor (_20355_, _13234_, _09215_);
  nor (_20356_, _20355_, _20343_);
  nor (_20357_, _20356_, _04630_);
  or (_20358_, _20357_, _20354_);
  and (_20359_, _20358_, _04537_);
  nor (_20360_, _06013_, _09215_);
  nor (_20361_, _20360_, _20343_);
  nor (_20363_, _20361_, _04537_);
  nor (_20364_, _20363_, _20359_);
  nor (_20365_, _20364_, _03750_);
  or (_20366_, _20365_, _07544_);
  nor (_20367_, _20366_, _20349_);
  and (_20368_, _20361_, _07544_);
  nor (_20369_, _20368_, _20367_);
  nor (_20370_, _20369_, _04678_);
  and (_20371_, _06933_, _05411_);
  nor (_20372_, _20343_, _04679_);
  not (_20374_, _20372_);
  nor (_20375_, _20374_, _20371_);
  or (_20376_, _20375_, _07559_);
  nor (_20377_, _20376_, _20370_);
  nor (_20378_, _13326_, _09215_);
  nor (_20379_, _20378_, _20343_);
  nor (_20380_, _20379_, _03415_);
  or (_20381_, _20380_, _03839_);
  nor (_20382_, _20381_, _20377_);
  nor (_20383_, _20382_, _20346_);
  or (_20385_, _20383_, _03838_);
  and (_20386_, _13341_, _05411_);
  or (_20387_, _20343_, _04703_);
  nor (_20388_, _20387_, _20386_);
  nor (_20389_, _20388_, _03959_);
  and (_20390_, _20389_, _20385_);
  and (_20391_, _08695_, _05411_);
  nor (_20392_, _20391_, _20343_);
  nor (_20393_, _20392_, _04701_);
  nor (_20394_, _20393_, _20390_);
  nor (_20396_, _20394_, _03866_);
  nor (_20397_, _20343_, _08289_);
  not (_20398_, _20397_);
  nor (_20399_, _20345_, _04708_);
  and (_20400_, _20399_, _20398_);
  nor (_20401_, _20400_, _20396_);
  nor (_20402_, _20401_, _03967_);
  nor (_20403_, _20348_, _04706_);
  and (_20404_, _20403_, _20398_);
  nor (_20405_, _20404_, _03835_);
  not (_20407_, _20405_);
  nor (_20408_, _20407_, _20402_);
  nor (_20409_, _13340_, _09215_);
  or (_20410_, _20343_, _06532_);
  nor (_20411_, _20410_, _20409_);
  or (_20412_, _20411_, _03954_);
  nor (_20413_, _20412_, _20408_);
  nor (_20414_, _08694_, _09215_);
  nor (_20415_, _20414_, _20343_);
  nor (_20416_, _20415_, _06537_);
  or (_20418_, _20416_, _03703_);
  nor (_20419_, _20418_, _20413_);
  and (_20420_, _20356_, _03703_);
  or (_20421_, _20420_, _03701_);
  nor (_20422_, _20421_, _20419_);
  nor (_20423_, _13399_, _09215_);
  nor (_20424_, _20423_, _20343_);
  nor (_20425_, _20424_, _03702_);
  or (_20426_, _20425_, _20422_);
  or (_20427_, _20426_, _42912_);
  or (_20429_, _42908_, \oc8051_golden_model_1.TL0 [6]);
  and (_20430_, _20429_, _41654_);
  and (_43196_, _20430_, _20427_);
  not (_20431_, \oc8051_golden_model_1.TL1 [0]);
  nor (_20432_, _05516_, _20431_);
  nor (_20433_, _05652_, _09295_);
  nor (_20434_, _20433_, _20432_);
  and (_20435_, _20434_, _17066_);
  and (_20436_, _05516_, \oc8051_golden_model_1.ACC [0]);
  nor (_20437_, _20436_, _20432_);
  nor (_20439_, _20437_, _03751_);
  nor (_20440_, _20437_, _04616_);
  nor (_20441_, _04615_, _20431_);
  or (_20442_, _20441_, _20440_);
  and (_20443_, _20442_, _04630_);
  nor (_20444_, _20434_, _04630_);
  or (_20445_, _20444_, _20443_);
  and (_20446_, _20445_, _04537_);
  and (_20447_, _05428_, _04608_);
  nor (_20448_, _20447_, _20432_);
  nor (_20450_, _20448_, _04537_);
  nor (_20451_, _20450_, _20446_);
  nor (_20452_, _20451_, _03750_);
  or (_20453_, _20452_, _07544_);
  nor (_20454_, _20453_, _20439_);
  and (_20455_, _20448_, _07544_);
  nor (_20456_, _20455_, _20454_);
  nor (_20457_, _20456_, _04678_);
  nor (_20458_, _20432_, _04679_);
  or (_20459_, _06698_, _09295_);
  and (_20461_, _20459_, _20458_);
  nor (_20462_, _20461_, _20457_);
  and (_20463_, _20462_, _03415_);
  not (_20464_, _05516_);
  nor (_20465_, _12119_, _20464_);
  nor (_20466_, _20465_, _20432_);
  nor (_20467_, _20466_, _03415_);
  or (_20468_, _20467_, _20463_);
  and (_20469_, _20468_, _04694_);
  and (_20470_, _05516_, _06428_);
  nor (_20472_, _20470_, _20432_);
  nor (_20473_, _20472_, _04694_);
  or (_20474_, _20473_, _20469_);
  and (_20475_, _20474_, _04703_);
  and (_20476_, _12133_, _05516_);
  nor (_20477_, _20476_, _20432_);
  nor (_20478_, _20477_, _04703_);
  or (_20479_, _20478_, _20475_);
  and (_20480_, _20479_, _04701_);
  nor (_20481_, _10458_, _09295_);
  nor (_20483_, _20481_, _20432_);
  and (_20484_, _20436_, _05652_);
  or (_20485_, _20484_, _04701_);
  nor (_20486_, _20485_, _20483_);
  nor (_20487_, _20486_, _20480_);
  nor (_20488_, _20487_, _03866_);
  and (_20489_, _12013_, _05516_);
  or (_20490_, _20489_, _20432_);
  and (_20491_, _20490_, _03866_);
  or (_20492_, _20491_, _20488_);
  and (_20494_, _20492_, _04706_);
  nor (_20495_, _20484_, _20432_);
  nor (_20496_, _20495_, _04706_);
  or (_20497_, _20496_, _20494_);
  and (_20498_, _20497_, _06532_);
  nor (_20499_, _12132_, _20464_);
  nor (_20500_, _20499_, _20432_);
  nor (_20501_, _20500_, _06532_);
  or (_20502_, _20501_, _20498_);
  and (_20503_, _20502_, _06537_);
  nor (_20505_, _20483_, _06537_);
  nor (_20506_, _20505_, _17066_);
  not (_20507_, _20506_);
  nor (_20508_, _20507_, _20503_);
  nor (_20509_, _20508_, _20435_);
  or (_20510_, _20509_, _42912_);
  or (_20511_, _42908_, \oc8051_golden_model_1.TL1 [0]);
  and (_20512_, _20511_, _41654_);
  and (_43197_, _20512_, _20510_);
  not (_20513_, \oc8051_golden_model_1.TL1 [1]);
  nor (_20515_, _05516_, _20513_);
  nor (_20516_, _20515_, _04679_);
  or (_20517_, _06653_, _09295_);
  and (_20518_, _20517_, _20516_);
  not (_20519_, _20518_);
  and (_20520_, _05428_, _04813_);
  nor (_20521_, _20520_, _20515_);
  and (_20522_, _20521_, _07544_);
  and (_20523_, _05516_, \oc8051_golden_model_1.ACC [1]);
  nor (_20524_, _20523_, _20515_);
  nor (_20526_, _20524_, _04616_);
  nor (_20527_, _04615_, _20513_);
  or (_20528_, _20527_, _20526_);
  and (_20529_, _20528_, _04630_);
  nor (_20530_, _05516_, \oc8051_golden_model_1.TL1 [1]);
  and (_20531_, _12225_, _05428_);
  nor (_20532_, _20531_, _20530_);
  and (_20533_, _20532_, _03757_);
  or (_20534_, _20533_, _20529_);
  and (_20535_, _20534_, _04537_);
  nor (_20537_, _20521_, _04537_);
  nor (_20538_, _20537_, _20535_);
  nor (_20539_, _20538_, _03750_);
  nor (_20540_, _20524_, _03751_);
  nor (_20541_, _20540_, _07544_);
  not (_20542_, _20541_);
  nor (_20543_, _20542_, _20539_);
  nor (_20544_, _20543_, _20522_);
  nor (_20545_, _20544_, _04678_);
  nor (_20546_, _20545_, _07559_);
  and (_20548_, _20546_, _20519_);
  nor (_20549_, _12313_, _20464_);
  nor (_20550_, _20549_, _20515_);
  nor (_20551_, _20550_, _03415_);
  nor (_20552_, _20551_, _20548_);
  nor (_20553_, _20552_, _08854_);
  nor (_20554_, _12207_, _09295_);
  or (_20555_, _20554_, _04703_);
  and (_20556_, _05428_, _04515_);
  or (_20557_, _20556_, _04694_);
  and (_20559_, _20557_, _20555_);
  nor (_20560_, _20559_, _20530_);
  or (_20561_, _20560_, _03959_);
  nor (_20562_, _20561_, _20553_);
  nor (_20563_, _08710_, _09295_);
  nor (_20564_, _20563_, _20515_);
  and (_20565_, _20523_, _05603_);
  nor (_20566_, _20565_, _20564_);
  nor (_20567_, _20566_, _04701_);
  nor (_20568_, _20567_, _03866_);
  not (_20570_, _20568_);
  nor (_20571_, _20570_, _20562_);
  and (_20572_, _12206_, _05516_);
  or (_20573_, _20572_, _20515_);
  and (_20574_, _20573_, _03866_);
  or (_20575_, _20574_, _20571_);
  and (_20576_, _20575_, _04706_);
  nor (_20577_, _20565_, _20515_);
  nor (_20578_, _20577_, _04706_);
  or (_20579_, _20578_, _20576_);
  and (_20581_, _20579_, _06532_);
  nor (_20582_, _12205_, _20464_);
  or (_20583_, _20582_, _20515_);
  and (_20584_, _20583_, _03835_);
  or (_20585_, _20584_, _20581_);
  and (_20586_, _20585_, _06537_);
  nor (_20587_, _20564_, _06537_);
  or (_20588_, _20587_, _20586_);
  and (_20589_, _20588_, _03704_);
  and (_20590_, _20532_, _03703_);
  or (_20592_, _20590_, _20589_);
  and (_20593_, _20592_, _03702_);
  nor (_20594_, _20531_, _20515_);
  nor (_20595_, _20594_, _03702_);
  nor (_20596_, _20595_, _20593_);
  nand (_20597_, _20596_, _42908_);
  or (_20598_, _42908_, \oc8051_golden_model_1.TL1 [1]);
  and (_20599_, _20598_, _41654_);
  and (_43199_, _20599_, _20597_);
  not (_20600_, \oc8051_golden_model_1.TL1 [2]);
  nor (_20602_, _05516_, _20600_);
  and (_20603_, _05516_, \oc8051_golden_model_1.ACC [2]);
  nor (_20604_, _20603_, _20602_);
  nor (_20605_, _20604_, _03751_);
  nor (_20606_, _20604_, _04616_);
  nor (_20607_, _04615_, _20600_);
  or (_20608_, _20607_, _20606_);
  and (_20609_, _20608_, _04630_);
  nor (_20610_, _12427_, _09295_);
  nor (_20611_, _20610_, _20602_);
  nor (_20613_, _20611_, _04630_);
  or (_20614_, _20613_, _20609_);
  and (_20615_, _20614_, _04537_);
  nor (_20616_, _09295_, _05236_);
  nor (_20617_, _20616_, _20602_);
  nor (_20618_, _20617_, _04537_);
  nor (_20619_, _20618_, _20615_);
  nor (_20620_, _20619_, _03750_);
  or (_20621_, _20620_, _07544_);
  nor (_20622_, _20621_, _20605_);
  and (_20624_, _20617_, _07544_);
  nor (_20625_, _20624_, _20622_);
  nor (_20626_, _20625_, _04678_);
  nor (_20627_, _20602_, _04679_);
  or (_20628_, _06789_, _09295_);
  and (_20629_, _20628_, _20627_);
  or (_20630_, _20629_, _07559_);
  nor (_20631_, _20630_, _20626_);
  nor (_20632_, _12523_, _09295_);
  nor (_20633_, _20632_, _20602_);
  nor (_20635_, _20633_, _03415_);
  or (_20636_, _20635_, _08854_);
  or (_20637_, _20636_, _20631_);
  and (_20638_, _12537_, _05428_);
  or (_20639_, _20602_, _04703_);
  or (_20640_, _20639_, _20638_);
  and (_20641_, _05516_, _06457_);
  nor (_20642_, _20641_, _20602_);
  and (_20643_, _20642_, _03839_);
  nor (_20644_, _20643_, _03959_);
  and (_20646_, _20644_, _20640_);
  and (_20647_, _20646_, _20637_);
  and (_20648_, _08707_, _05516_);
  nor (_20649_, _20648_, _20602_);
  nor (_20650_, _20649_, _04701_);
  nor (_20651_, _20650_, _20647_);
  nor (_20652_, _20651_, _03866_);
  nor (_20653_, _20602_, _05700_);
  not (_20654_, _20653_);
  nor (_20655_, _20642_, _04708_);
  and (_20657_, _20655_, _20654_);
  nor (_20658_, _20657_, _20652_);
  nor (_20659_, _20658_, _03967_);
  nor (_20660_, _20604_, _04706_);
  and (_20661_, _20660_, _20654_);
  or (_20662_, _20661_, _20659_);
  and (_20663_, _20662_, _06532_);
  nor (_20664_, _12536_, _20464_);
  nor (_20665_, _20664_, _20602_);
  nor (_20666_, _20665_, _06532_);
  or (_20668_, _20666_, _20663_);
  and (_20669_, _20668_, _06537_);
  nor (_20670_, _08706_, _09295_);
  nor (_20671_, _20670_, _20602_);
  nor (_20672_, _20671_, _06537_);
  or (_20673_, _20672_, _03703_);
  nor (_20674_, _20673_, _20669_);
  and (_20675_, _20611_, _03703_);
  or (_20676_, _20675_, _03701_);
  nor (_20677_, _20676_, _20674_);
  and (_20679_, _12596_, _05516_);
  nor (_20680_, _20679_, _20602_);
  nor (_20681_, _20680_, _03702_);
  or (_20682_, _20681_, _20677_);
  or (_20683_, _20682_, _42912_);
  or (_20684_, _42908_, \oc8051_golden_model_1.TL1 [2]);
  and (_20685_, _20684_, _41654_);
  and (_43200_, _20685_, _20683_);
  and (_20686_, _20464_, \oc8051_golden_model_1.TL1 [3]);
  nor (_20687_, _12610_, _09295_);
  or (_20689_, _20687_, _20686_);
  or (_20690_, _20689_, _04630_);
  and (_20691_, _05516_, \oc8051_golden_model_1.ACC [3]);
  or (_20692_, _20691_, _20686_);
  and (_20693_, _20692_, _04615_);
  and (_20694_, _04616_, \oc8051_golden_model_1.TL1 [3]);
  or (_20695_, _20694_, _03757_);
  or (_20696_, _20695_, _20693_);
  and (_20697_, _20696_, _04537_);
  and (_20698_, _20697_, _20690_);
  nor (_20700_, _09295_, _05050_);
  or (_20701_, _20700_, _20686_);
  and (_20702_, _20701_, _03755_);
  or (_20703_, _20702_, _20698_);
  and (_20704_, _20703_, _03751_);
  and (_20705_, _20692_, _03750_);
  or (_20706_, _20705_, _07544_);
  or (_20707_, _20706_, _20704_);
  or (_20708_, _20701_, _06994_);
  and (_20709_, _20708_, _20707_);
  or (_20711_, _20709_, _04678_);
  and (_20712_, _06937_, _05516_);
  or (_20713_, _20686_, _04679_);
  or (_20714_, _20713_, _20712_);
  and (_20715_, _20714_, _03415_);
  and (_20716_, _20715_, _20711_);
  nor (_20717_, _12724_, _09295_);
  or (_20718_, _20717_, _20686_);
  and (_20719_, _20718_, _07559_);
  or (_20720_, _20719_, _08854_);
  or (_20722_, _20720_, _20716_);
  and (_20723_, _12738_, _05428_);
  or (_20724_, _20686_, _04703_);
  or (_20725_, _20724_, _20723_);
  and (_20726_, _05516_, _06415_);
  or (_20727_, _20726_, _20686_);
  or (_20728_, _20727_, _04694_);
  and (_20729_, _20728_, _04701_);
  and (_20730_, _20729_, _20725_);
  and (_20731_, _20730_, _20722_);
  and (_20733_, _10455_, _05516_);
  or (_20734_, _20733_, _20686_);
  and (_20735_, _20734_, _03959_);
  or (_20736_, _20735_, _20731_);
  and (_20737_, _20736_, _04708_);
  or (_20738_, _20686_, _05554_);
  and (_20739_, _20727_, _03866_);
  and (_20740_, _20739_, _20738_);
  or (_20741_, _20740_, _20737_);
  and (_20742_, _20741_, _04706_);
  and (_20744_, _20692_, _03967_);
  and (_20745_, _20744_, _20738_);
  or (_20746_, _20745_, _03835_);
  or (_20747_, _20746_, _20742_);
  nor (_20748_, _12737_, _09295_);
  or (_20749_, _20686_, _06532_);
  or (_20750_, _20749_, _20748_);
  and (_20751_, _20750_, _06537_);
  and (_20752_, _20751_, _20747_);
  nor (_20753_, _08701_, _09295_);
  or (_20755_, _20753_, _20686_);
  and (_20756_, _20755_, _03954_);
  or (_20757_, _20756_, _03703_);
  or (_20758_, _20757_, _20752_);
  or (_20759_, _20689_, _03704_);
  and (_20760_, _20759_, _03702_);
  and (_20761_, _20760_, _20758_);
  and (_20762_, _12792_, _05516_);
  or (_20763_, _20762_, _20686_);
  and (_20764_, _20763_, _03701_);
  or (_20766_, _20764_, _20761_);
  or (_20767_, _20766_, _42912_);
  or (_20768_, _42908_, \oc8051_golden_model_1.TL1 [3]);
  and (_20769_, _20768_, _41654_);
  and (_43201_, _20769_, _20767_);
  not (_20770_, \oc8051_golden_model_1.TL1 [4]);
  nor (_20771_, _05516_, _20770_);
  and (_20772_, _06422_, _05516_);
  nor (_20773_, _20772_, _20771_);
  and (_20774_, _20773_, _03839_);
  nor (_20776_, _05898_, _09295_);
  nor (_20777_, _20776_, _20771_);
  and (_20778_, _20777_, _07544_);
  and (_20779_, _05516_, \oc8051_golden_model_1.ACC [4]);
  nor (_20780_, _20779_, _20771_);
  nor (_20781_, _20780_, _04616_);
  nor (_20782_, _04615_, _20770_);
  or (_20783_, _20782_, _20781_);
  and (_20784_, _20783_, _04630_);
  nor (_20785_, _12828_, _09295_);
  nor (_20787_, _20785_, _20771_);
  nor (_20788_, _20787_, _04630_);
  or (_20789_, _20788_, _20784_);
  and (_20790_, _20789_, _04537_);
  nor (_20791_, _20777_, _04537_);
  nor (_20792_, _20791_, _20790_);
  nor (_20793_, _20792_, _03750_);
  nor (_20794_, _20780_, _03751_);
  nor (_20795_, _20794_, _07544_);
  not (_20796_, _20795_);
  nor (_20798_, _20796_, _20793_);
  nor (_20799_, _20798_, _20778_);
  nor (_20800_, _20799_, _04678_);
  nor (_20801_, _20771_, _04679_);
  or (_20802_, _06881_, _09295_);
  and (_20803_, _20802_, _20801_);
  or (_20804_, _20803_, _07559_);
  nor (_20805_, _20804_, _20800_);
  nor (_20806_, _12919_, _20464_);
  nor (_20807_, _20806_, _20771_);
  nor (_20809_, _20807_, _03415_);
  or (_20810_, _20809_, _03839_);
  nor (_20811_, _20810_, _20805_);
  nor (_20812_, _20811_, _20774_);
  or (_20813_, _20812_, _03838_);
  and (_20814_, _12933_, _05516_);
  or (_20815_, _20814_, _20771_);
  or (_20816_, _20815_, _04703_);
  and (_20817_, _20816_, _04701_);
  and (_20818_, _20817_, _20813_);
  and (_20820_, _08700_, _05516_);
  nor (_20821_, _20820_, _20771_);
  nor (_20822_, _20821_, _04701_);
  nor (_20823_, _20822_, _20818_);
  nor (_20824_, _20823_, _03866_);
  nor (_20825_, _20771_, _08303_);
  not (_20826_, _20825_);
  nor (_20827_, _20773_, _04708_);
  and (_20828_, _20827_, _20826_);
  nor (_20829_, _20828_, _20824_);
  nor (_20831_, _20829_, _03967_);
  nor (_20832_, _20780_, _04706_);
  and (_20833_, _20832_, _20826_);
  or (_20834_, _20833_, _20831_);
  and (_20835_, _20834_, _06532_);
  nor (_20836_, _12931_, _20464_);
  nor (_20837_, _20836_, _20771_);
  nor (_20838_, _20837_, _06532_);
  or (_20839_, _20838_, _20835_);
  and (_20840_, _20839_, _06537_);
  nor (_20842_, _08699_, _09295_);
  nor (_20843_, _20842_, _20771_);
  nor (_20844_, _20843_, _06537_);
  or (_20845_, _20844_, _03703_);
  nor (_20846_, _20845_, _20840_);
  and (_20847_, _20787_, _03703_);
  or (_20848_, _20847_, _03701_);
  nor (_20849_, _20848_, _20846_);
  and (_20850_, _12991_, _05516_);
  nor (_20851_, _20850_, _20771_);
  nor (_20853_, _20851_, _03702_);
  or (_20854_, _20853_, _20849_);
  or (_20855_, _20854_, _42912_);
  or (_20856_, _42908_, \oc8051_golden_model_1.TL1 [4]);
  and (_20857_, _20856_, _41654_);
  and (_43202_, _20857_, _20855_);
  and (_20858_, _20464_, \oc8051_golden_model_1.TL1 [5]);
  nor (_20859_, _13025_, _09295_);
  or (_20860_, _20859_, _20858_);
  or (_20861_, _20860_, _04630_);
  and (_20863_, _05516_, \oc8051_golden_model_1.ACC [5]);
  or (_20864_, _20863_, _20858_);
  and (_20865_, _20864_, _04615_);
  and (_20866_, _04616_, \oc8051_golden_model_1.TL1 [5]);
  or (_20867_, _20866_, _03757_);
  or (_20868_, _20867_, _20865_);
  and (_20869_, _20868_, _04537_);
  and (_20870_, _20869_, _20861_);
  nor (_20871_, _05799_, _09295_);
  or (_20872_, _20871_, _20858_);
  and (_20874_, _20872_, _03755_);
  or (_20875_, _20874_, _20870_);
  and (_20876_, _20875_, _03751_);
  and (_20877_, _20864_, _03750_);
  or (_20878_, _20877_, _07544_);
  or (_20879_, _20878_, _20876_);
  or (_20880_, _20872_, _06994_);
  and (_20881_, _20880_, _20879_);
  or (_20882_, _20881_, _04678_);
  and (_20883_, _06941_, _05516_);
  or (_20885_, _20858_, _04679_);
  or (_20886_, _20885_, _20883_);
  and (_20887_, _20886_, _03415_);
  and (_20888_, _20887_, _20882_);
  nor (_20889_, _13118_, _09295_);
  or (_20890_, _20889_, _20858_);
  and (_20891_, _20890_, _07559_);
  or (_20892_, _20891_, _08854_);
  or (_20893_, _20892_, _20888_);
  and (_20894_, _13133_, _05428_);
  or (_20896_, _20858_, _04703_);
  or (_20897_, _20896_, _20894_);
  and (_20898_, _06371_, _05516_);
  or (_20899_, _20898_, _20858_);
  or (_20900_, _20899_, _04694_);
  and (_20901_, _20900_, _04701_);
  and (_20902_, _20901_, _20897_);
  and (_20903_, _20902_, _20893_);
  and (_20904_, _10451_, _05516_);
  or (_20905_, _20904_, _20858_);
  and (_20907_, _20905_, _03959_);
  or (_20908_, _20907_, _20903_);
  and (_20909_, _20908_, _04708_);
  or (_20910_, _20858_, _08302_);
  and (_20911_, _20899_, _03866_);
  and (_20912_, _20911_, _20910_);
  or (_20913_, _20912_, _20909_);
  and (_20914_, _20913_, _04706_);
  and (_20915_, _20864_, _03967_);
  and (_20916_, _20915_, _20910_);
  or (_20918_, _20916_, _03835_);
  or (_20919_, _20918_, _20914_);
  nor (_20920_, _13131_, _09295_);
  or (_20921_, _20858_, _06532_);
  or (_20922_, _20921_, _20920_);
  and (_20923_, _20922_, _06537_);
  and (_20924_, _20923_, _20919_);
  nor (_20925_, _08697_, _09295_);
  or (_20926_, _20925_, _20858_);
  and (_20927_, _20926_, _03954_);
  or (_20928_, _20927_, _20924_);
  and (_20929_, _20928_, _03704_);
  and (_20930_, _20860_, _03703_);
  or (_20931_, _20930_, _03701_);
  or (_20932_, _20931_, _20929_);
  and (_20933_, _13193_, _05516_);
  or (_20934_, _20933_, _20858_);
  or (_20935_, _20934_, _03702_);
  and (_20936_, _20935_, _20932_);
  or (_20937_, _20936_, _42912_);
  or (_20939_, _42908_, \oc8051_golden_model_1.TL1 [5]);
  and (_20940_, _20939_, _41654_);
  and (_43203_, _20940_, _20937_);
  not (_20941_, \oc8051_golden_model_1.TL1 [6]);
  nor (_20942_, _05516_, _20941_);
  and (_20943_, _13333_, _05516_);
  nor (_20944_, _20943_, _20942_);
  and (_20945_, _20944_, _03839_);
  nor (_20946_, _06013_, _09295_);
  nor (_20947_, _20946_, _20942_);
  and (_20949_, _20947_, _07544_);
  and (_20950_, _05516_, \oc8051_golden_model_1.ACC [6]);
  nor (_20951_, _20950_, _20942_);
  nor (_20952_, _20951_, _04616_);
  nor (_20953_, _04615_, _20941_);
  or (_20954_, _20953_, _20952_);
  and (_20955_, _20954_, _04630_);
  nor (_20956_, _13234_, _09295_);
  nor (_20957_, _20956_, _20942_);
  nor (_20958_, _20957_, _04630_);
  or (_20960_, _20958_, _20955_);
  and (_20961_, _20960_, _04537_);
  nor (_20962_, _20947_, _04537_);
  nor (_20963_, _20962_, _20961_);
  nor (_20964_, _20963_, _03750_);
  nor (_20965_, _20951_, _03751_);
  nor (_20966_, _20965_, _07544_);
  not (_20967_, _20966_);
  nor (_20968_, _20967_, _20964_);
  nor (_20969_, _20968_, _20949_);
  nor (_20970_, _20969_, _04678_);
  nor (_20971_, _20942_, _04679_);
  or (_20972_, _06607_, _09295_);
  and (_20973_, _20972_, _20971_);
  or (_20974_, _20973_, _07559_);
  nor (_20975_, _20974_, _20970_);
  nor (_20976_, _13326_, _20464_);
  nor (_20977_, _20976_, _20942_);
  nor (_20978_, _20977_, _03415_);
  or (_20979_, _20978_, _03839_);
  nor (_20981_, _20979_, _20975_);
  nor (_20982_, _20981_, _20945_);
  or (_20983_, _20982_, _03838_);
  and (_20984_, _13341_, _05516_);
  or (_20985_, _20984_, _20942_);
  or (_20986_, _20985_, _04703_);
  and (_20987_, _20986_, _04701_);
  and (_20988_, _20987_, _20983_);
  and (_20989_, _08695_, _05516_);
  nor (_20990_, _20989_, _20942_);
  nor (_20991_, _20990_, _04701_);
  nor (_20992_, _20991_, _20988_);
  nor (_20993_, _20992_, _03866_);
  nor (_20994_, _20942_, _08289_);
  not (_20995_, _20994_);
  nor (_20996_, _20944_, _04708_);
  and (_20997_, _20996_, _20995_);
  nor (_20998_, _20997_, _20993_);
  nor (_20999_, _20998_, _03967_);
  nor (_21000_, _20951_, _04706_);
  and (_21002_, _21000_, _20995_);
  nor (_21003_, _21002_, _03835_);
  not (_21004_, _21003_);
  nor (_21005_, _21004_, _20999_);
  or (_21006_, _13340_, _09295_);
  nor (_21007_, _20942_, _06532_);
  and (_21008_, _21007_, _21006_);
  or (_21009_, _21008_, _03954_);
  nor (_21010_, _21009_, _21005_);
  nor (_21011_, _08694_, _09295_);
  nor (_21013_, _21011_, _20942_);
  nor (_21014_, _21013_, _06537_);
  or (_21015_, _21014_, _03703_);
  nor (_21016_, _21015_, _21010_);
  and (_21017_, _20957_, _03703_);
  or (_21018_, _21017_, _03701_);
  nor (_21019_, _21018_, _21016_);
  nor (_21020_, _13399_, _20464_);
  nor (_21021_, _21020_, _20942_);
  nor (_21022_, _21021_, _03702_);
  or (_21023_, _21022_, _21019_);
  or (_21024_, _21023_, _42912_);
  or (_21025_, _42908_, \oc8051_golden_model_1.TL1 [6]);
  and (_21026_, _21025_, _41654_);
  and (_43204_, _21026_, _21024_);
  not (_21027_, \oc8051_golden_model_1.TH0 [0]);
  nor (_21028_, _05426_, _21027_);
  nor (_21029_, _05652_, _09375_);
  nor (_21030_, _21029_, _21028_);
  and (_21031_, _21030_, _17066_);
  and (_21033_, _05426_, \oc8051_golden_model_1.ACC [0]);
  nor (_21034_, _21033_, _21028_);
  nor (_21035_, _21034_, _03751_);
  nor (_21036_, _21035_, _07544_);
  nor (_21037_, _21030_, _04630_);
  nor (_21038_, _04615_, _21027_);
  nor (_21039_, _21034_, _04616_);
  nor (_21040_, _21039_, _21038_);
  nor (_21041_, _21040_, _03757_);
  or (_21042_, _21041_, _03755_);
  nor (_21044_, _21042_, _21037_);
  or (_21045_, _21044_, _03750_);
  and (_21046_, _21045_, _21036_);
  and (_21047_, _05426_, _04608_);
  or (_21048_, _21028_, _19847_);
  nor (_21049_, _21048_, _21047_);
  nor (_21050_, _21049_, _21046_);
  nor (_21051_, _21050_, _04678_);
  and (_21052_, _06935_, _05426_);
  nor (_21053_, _21028_, _04679_);
  not (_21054_, _21053_);
  nor (_21055_, _21054_, _21052_);
  nor (_21056_, _21055_, _21051_);
  and (_21057_, _21056_, _03415_);
  nor (_21058_, _12119_, _09375_);
  nor (_21059_, _21058_, _21028_);
  nor (_21060_, _21059_, _03415_);
  or (_21061_, _21060_, _21057_);
  and (_21062_, _21061_, _04694_);
  and (_21063_, _05426_, _06428_);
  nor (_21065_, _21063_, _21028_);
  nor (_21066_, _21065_, _04694_);
  or (_21067_, _21066_, _21062_);
  and (_21068_, _21067_, _04703_);
  and (_21069_, _12133_, _05426_);
  nor (_21070_, _21069_, _21028_);
  nor (_21071_, _21070_, _04703_);
  or (_21072_, _21071_, _21068_);
  and (_21073_, _21072_, _04701_);
  nor (_21074_, _10458_, _09375_);
  nor (_21076_, _21074_, _21028_);
  not (_21077_, _21076_);
  and (_21078_, _08712_, _05426_);
  nor (_21079_, _21078_, _04701_);
  and (_21080_, _21079_, _21077_);
  nor (_21081_, _21080_, _21073_);
  nor (_21082_, _21081_, _03866_);
  and (_21083_, _12013_, _05426_);
  or (_21084_, _21083_, _21028_);
  and (_21085_, _21084_, _03866_);
  or (_21086_, _21085_, _21082_);
  and (_21087_, _21086_, _04706_);
  nor (_21088_, _21078_, _21028_);
  nor (_21089_, _21088_, _04706_);
  or (_21090_, _21089_, _21087_);
  and (_21091_, _21090_, _06532_);
  nor (_21092_, _12132_, _09375_);
  nor (_21093_, _21092_, _21028_);
  nor (_21094_, _21093_, _06532_);
  or (_21095_, _21094_, _21091_);
  and (_21097_, _21095_, _06537_);
  nor (_21098_, _21076_, _06537_);
  nor (_21099_, _21098_, _17066_);
  not (_21100_, _21099_);
  nor (_21101_, _21100_, _21097_);
  nor (_21102_, _21101_, _21031_);
  or (_21103_, _21102_, _42912_);
  or (_21104_, _42908_, \oc8051_golden_model_1.TH0 [0]);
  and (_21105_, _21104_, _41654_);
  and (_43207_, _21105_, _21103_);
  and (_21107_, _06934_, _05426_);
  not (_21108_, \oc8051_golden_model_1.TH0 [1]);
  nor (_21109_, _05426_, _21108_);
  nor (_21110_, _21109_, _04679_);
  not (_21111_, _21110_);
  nor (_21112_, _21111_, _21107_);
  not (_21113_, _21112_);
  and (_21114_, _05426_, \oc8051_golden_model_1.ACC [1]);
  nor (_21115_, _21114_, _21109_);
  nor (_21116_, _21115_, _03751_);
  nor (_21117_, _21115_, _04616_);
  nor (_21118_, _04615_, _21108_);
  or (_21119_, _21118_, _21117_);
  and (_21120_, _21119_, _04630_);
  nor (_21121_, _05426_, \oc8051_golden_model_1.TH0 [1]);
  and (_21122_, _12225_, _05426_);
  nor (_21123_, _21122_, _21121_);
  and (_21124_, _21123_, _03757_);
  or (_21125_, _21124_, _21120_);
  and (_21126_, _21125_, _04537_);
  and (_21128_, _05426_, _04813_);
  nor (_21129_, _21128_, _21109_);
  nor (_21130_, _21129_, _04537_);
  nor (_21131_, _21130_, _21126_);
  nor (_21132_, _21131_, _03750_);
  or (_21133_, _21132_, _07544_);
  nor (_21134_, _21133_, _21116_);
  and (_21135_, _21129_, _07544_);
  nor (_21136_, _21135_, _21134_);
  nor (_21137_, _21136_, _04678_);
  nor (_21139_, _21137_, _07559_);
  and (_21140_, _21139_, _21113_);
  and (_21141_, _12313_, _05426_);
  or (_21142_, _21141_, _03415_);
  nor (_21143_, _21142_, _21121_);
  nor (_21144_, _21143_, _21140_);
  nor (_21145_, _21144_, _08854_);
  nor (_21146_, _12207_, _09375_);
  or (_21147_, _21146_, _04703_);
  and (_21148_, _05426_, _04515_);
  or (_21149_, _21148_, _04694_);
  and (_21150_, _21149_, _21147_);
  nor (_21151_, _21150_, _21121_);
  or (_21152_, _21151_, _03959_);
  nor (_21153_, _21152_, _21145_);
  nor (_21154_, _08710_, _09375_);
  nor (_21155_, _21154_, _21109_);
  and (_21156_, _08709_, _05426_);
  nor (_21157_, _21156_, _21155_);
  nor (_21158_, _21157_, _04701_);
  nor (_21160_, _21158_, _03866_);
  not (_21161_, _21160_);
  nor (_21162_, _21161_, _21153_);
  and (_21163_, _12206_, _05426_);
  or (_21164_, _21163_, _21109_);
  and (_21165_, _21164_, _03866_);
  or (_21166_, _21165_, _21162_);
  and (_21167_, _21166_, _04706_);
  nor (_21168_, _21156_, _21109_);
  nor (_21169_, _21168_, _04706_);
  or (_21171_, _21169_, _21167_);
  and (_21172_, _21171_, _06532_);
  nor (_21173_, _12205_, _09375_);
  or (_21174_, _21173_, _21109_);
  and (_21175_, _21174_, _03835_);
  or (_21176_, _21175_, _21172_);
  and (_21177_, _21176_, _06537_);
  nor (_21178_, _21155_, _06537_);
  or (_21179_, _21178_, _21177_);
  and (_21180_, _21179_, _03704_);
  and (_21181_, _21123_, _03703_);
  or (_21182_, _21181_, _21180_);
  and (_21183_, _21182_, _03702_);
  nor (_21184_, _21122_, _21109_);
  nor (_21185_, _21184_, _03702_);
  nor (_21186_, _21185_, _21183_);
  nand (_21187_, _21186_, _42908_);
  or (_21188_, _42908_, \oc8051_golden_model_1.TH0 [1]);
  and (_21189_, _21188_, _41654_);
  and (_43208_, _21189_, _21187_);
  not (_21191_, \oc8051_golden_model_1.TH0 [2]);
  nor (_21192_, _05426_, _21191_);
  nor (_21193_, _09375_, _05236_);
  nor (_21194_, _21193_, _21192_);
  and (_21195_, _21194_, _07544_);
  and (_21196_, _05426_, \oc8051_golden_model_1.ACC [2]);
  nor (_21197_, _21196_, _21192_);
  nor (_21198_, _21197_, _03751_);
  nor (_21199_, _21197_, _04616_);
  nor (_21200_, _04615_, _21191_);
  or (_21202_, _21200_, _21199_);
  and (_21203_, _21202_, _04630_);
  nor (_21204_, _12427_, _09375_);
  nor (_21205_, _21204_, _21192_);
  nor (_21206_, _21205_, _04630_);
  or (_21207_, _21206_, _21203_);
  and (_21208_, _21207_, _04537_);
  nor (_21209_, _21194_, _04537_);
  nor (_21210_, _21209_, _21208_);
  nor (_21211_, _21210_, _03750_);
  or (_21212_, _21211_, _07544_);
  nor (_21213_, _21212_, _21198_);
  nor (_21214_, _21213_, _21195_);
  nor (_21215_, _21214_, _04678_);
  and (_21216_, _06938_, _05426_);
  nor (_21217_, _21192_, _04679_);
  not (_21218_, _21217_);
  nor (_21219_, _21218_, _21216_);
  nor (_21220_, _21219_, _07559_);
  not (_21221_, _21220_);
  nor (_21223_, _21221_, _21215_);
  nor (_21224_, _12523_, _09375_);
  nor (_21225_, _21224_, _21192_);
  nor (_21226_, _21225_, _03415_);
  or (_21227_, _21226_, _08854_);
  or (_21228_, _21227_, _21223_);
  and (_21229_, _12537_, _05426_);
  or (_21230_, _21192_, _04703_);
  nor (_21231_, _21230_, _21229_);
  and (_21232_, _05426_, _06457_);
  nor (_21234_, _21232_, _21192_);
  and (_21235_, _21234_, _03839_);
  or (_21236_, _21235_, _03959_);
  nor (_21237_, _21236_, _21231_);
  and (_21238_, _21237_, _21228_);
  and (_21239_, _08707_, _05426_);
  nor (_21240_, _21239_, _21192_);
  nor (_21241_, _21240_, _04701_);
  nor (_21242_, _21241_, _21238_);
  nor (_21243_, _21242_, _03866_);
  nor (_21244_, _21192_, _05700_);
  not (_21245_, _21244_);
  nor (_21246_, _21234_, _04708_);
  and (_21247_, _21246_, _21245_);
  nor (_21248_, _21247_, _21243_);
  nor (_21249_, _21248_, _03967_);
  nor (_21250_, _21197_, _04706_);
  and (_21251_, _21250_, _21245_);
  or (_21252_, _21251_, _21249_);
  and (_21253_, _21252_, _06532_);
  nor (_21255_, _12536_, _09375_);
  nor (_21256_, _21255_, _21192_);
  nor (_21257_, _21256_, _06532_);
  or (_21258_, _21257_, _21253_);
  and (_21259_, _21258_, _06537_);
  nor (_21260_, _08706_, _09375_);
  nor (_21261_, _21260_, _21192_);
  nor (_21262_, _21261_, _06537_);
  or (_21263_, _21262_, _03703_);
  nor (_21264_, _21263_, _21259_);
  and (_21266_, _21205_, _03703_);
  or (_21267_, _21266_, _03701_);
  nor (_21268_, _21267_, _21264_);
  and (_21269_, _12596_, _05426_);
  nor (_21270_, _21269_, _21192_);
  nor (_21271_, _21270_, _03702_);
  or (_21272_, _21271_, _21268_);
  or (_21273_, _21272_, _42912_);
  or (_21274_, _42908_, \oc8051_golden_model_1.TH0 [2]);
  and (_21275_, _21274_, _41654_);
  and (_43209_, _21275_, _21273_);
  and (_21276_, _09375_, \oc8051_golden_model_1.TH0 [3]);
  nor (_21277_, _12610_, _09375_);
  or (_21278_, _21277_, _21276_);
  or (_21279_, _21278_, _04630_);
  and (_21280_, _05426_, \oc8051_golden_model_1.ACC [3]);
  or (_21281_, _21280_, _21276_);
  and (_21282_, _21281_, _04615_);
  and (_21283_, _04616_, \oc8051_golden_model_1.TH0 [3]);
  or (_21284_, _21283_, _03757_);
  or (_21286_, _21284_, _21282_);
  and (_21287_, _21286_, _04537_);
  and (_21288_, _21287_, _21279_);
  nor (_21289_, _09375_, _05050_);
  or (_21290_, _21289_, _21276_);
  and (_21291_, _21290_, _03755_);
  or (_21292_, _21291_, _21288_);
  and (_21293_, _21292_, _03751_);
  and (_21294_, _21281_, _03750_);
  or (_21295_, _21294_, _07544_);
  or (_21297_, _21295_, _21293_);
  or (_21298_, _21290_, _06994_);
  and (_21299_, _21298_, _21297_);
  or (_21300_, _21299_, _04678_);
  and (_21301_, _06937_, _05426_);
  or (_21302_, _21276_, _04679_);
  or (_21303_, _21302_, _21301_);
  and (_21304_, _21303_, _03415_);
  and (_21305_, _21304_, _21300_);
  nor (_21306_, _12724_, _09375_);
  or (_21307_, _21306_, _21276_);
  and (_21308_, _21307_, _07559_);
  or (_21309_, _21308_, _08854_);
  or (_21310_, _21309_, _21305_);
  and (_21311_, _12738_, _05426_);
  or (_21312_, _21276_, _04703_);
  or (_21313_, _21312_, _21311_);
  and (_21314_, _05426_, _06415_);
  or (_21315_, _21314_, _21276_);
  or (_21316_, _21315_, _04694_);
  and (_21318_, _21316_, _04701_);
  and (_21319_, _21318_, _21313_);
  and (_21320_, _21319_, _21310_);
  and (_21321_, _10455_, _05426_);
  or (_21322_, _21321_, _21276_);
  and (_21323_, _21322_, _03959_);
  or (_21324_, _21323_, _21320_);
  and (_21325_, _21324_, _04708_);
  or (_21326_, _21276_, _05554_);
  and (_21327_, _21315_, _03866_);
  and (_21329_, _21327_, _21326_);
  or (_21330_, _21329_, _21325_);
  and (_21331_, _21330_, _04706_);
  and (_21332_, _21281_, _03967_);
  and (_21333_, _21332_, _21326_);
  or (_21334_, _21333_, _03835_);
  or (_21335_, _21334_, _21331_);
  nor (_21336_, _12737_, _09375_);
  or (_21337_, _21276_, _06532_);
  or (_21338_, _21337_, _21336_);
  and (_21340_, _21338_, _06537_);
  and (_21341_, _21340_, _21335_);
  nor (_21342_, _08701_, _09375_);
  or (_21343_, _21342_, _21276_);
  and (_21344_, _21343_, _03954_);
  or (_21345_, _21344_, _03703_);
  or (_21346_, _21345_, _21341_);
  or (_21347_, _21278_, _03704_);
  and (_21348_, _21347_, _03702_);
  and (_21349_, _21348_, _21346_);
  and (_21350_, _12792_, _05426_);
  or (_21351_, _21350_, _21276_);
  and (_21352_, _21351_, _03701_);
  or (_21353_, _21352_, _21349_);
  or (_21354_, _21353_, _42912_);
  or (_21355_, _42908_, \oc8051_golden_model_1.TH0 [3]);
  and (_21356_, _21355_, _41654_);
  and (_43210_, _21356_, _21354_);
  not (_21357_, \oc8051_golden_model_1.TH0 [4]);
  nor (_21358_, _05426_, _21357_);
  and (_21360_, _06422_, _05426_);
  nor (_21361_, _21360_, _21358_);
  and (_21362_, _21361_, _03839_);
  and (_21363_, _05426_, \oc8051_golden_model_1.ACC [4]);
  nor (_21364_, _21363_, _21358_);
  nor (_21365_, _21364_, _03751_);
  nor (_21366_, _21364_, _04616_);
  nor (_21367_, _04615_, _21357_);
  or (_21368_, _21367_, _21366_);
  and (_21369_, _21368_, _04630_);
  nor (_21371_, _12828_, _09375_);
  nor (_21372_, _21371_, _21358_);
  nor (_21373_, _21372_, _04630_);
  or (_21374_, _21373_, _21369_);
  and (_21375_, _21374_, _04537_);
  nor (_21376_, _05898_, _09375_);
  nor (_21377_, _21376_, _21358_);
  nor (_21378_, _21377_, _04537_);
  nor (_21379_, _21378_, _21375_);
  nor (_21380_, _21379_, _03750_);
  or (_21382_, _21380_, _07544_);
  nor (_21383_, _21382_, _21365_);
  and (_21384_, _21377_, _07544_);
  nor (_21385_, _21384_, _21383_);
  nor (_21386_, _21385_, _04678_);
  and (_21387_, _06942_, _05426_);
  nor (_21388_, _21358_, _04679_);
  not (_21389_, _21388_);
  nor (_21390_, _21389_, _21387_);
  or (_21391_, _21390_, _07559_);
  nor (_21393_, _21391_, _21386_);
  nor (_21394_, _12919_, _09375_);
  nor (_21395_, _21394_, _21358_);
  nor (_21396_, _21395_, _03415_);
  or (_21397_, _21396_, _03839_);
  nor (_21398_, _21397_, _21393_);
  nor (_21399_, _21398_, _21362_);
  or (_21400_, _21399_, _03838_);
  and (_21401_, _12933_, _05426_);
  or (_21402_, _21401_, _21358_);
  or (_21405_, _21402_, _04703_);
  and (_21406_, _21405_, _04701_);
  and (_21407_, _21406_, _21400_);
  and (_21408_, _08700_, _05426_);
  nor (_21409_, _21408_, _21358_);
  nor (_21410_, _21409_, _04701_);
  nor (_21411_, _21410_, _21407_);
  nor (_21412_, _21411_, _03866_);
  nor (_21413_, _21358_, _08303_);
  not (_21414_, _21413_);
  nor (_21417_, _21361_, _04708_);
  and (_21418_, _21417_, _21414_);
  nor (_21419_, _21418_, _21412_);
  nor (_21420_, _21419_, _03967_);
  nor (_21421_, _21364_, _04706_);
  and (_21422_, _21421_, _21414_);
  or (_21423_, _21422_, _21420_);
  and (_21424_, _21423_, _06532_);
  nor (_21425_, _12931_, _09375_);
  nor (_21426_, _21425_, _21358_);
  nor (_21429_, _21426_, _06532_);
  or (_21430_, _21429_, _21424_);
  and (_21431_, _21430_, _06537_);
  nor (_21432_, _08699_, _09375_);
  nor (_21433_, _21432_, _21358_);
  nor (_21434_, _21433_, _06537_);
  or (_21435_, _21434_, _03703_);
  nor (_21436_, _21435_, _21431_);
  and (_21437_, _21372_, _03703_);
  or (_21438_, _21437_, _03701_);
  nor (_21440_, _21438_, _21436_);
  and (_21441_, _12991_, _05426_);
  nor (_21442_, _21441_, _21358_);
  nor (_21443_, _21442_, _03702_);
  or (_21444_, _21443_, _21440_);
  or (_21445_, _21444_, _42912_);
  or (_21446_, _42908_, \oc8051_golden_model_1.TH0 [4]);
  and (_21447_, _21446_, _41654_);
  and (_43211_, _21447_, _21445_);
  not (_21448_, \oc8051_golden_model_1.TH0 [5]);
  nor (_21451_, _05426_, _21448_);
  and (_21452_, _06941_, _05426_);
  or (_21453_, _21452_, _21451_);
  and (_21454_, _21453_, _04678_);
  and (_21455_, _05426_, \oc8051_golden_model_1.ACC [5]);
  nor (_21456_, _21455_, _21451_);
  nor (_21457_, _21456_, _04616_);
  nor (_21458_, _04615_, _21448_);
  or (_21459_, _21458_, _21457_);
  and (_21460_, _21459_, _04630_);
  nor (_21461_, _13025_, _09375_);
  nor (_21462_, _21461_, _21451_);
  nor (_21463_, _21462_, _04630_);
  or (_21464_, _21463_, _21460_);
  and (_21465_, _21464_, _04537_);
  nor (_21466_, _05799_, _09375_);
  nor (_21467_, _21466_, _21451_);
  nor (_21468_, _21467_, _04537_);
  nor (_21469_, _21468_, _21465_);
  nor (_21470_, _21469_, _03750_);
  nor (_21472_, _21456_, _03751_);
  nor (_21473_, _21472_, _07544_);
  not (_21474_, _21473_);
  nor (_21475_, _21474_, _21470_);
  and (_21476_, _21467_, _07544_);
  or (_21477_, _21476_, _04678_);
  nor (_21478_, _21477_, _21475_);
  or (_21479_, _21478_, _21454_);
  and (_21480_, _21479_, _03415_);
  nor (_21481_, _13118_, _09375_);
  nor (_21483_, _21481_, _21451_);
  nor (_21484_, _21483_, _03415_);
  or (_21485_, _21484_, _08854_);
  or (_21486_, _21485_, _21480_);
  and (_21487_, _13133_, _05426_);
  or (_21488_, _21451_, _04703_);
  nor (_21489_, _21488_, _21487_);
  and (_21490_, _06371_, _05426_);
  nor (_21491_, _21490_, _21451_);
  and (_21492_, _21491_, _03839_);
  or (_21494_, _21492_, _03959_);
  nor (_21495_, _21494_, _21489_);
  and (_21496_, _21495_, _21486_);
  and (_21497_, _10451_, _05426_);
  nor (_21498_, _21497_, _21451_);
  nor (_21499_, _21498_, _04701_);
  nor (_21500_, _21499_, _21496_);
  nor (_21501_, _21500_, _03866_);
  nor (_21502_, _21451_, _08302_);
  not (_21503_, _21502_);
  nor (_21505_, _21491_, _04708_);
  and (_21506_, _21505_, _21503_);
  nor (_21507_, _21506_, _21501_);
  nor (_21508_, _21507_, _03967_);
  nor (_21509_, _21456_, _04706_);
  and (_21510_, _21509_, _21503_);
  or (_21511_, _21510_, _21508_);
  and (_21512_, _21511_, _06532_);
  nor (_21513_, _13131_, _09375_);
  nor (_21514_, _21513_, _21451_);
  nor (_21516_, _21514_, _06532_);
  or (_21517_, _21516_, _21512_);
  and (_21518_, _21517_, _06537_);
  nor (_21519_, _08697_, _09375_);
  nor (_21520_, _21519_, _21451_);
  nor (_21521_, _21520_, _06537_);
  nor (_21522_, _21521_, _21518_);
  nor (_21523_, _21522_, _03703_);
  nor (_21524_, _21462_, _03704_);
  or (_21525_, _21524_, _03701_);
  nor (_21527_, _21525_, _21523_);
  and (_21528_, _13193_, _05426_);
  nor (_21529_, _21528_, _21451_);
  and (_21530_, _21529_, _03701_);
  nor (_21531_, _21530_, _21527_);
  or (_21532_, _21531_, _42912_);
  or (_21533_, _42908_, \oc8051_golden_model_1.TH0 [5]);
  and (_21534_, _21533_, _41654_);
  and (_43212_, _21534_, _21532_);
  not (_21535_, \oc8051_golden_model_1.TH0 [6]);
  nor (_21537_, _05426_, _21535_);
  and (_21538_, _13333_, _05426_);
  nor (_21539_, _21538_, _21537_);
  and (_21540_, _21539_, _03839_);
  nor (_21541_, _06013_, _09375_);
  nor (_21542_, _21541_, _21537_);
  and (_21543_, _21542_, _07544_);
  and (_21544_, _05426_, \oc8051_golden_model_1.ACC [6]);
  nor (_21545_, _21544_, _21537_);
  nor (_21546_, _21545_, _03751_);
  nor (_21548_, _21545_, _04616_);
  nor (_21549_, _04615_, _21535_);
  or (_21550_, _21549_, _21548_);
  and (_21551_, _21550_, _04630_);
  nor (_21552_, _13234_, _09375_);
  nor (_21553_, _21552_, _21537_);
  nor (_21554_, _21553_, _04630_);
  or (_21555_, _21554_, _21551_);
  and (_21556_, _21555_, _04537_);
  nor (_21557_, _21542_, _04537_);
  nor (_21559_, _21557_, _21556_);
  nor (_21560_, _21559_, _03750_);
  or (_21561_, _21560_, _07544_);
  nor (_21562_, _21561_, _21546_);
  nor (_21563_, _21562_, _21543_);
  nor (_21564_, _21563_, _04678_);
  and (_21565_, _06933_, _05426_);
  nor (_21566_, _21537_, _04679_);
  not (_21567_, _21566_);
  nor (_21568_, _21567_, _21565_);
  or (_21569_, _21568_, _07559_);
  nor (_21570_, _21569_, _21564_);
  nor (_21571_, _13326_, _09375_);
  nor (_21572_, _21571_, _21537_);
  nor (_21573_, _21572_, _03415_);
  or (_21574_, _21573_, _03839_);
  nor (_21575_, _21574_, _21570_);
  nor (_21576_, _21575_, _21540_);
  or (_21577_, _21576_, _03838_);
  and (_21578_, _13341_, _05426_);
  or (_21579_, _21537_, _04703_);
  nor (_21580_, _21579_, _21578_);
  nor (_21581_, _21580_, _03959_);
  and (_21582_, _21581_, _21577_);
  and (_21583_, _08695_, _05426_);
  nor (_21584_, _21583_, _21537_);
  nor (_21585_, _21584_, _04701_);
  nor (_21586_, _21585_, _21582_);
  nor (_21587_, _21586_, _03866_);
  nor (_21588_, _21537_, _08289_);
  not (_21590_, _21588_);
  nor (_21591_, _21539_, _04708_);
  and (_21592_, _21591_, _21590_);
  nor (_21593_, _21592_, _21587_);
  nor (_21594_, _21593_, _03967_);
  nor (_21595_, _21545_, _04706_);
  and (_21596_, _21595_, _21590_);
  or (_21597_, _21596_, _21594_);
  and (_21598_, _21597_, _06532_);
  nor (_21599_, _13340_, _09375_);
  nor (_21601_, _21599_, _21537_);
  nor (_21602_, _21601_, _06532_);
  or (_21603_, _21602_, _21598_);
  and (_21604_, _21603_, _06537_);
  nor (_21605_, _08694_, _09375_);
  nor (_21606_, _21605_, _21537_);
  nor (_21607_, _21606_, _06537_);
  or (_21608_, _21607_, _03703_);
  nor (_21609_, _21608_, _21604_);
  and (_21610_, _21553_, _03703_);
  or (_21612_, _21610_, _03701_);
  nor (_21613_, _21612_, _21609_);
  nor (_21614_, _13399_, _09375_);
  nor (_21615_, _21614_, _21537_);
  nor (_21616_, _21615_, _03702_);
  or (_21617_, _21616_, _21613_);
  or (_21618_, _21617_, _42912_);
  or (_21619_, _42908_, \oc8051_golden_model_1.TH0 [6]);
  and (_21620_, _21619_, _41654_);
  and (_43213_, _21620_, _21618_);
  not (_21622_, \oc8051_golden_model_1.TH1 [0]);
  nor (_21623_, _05404_, _21622_);
  nor (_21624_, _05652_, _09454_);
  nor (_21625_, _21624_, _21623_);
  and (_21626_, _21625_, _17066_);
  and (_21627_, _05404_, _04608_);
  nor (_21628_, _21627_, _21623_);
  and (_21629_, _21628_, _07544_);
  and (_21630_, _05404_, \oc8051_golden_model_1.ACC [0]);
  nor (_21631_, _21630_, _21623_);
  nor (_21633_, _21631_, _04616_);
  nor (_21634_, _04615_, _21622_);
  or (_21635_, _21634_, _21633_);
  and (_21636_, _21635_, _04630_);
  nor (_21637_, _21625_, _04630_);
  or (_21638_, _21637_, _21636_);
  and (_21639_, _21638_, _04537_);
  nor (_21640_, _21628_, _04537_);
  nor (_21641_, _21640_, _21639_);
  nor (_21642_, _21641_, _03750_);
  nor (_21644_, _21631_, _03751_);
  nor (_21645_, _21644_, _07544_);
  not (_21646_, _21645_);
  nor (_21647_, _21646_, _21642_);
  nor (_21648_, _21647_, _21629_);
  nor (_21649_, _21648_, _04678_);
  and (_21650_, _06935_, _05404_);
  nor (_21651_, _21623_, _04679_);
  not (_21652_, _21651_);
  nor (_21653_, _21652_, _21650_);
  nor (_21655_, _21653_, _21649_);
  and (_21656_, _21655_, _03415_);
  nor (_21657_, _12119_, _09454_);
  nor (_21658_, _21657_, _21623_);
  nor (_21659_, _21658_, _03415_);
  or (_21660_, _21659_, _21656_);
  and (_21661_, _21660_, _04694_);
  and (_21662_, _05404_, _06428_);
  nor (_21663_, _21662_, _21623_);
  nor (_21664_, _21663_, _04694_);
  or (_21666_, _21664_, _03838_);
  nor (_21667_, _21666_, _21661_);
  and (_21668_, _12133_, _05404_);
  or (_21669_, _21623_, _04703_);
  nor (_21670_, _21669_, _21668_);
  or (_21671_, _21670_, _03959_);
  nor (_21672_, _21671_, _21667_);
  nor (_21673_, _10458_, _09454_);
  nor (_21674_, _21673_, _21623_);
  not (_21675_, _21674_);
  and (_21677_, _08712_, _05404_);
  nor (_21678_, _21677_, _04701_);
  and (_21679_, _21678_, _21675_);
  nor (_21680_, _21679_, _21672_);
  nor (_21681_, _21680_, _03866_);
  and (_21682_, _12013_, _05404_);
  or (_21683_, _21682_, _21623_);
  and (_21684_, _21683_, _03866_);
  or (_21685_, _21684_, _21681_);
  and (_21686_, _21685_, _04706_);
  nor (_21688_, _21677_, _21623_);
  nor (_21689_, _21688_, _04706_);
  or (_21690_, _21689_, _21686_);
  and (_21691_, _21690_, _06532_);
  nor (_21692_, _12132_, _09454_);
  nor (_21693_, _21692_, _21623_);
  nor (_21694_, _21693_, _06532_);
  or (_21695_, _21694_, _21691_);
  and (_21696_, _21695_, _06537_);
  nor (_21697_, _21674_, _06537_);
  nor (_21699_, _21697_, _17066_);
  not (_21700_, _21699_);
  nor (_21701_, _21700_, _21696_);
  nor (_21702_, _21701_, _21626_);
  or (_21703_, _21702_, _42912_);
  or (_21704_, _42908_, \oc8051_golden_model_1.TH1 [0]);
  and (_21705_, _21704_, _41654_);
  and (_43215_, _21705_, _21703_);
  and (_21706_, _06934_, _05404_);
  not (_21707_, \oc8051_golden_model_1.TH1 [1]);
  nor (_21709_, _05404_, _21707_);
  nor (_21710_, _21709_, _04679_);
  not (_21711_, _21710_);
  nor (_21712_, _21711_, _21706_);
  not (_21713_, _21712_);
  and (_21714_, _05404_, \oc8051_golden_model_1.ACC [1]);
  nor (_21715_, _21714_, _21709_);
  nor (_21716_, _21715_, _03751_);
  nor (_21717_, _21715_, _04616_);
  nor (_21718_, _04615_, _21707_);
  or (_21720_, _21718_, _21717_);
  and (_21721_, _21720_, _04630_);
  nor (_21722_, _05404_, \oc8051_golden_model_1.TH1 [1]);
  and (_21723_, _12225_, _05404_);
  nor (_21724_, _21723_, _21722_);
  and (_21725_, _21724_, _03757_);
  or (_21726_, _21725_, _21721_);
  and (_21727_, _21726_, _04537_);
  and (_21728_, _05404_, _04813_);
  nor (_21729_, _21728_, _21709_);
  nor (_21731_, _21729_, _04537_);
  nor (_21732_, _21731_, _21727_);
  nor (_21733_, _21732_, _03750_);
  or (_21734_, _21733_, _07544_);
  nor (_21735_, _21734_, _21716_);
  and (_21736_, _21729_, _07544_);
  nor (_21737_, _21736_, _21735_);
  nor (_21738_, _21737_, _04678_);
  nor (_21739_, _21738_, _07559_);
  and (_21740_, _21739_, _21713_);
  and (_21742_, _12313_, _05404_);
  or (_21743_, _21742_, _03415_);
  nor (_21744_, _21743_, _21722_);
  nor (_21745_, _21744_, _21740_);
  nor (_21746_, _21745_, _08854_);
  nor (_21747_, _12207_, _09454_);
  or (_21748_, _21747_, _04703_);
  and (_21749_, _05404_, _04515_);
  or (_21750_, _21749_, _04694_);
  and (_21751_, _21750_, _21748_);
  nor (_21753_, _21751_, _21722_);
  or (_21754_, _21753_, _03959_);
  nor (_21755_, _21754_, _21746_);
  nor (_21756_, _08710_, _09454_);
  nor (_21757_, _21756_, _21709_);
  and (_21758_, _08709_, _05404_);
  nor (_21759_, _21758_, _21757_);
  nor (_21760_, _21759_, _04701_);
  nor (_21761_, _21760_, _03866_);
  not (_21762_, _21761_);
  nor (_21764_, _21762_, _21755_);
  and (_21765_, _12206_, _05404_);
  or (_21766_, _21765_, _21709_);
  and (_21767_, _21766_, _03866_);
  or (_21768_, _21767_, _21764_);
  and (_21769_, _21768_, _04706_);
  nor (_21770_, _21758_, _21709_);
  nor (_21771_, _21770_, _04706_);
  or (_21772_, _21771_, _21769_);
  and (_21773_, _21772_, _06532_);
  and (_21775_, _21749_, _05602_);
  or (_21776_, _21775_, _06532_);
  nor (_21777_, _21776_, _21722_);
  or (_21778_, _21777_, _21773_);
  and (_21779_, _21778_, _06537_);
  nor (_21780_, _21757_, _06537_);
  or (_21781_, _21780_, _21779_);
  and (_21782_, _21781_, _03704_);
  and (_21783_, _21724_, _03703_);
  or (_21784_, _21783_, _21782_);
  and (_21786_, _21784_, _03702_);
  nor (_21787_, _21723_, _21709_);
  nor (_21788_, _21787_, _03702_);
  nor (_21789_, _21788_, _21786_);
  nand (_21790_, _21789_, _42908_);
  or (_21791_, _42908_, \oc8051_golden_model_1.TH1 [1]);
  and (_21792_, _21791_, _41654_);
  and (_43216_, _21792_, _21790_);
  and (_21793_, _09454_, \oc8051_golden_model_1.TH1 [2]);
  and (_21794_, _06938_, _05404_);
  or (_21796_, _21794_, _21793_);
  and (_21797_, _21796_, _04678_);
  nor (_21798_, _12427_, _09454_);
  or (_21799_, _21798_, _21793_);
  or (_21800_, _21799_, _04630_);
  and (_21801_, _05404_, \oc8051_golden_model_1.ACC [2]);
  or (_21802_, _21801_, _21793_);
  and (_21803_, _21802_, _04615_);
  and (_21804_, _04616_, \oc8051_golden_model_1.TH1 [2]);
  or (_21805_, _21804_, _03757_);
  or (_21807_, _21805_, _21803_);
  and (_21808_, _21807_, _04537_);
  and (_21809_, _21808_, _21800_);
  nor (_21810_, _09454_, _05236_);
  or (_21811_, _21810_, _21793_);
  and (_21812_, _21811_, _03755_);
  or (_21813_, _21812_, _21809_);
  and (_21814_, _21813_, _03751_);
  and (_21815_, _21802_, _03750_);
  or (_21816_, _21815_, _07544_);
  or (_21818_, _21816_, _21814_);
  or (_21819_, _21811_, _06994_);
  and (_21820_, _21819_, _04679_);
  and (_21821_, _21820_, _21818_);
  or (_21822_, _21821_, _07559_);
  or (_21823_, _21822_, _21797_);
  nor (_21824_, _12523_, _09454_);
  or (_21825_, _21793_, _03415_);
  or (_21826_, _21825_, _21824_);
  and (_21827_, _21826_, _04694_);
  and (_21829_, _21827_, _21823_);
  and (_21830_, _05404_, _06457_);
  or (_21831_, _21830_, _21793_);
  and (_21832_, _21831_, _03839_);
  or (_21833_, _21832_, _03838_);
  or (_21834_, _21833_, _21829_);
  and (_21835_, _12537_, _05404_);
  or (_21836_, _21835_, _21793_);
  or (_21837_, _21836_, _04703_);
  and (_21838_, _21837_, _04701_);
  and (_21840_, _21838_, _21834_);
  and (_21841_, _08707_, _05404_);
  or (_21842_, _21841_, _21793_);
  and (_21843_, _21842_, _03959_);
  or (_21844_, _21843_, _21840_);
  and (_21845_, _21844_, _04708_);
  or (_21846_, _21793_, _05700_);
  and (_21847_, _21831_, _03866_);
  and (_21848_, _21847_, _21846_);
  or (_21849_, _21848_, _21845_);
  and (_21851_, _21849_, _04706_);
  and (_21852_, _21802_, _03967_);
  and (_21853_, _21852_, _21846_);
  or (_21854_, _21853_, _03835_);
  or (_21855_, _21854_, _21851_);
  nor (_21856_, _12536_, _09454_);
  or (_21857_, _21793_, _06532_);
  or (_21858_, _21857_, _21856_);
  and (_21859_, _21858_, _06537_);
  and (_21860_, _21859_, _21855_);
  nor (_21862_, _08706_, _09454_);
  or (_21863_, _21862_, _21793_);
  and (_21864_, _21863_, _03954_);
  or (_21865_, _21864_, _03703_);
  or (_21866_, _21865_, _21860_);
  or (_21867_, _21799_, _03704_);
  and (_21868_, _21867_, _03702_);
  and (_21869_, _21868_, _21866_);
  and (_21870_, _12596_, _05404_);
  or (_21871_, _21870_, _21793_);
  and (_21873_, _21871_, _03701_);
  or (_21874_, _21873_, _21869_);
  or (_21875_, _21874_, _42912_);
  or (_21876_, _42908_, \oc8051_golden_model_1.TH1 [2]);
  and (_21877_, _21876_, _41654_);
  and (_43217_, _21877_, _21875_);
  and (_21878_, _09454_, \oc8051_golden_model_1.TH1 [3]);
  nor (_21879_, _12610_, _09454_);
  or (_21880_, _21879_, _21878_);
  or (_21881_, _21880_, _04630_);
  and (_21883_, _05404_, \oc8051_golden_model_1.ACC [3]);
  or (_21884_, _21883_, _21878_);
  and (_21885_, _21884_, _04615_);
  and (_21886_, _04616_, \oc8051_golden_model_1.TH1 [3]);
  or (_21887_, _21886_, _03757_);
  or (_21888_, _21887_, _21885_);
  and (_21889_, _21888_, _04537_);
  and (_21890_, _21889_, _21881_);
  nor (_21891_, _09454_, _05050_);
  or (_21892_, _21891_, _21878_);
  and (_21894_, _21892_, _03755_);
  or (_21895_, _21894_, _21890_);
  and (_21896_, _21895_, _03751_);
  and (_21897_, _21884_, _03750_);
  or (_21898_, _21897_, _07544_);
  or (_21899_, _21898_, _21896_);
  or (_21900_, _21892_, _06994_);
  and (_21901_, _21900_, _21899_);
  or (_21902_, _21901_, _04678_);
  and (_21903_, _06937_, _05404_);
  or (_21905_, _21878_, _04679_);
  or (_21906_, _21905_, _21903_);
  and (_21907_, _21906_, _03415_);
  and (_21908_, _21907_, _21902_);
  nor (_21909_, _12724_, _09454_);
  or (_21910_, _21909_, _21878_);
  and (_21911_, _21910_, _07559_);
  or (_21912_, _21911_, _08854_);
  or (_21913_, _21912_, _21908_);
  and (_21914_, _12738_, _05404_);
  or (_21916_, _21878_, _04703_);
  or (_21917_, _21916_, _21914_);
  and (_21918_, _05404_, _06415_);
  or (_21919_, _21918_, _21878_);
  or (_21920_, _21919_, _04694_);
  and (_21921_, _21920_, _04701_);
  and (_21922_, _21921_, _21917_);
  and (_21923_, _21922_, _21913_);
  and (_21924_, _10455_, _05404_);
  or (_21925_, _21924_, _21878_);
  and (_21927_, _21925_, _03959_);
  or (_21928_, _21927_, _21923_);
  and (_21929_, _21928_, _04708_);
  or (_21930_, _21878_, _05554_);
  and (_21931_, _21919_, _03866_);
  and (_21932_, _21931_, _21930_);
  or (_21933_, _21932_, _21929_);
  and (_21934_, _21933_, _04706_);
  and (_21935_, _21884_, _03967_);
  and (_21936_, _21935_, _21930_);
  or (_21938_, _21936_, _03835_);
  or (_21939_, _21938_, _21934_);
  nor (_21940_, _12737_, _09454_);
  or (_21941_, _21878_, _06532_);
  or (_21942_, _21941_, _21940_);
  and (_21943_, _21942_, _06537_);
  and (_21944_, _21943_, _21939_);
  nor (_21945_, _08701_, _09454_);
  or (_21946_, _21945_, _21878_);
  and (_21947_, _21946_, _03954_);
  or (_21948_, _21947_, _03703_);
  or (_21949_, _21948_, _21944_);
  or (_21950_, _21880_, _03704_);
  and (_21951_, _21950_, _03702_);
  and (_21952_, _21951_, _21949_);
  and (_21953_, _12792_, _05404_);
  or (_21954_, _21953_, _21878_);
  and (_21955_, _21954_, _03701_);
  or (_21956_, _21955_, _21952_);
  or (_21957_, _21956_, _42912_);
  or (_21960_, _42908_, \oc8051_golden_model_1.TH1 [3]);
  and (_21961_, _21960_, _41654_);
  and (_43218_, _21961_, _21957_);
  not (_21962_, \oc8051_golden_model_1.TH1 [4]);
  nor (_21963_, _05404_, _21962_);
  and (_21964_, _06422_, _05404_);
  nor (_21965_, _21964_, _21963_);
  and (_21966_, _21965_, _03839_);
  and (_21967_, _05404_, \oc8051_golden_model_1.ACC [4]);
  nor (_21968_, _21967_, _21963_);
  nor (_21970_, _21968_, _03751_);
  nor (_21971_, _21968_, _04616_);
  nor (_21972_, _04615_, _21962_);
  or (_21973_, _21972_, _21971_);
  and (_21974_, _21973_, _04630_);
  nor (_21975_, _12828_, _09454_);
  nor (_21976_, _21975_, _21963_);
  nor (_21977_, _21976_, _04630_);
  or (_21978_, _21977_, _21974_);
  and (_21979_, _21978_, _04537_);
  nor (_21981_, _05898_, _09454_);
  nor (_21982_, _21981_, _21963_);
  nor (_21983_, _21982_, _04537_);
  nor (_21984_, _21983_, _21979_);
  nor (_21985_, _21984_, _03750_);
  or (_21986_, _21985_, _07544_);
  nor (_21987_, _21986_, _21970_);
  and (_21988_, _21982_, _07544_);
  nor (_21989_, _21988_, _21987_);
  nor (_21990_, _21989_, _04678_);
  and (_21992_, _06942_, _05404_);
  nor (_21993_, _21963_, _04679_);
  not (_21994_, _21993_);
  nor (_21995_, _21994_, _21992_);
  or (_21996_, _21995_, _07559_);
  nor (_21997_, _21996_, _21990_);
  nor (_21998_, _12919_, _09454_);
  nor (_21999_, _21998_, _21963_);
  nor (_22000_, _21999_, _03415_);
  or (_22001_, _22000_, _03839_);
  nor (_22003_, _22001_, _21997_);
  nor (_22004_, _22003_, _21966_);
  or (_22005_, _22004_, _03838_);
  and (_22006_, _12933_, _05404_);
  or (_22007_, _21963_, _04703_);
  nor (_22008_, _22007_, _22006_);
  nor (_22009_, _22008_, _03959_);
  and (_22010_, _22009_, _22005_);
  and (_22011_, _08700_, _05404_);
  nor (_22012_, _22011_, _21963_);
  nor (_22014_, _22012_, _04701_);
  nor (_22015_, _22014_, _22010_);
  nor (_22016_, _22015_, _03866_);
  nor (_22017_, _21963_, _08303_);
  not (_22018_, _22017_);
  nor (_22019_, _21965_, _04708_);
  and (_22020_, _22019_, _22018_);
  nor (_22021_, _22020_, _22016_);
  nor (_22022_, _22021_, _03967_);
  nor (_22023_, _21968_, _04706_);
  and (_22025_, _22023_, _22018_);
  nor (_22026_, _22025_, _03835_);
  not (_22027_, _22026_);
  nor (_22028_, _22027_, _22022_);
  nor (_22029_, _12931_, _09454_);
  or (_22030_, _21963_, _06532_);
  nor (_22031_, _22030_, _22029_);
  or (_22032_, _22031_, _03954_);
  nor (_22033_, _22032_, _22028_);
  nor (_22034_, _08699_, _09454_);
  nor (_22036_, _22034_, _21963_);
  nor (_22037_, _22036_, _06537_);
  or (_22038_, _22037_, _03703_);
  nor (_22039_, _22038_, _22033_);
  and (_22040_, _21976_, _03703_);
  or (_22041_, _22040_, _03701_);
  nor (_22042_, _22041_, _22039_);
  and (_22043_, _12991_, _05404_);
  nor (_22044_, _22043_, _21963_);
  nor (_22045_, _22044_, _03702_);
  or (_22047_, _22045_, _22042_);
  or (_22048_, _22047_, _42912_);
  or (_22049_, _42908_, \oc8051_golden_model_1.TH1 [4]);
  and (_22050_, _22049_, _41654_);
  and (_43219_, _22050_, _22048_);
  not (_22051_, \oc8051_golden_model_1.TH1 [5]);
  nor (_22052_, _05404_, _22051_);
  and (_22053_, _06941_, _05404_);
  or (_22054_, _22053_, _22052_);
  and (_22055_, _22054_, _04678_);
  and (_22057_, _05404_, \oc8051_golden_model_1.ACC [5]);
  nor (_22058_, _22057_, _22052_);
  nor (_22059_, _22058_, _04616_);
  nor (_22060_, _04615_, _22051_);
  or (_22061_, _22060_, _22059_);
  and (_22062_, _22061_, _04630_);
  nor (_22063_, _13025_, _09454_);
  nor (_22064_, _22063_, _22052_);
  nor (_22065_, _22064_, _04630_);
  or (_22066_, _22065_, _22062_);
  and (_22068_, _22066_, _04537_);
  nor (_22069_, _05799_, _09454_);
  nor (_22070_, _22069_, _22052_);
  nor (_22071_, _22070_, _04537_);
  nor (_22072_, _22071_, _22068_);
  nor (_22073_, _22072_, _03750_);
  nor (_22074_, _22058_, _03751_);
  nor (_22075_, _22074_, _07544_);
  not (_22076_, _22075_);
  nor (_22077_, _22076_, _22073_);
  and (_22079_, _22070_, _07544_);
  or (_22080_, _22079_, _04678_);
  nor (_22081_, _22080_, _22077_);
  or (_22082_, _22081_, _22055_);
  and (_22083_, _22082_, _03415_);
  nor (_22084_, _13118_, _09454_);
  nor (_22085_, _22084_, _22052_);
  nor (_22086_, _22085_, _03415_);
  or (_22087_, _22086_, _08854_);
  or (_22088_, _22087_, _22083_);
  and (_22090_, _13133_, _05404_);
  or (_22091_, _22052_, _04703_);
  nor (_22092_, _22091_, _22090_);
  and (_22093_, _06371_, _05404_);
  nor (_22094_, _22093_, _22052_);
  and (_22095_, _22094_, _03839_);
  or (_22096_, _22095_, _03959_);
  nor (_22097_, _22096_, _22092_);
  and (_22098_, _22097_, _22088_);
  and (_22099_, _10451_, _05404_);
  nor (_22101_, _22099_, _22052_);
  nor (_22102_, _22101_, _04701_);
  nor (_22103_, _22102_, _22098_);
  nor (_22104_, _22103_, _03866_);
  nor (_22105_, _22052_, _08302_);
  not (_22106_, _22105_);
  nor (_22107_, _22094_, _04708_);
  and (_22108_, _22107_, _22106_);
  nor (_22109_, _22108_, _22104_);
  nor (_22110_, _22109_, _03967_);
  nor (_22112_, _22058_, _04706_);
  and (_22113_, _22112_, _22106_);
  or (_22114_, _22113_, _22110_);
  and (_22115_, _22114_, _06532_);
  nor (_22116_, _13131_, _09454_);
  nor (_22117_, _22116_, _22052_);
  nor (_22118_, _22117_, _06532_);
  or (_22119_, _22118_, _22115_);
  and (_22120_, _22119_, _06537_);
  nor (_22121_, _08697_, _09454_);
  nor (_22123_, _22121_, _22052_);
  nor (_22124_, _22123_, _06537_);
  nor (_22125_, _22124_, _22120_);
  nor (_22126_, _22125_, _03703_);
  nor (_22127_, _22064_, _03704_);
  or (_22128_, _22127_, _03701_);
  nor (_22129_, _22128_, _22126_);
  and (_22130_, _13193_, _05404_);
  nor (_22131_, _22130_, _22052_);
  and (_22132_, _22131_, _03701_);
  nor (_22134_, _22132_, _22129_);
  or (_22135_, _22134_, _42912_);
  or (_22136_, _42908_, \oc8051_golden_model_1.TH1 [5]);
  and (_22137_, _22136_, _41654_);
  and (_43220_, _22137_, _22135_);
  not (_22138_, \oc8051_golden_model_1.TH1 [6]);
  nor (_22139_, _05404_, _22138_);
  and (_22140_, _13333_, _05404_);
  nor (_22141_, _22140_, _22139_);
  and (_22142_, _22141_, _03839_);
  nor (_22144_, _06013_, _09454_);
  nor (_22145_, _22144_, _22139_);
  and (_22146_, _22145_, _07544_);
  and (_22147_, _05404_, \oc8051_golden_model_1.ACC [6]);
  nor (_22148_, _22147_, _22139_);
  nor (_22149_, _22148_, _04616_);
  nor (_22150_, _04615_, _22138_);
  or (_22151_, _22150_, _22149_);
  and (_22152_, _22151_, _04630_);
  nor (_22153_, _13234_, _09454_);
  nor (_22155_, _22153_, _22139_);
  nor (_22156_, _22155_, _04630_);
  or (_22157_, _22156_, _22152_);
  and (_22158_, _22157_, _04537_);
  nor (_22159_, _22145_, _04537_);
  nor (_22160_, _22159_, _22158_);
  nor (_22161_, _22160_, _03750_);
  nor (_22162_, _22148_, _03751_);
  nor (_22163_, _22162_, _07544_);
  not (_22164_, _22163_);
  nor (_22166_, _22164_, _22161_);
  nor (_22167_, _22166_, _22146_);
  nor (_22168_, _22167_, _04678_);
  and (_22169_, _06933_, _05404_);
  nor (_22170_, _22139_, _04679_);
  not (_22171_, _22170_);
  nor (_22172_, _22171_, _22169_);
  or (_22173_, _22172_, _07559_);
  nor (_22174_, _22173_, _22168_);
  nor (_22175_, _13326_, _09454_);
  nor (_22177_, _22175_, _22139_);
  nor (_22178_, _22177_, _03415_);
  or (_22179_, _22178_, _03839_);
  nor (_22180_, _22179_, _22174_);
  nor (_22181_, _22180_, _22142_);
  or (_22182_, _22181_, _03838_);
  and (_22183_, _13341_, _05404_);
  or (_22184_, _22183_, _22139_);
  or (_22185_, _22184_, _04703_);
  and (_22186_, _22185_, _04701_);
  and (_22188_, _22186_, _22182_);
  and (_22189_, _08695_, _05404_);
  nor (_22190_, _22189_, _22139_);
  nor (_22191_, _22190_, _04701_);
  nor (_22192_, _22191_, _22188_);
  nor (_22193_, _22192_, _03866_);
  nor (_22194_, _22139_, _08289_);
  not (_22195_, _22194_);
  nor (_22196_, _22141_, _04708_);
  and (_22197_, _22196_, _22195_);
  nor (_22199_, _22197_, _22193_);
  nor (_22200_, _22199_, _03967_);
  nor (_22201_, _22148_, _04706_);
  and (_22202_, _22201_, _22195_);
  or (_22203_, _22202_, _22200_);
  and (_22204_, _22203_, _06532_);
  nor (_22205_, _13340_, _09454_);
  nor (_22206_, _22205_, _22139_);
  nor (_22207_, _22206_, _06532_);
  or (_22208_, _22207_, _22204_);
  and (_22210_, _22208_, _06537_);
  nor (_22211_, _08694_, _09454_);
  nor (_22212_, _22211_, _22139_);
  nor (_22213_, _22212_, _06537_);
  or (_22214_, _22213_, _03703_);
  nor (_22215_, _22214_, _22210_);
  and (_22216_, _22155_, _03703_);
  or (_22217_, _22216_, _03701_);
  nor (_22218_, _22217_, _22215_);
  nor (_22219_, _13399_, _09454_);
  nor (_22222_, _22219_, _22139_);
  nor (_22223_, _22222_, _03702_);
  or (_22224_, _22223_, _22218_);
  or (_22225_, _22224_, _42912_);
  or (_22226_, _42908_, \oc8051_golden_model_1.TH1 [6]);
  and (_22227_, _22226_, _41654_);
  and (_43221_, _22227_, _22225_);
  not (_22228_, \oc8051_golden_model_1.TMOD [0]);
  nor (_22229_, _05414_, _22228_);
  nor (_22230_, _05652_, _09536_);
  nor (_22232_, _22230_, _22229_);
  and (_22233_, _22232_, _17066_);
  and (_22234_, _05414_, \oc8051_golden_model_1.ACC [0]);
  nor (_22235_, _22234_, _22229_);
  nor (_22236_, _22235_, _03751_);
  nor (_22237_, _22236_, _07544_);
  nor (_22238_, _22232_, _04630_);
  nor (_22239_, _04615_, _22228_);
  nor (_22240_, _22235_, _04616_);
  nor (_22241_, _22240_, _22239_);
  nor (_22243_, _22241_, _03757_);
  or (_22244_, _22243_, _03755_);
  nor (_22245_, _22244_, _22238_);
  or (_22246_, _22245_, _03750_);
  and (_22247_, _22246_, _22237_);
  and (_22248_, _05414_, _04608_);
  or (_22249_, _22229_, _19847_);
  nor (_22250_, _22249_, _22248_);
  nor (_22251_, _22250_, _22247_);
  nor (_22252_, _22251_, _04678_);
  and (_22254_, _06935_, _05414_);
  nor (_22255_, _22229_, _04679_);
  not (_22256_, _22255_);
  nor (_22257_, _22256_, _22254_);
  nor (_22258_, _22257_, _22252_);
  and (_22259_, _22258_, _03415_);
  nor (_22260_, _12119_, _09536_);
  nor (_22261_, _22260_, _22229_);
  nor (_22262_, _22261_, _03415_);
  or (_22263_, _22262_, _22259_);
  and (_22265_, _22263_, _04694_);
  and (_22266_, _05414_, _06428_);
  nor (_22267_, _22266_, _22229_);
  nor (_22268_, _22267_, _04694_);
  or (_22269_, _22268_, _03838_);
  nor (_22270_, _22269_, _22265_);
  and (_22271_, _12133_, _05414_);
  or (_22272_, _22229_, _04703_);
  nor (_22273_, _22272_, _22271_);
  or (_22274_, _22273_, _03959_);
  nor (_22276_, _22274_, _22270_);
  nor (_22277_, _10458_, _09536_);
  nor (_22278_, _22277_, _22229_);
  not (_22279_, _22278_);
  and (_22280_, _08712_, _05414_);
  nor (_22281_, _22280_, _04701_);
  and (_22282_, _22281_, _22279_);
  nor (_22283_, _22282_, _22276_);
  nor (_22284_, _22283_, _03866_);
  and (_22285_, _12013_, _05414_);
  or (_22287_, _22285_, _22229_);
  and (_22288_, _22287_, _03866_);
  or (_22289_, _22288_, _22284_);
  and (_22290_, _22289_, _04706_);
  nor (_22291_, _22280_, _22229_);
  nor (_22292_, _22291_, _04706_);
  or (_22293_, _22292_, _22290_);
  and (_22294_, _22293_, _06532_);
  nor (_22295_, _12132_, _09536_);
  nor (_22296_, _22295_, _22229_);
  nor (_22298_, _22296_, _06532_);
  or (_22299_, _22298_, _22294_);
  and (_22300_, _22299_, _06537_);
  nor (_22301_, _22278_, _06537_);
  nor (_22302_, _22301_, _17066_);
  not (_22303_, _22302_);
  nor (_22304_, _22303_, _22300_);
  nor (_22305_, _22304_, _22233_);
  or (_22306_, _22305_, _42912_);
  or (_22307_, _42908_, \oc8051_golden_model_1.TMOD [0]);
  and (_22309_, _22307_, _41654_);
  and (_43224_, _22309_, _22306_);
  and (_22310_, _06934_, _05414_);
  not (_22311_, \oc8051_golden_model_1.TMOD [1]);
  nor (_22312_, _05414_, _22311_);
  nor (_22313_, _22312_, _04679_);
  not (_22314_, _22313_);
  nor (_22315_, _22314_, _22310_);
  not (_22316_, _22315_);
  and (_22317_, _05414_, \oc8051_golden_model_1.ACC [1]);
  nor (_22319_, _22317_, _22312_);
  nor (_22320_, _22319_, _03751_);
  nor (_22321_, _22319_, _04616_);
  nor (_22322_, _04615_, _22311_);
  or (_22323_, _22322_, _22321_);
  and (_22324_, _22323_, _04630_);
  nor (_22325_, _05414_, \oc8051_golden_model_1.TMOD [1]);
  and (_22326_, _12225_, _05414_);
  nor (_22327_, _22326_, _22325_);
  and (_22328_, _22327_, _03757_);
  or (_22331_, _22328_, _22324_);
  and (_22332_, _22331_, _04537_);
  and (_22333_, _05414_, _04813_);
  nor (_22334_, _22333_, _22312_);
  nor (_22335_, _22334_, _04537_);
  nor (_22336_, _22335_, _22332_);
  nor (_22337_, _22336_, _03750_);
  or (_22338_, _22337_, _07544_);
  nor (_22339_, _22338_, _22320_);
  and (_22340_, _22334_, _07544_);
  nor (_22342_, _22340_, _22339_);
  nor (_22343_, _22342_, _04678_);
  nor (_22344_, _22343_, _07559_);
  and (_22345_, _22344_, _22316_);
  and (_22346_, _12313_, _05414_);
  or (_22347_, _22346_, _03415_);
  nor (_22348_, _22347_, _22325_);
  nor (_22349_, _22348_, _22345_);
  nor (_22350_, _22349_, _08854_);
  nor (_22351_, _12207_, _09536_);
  or (_22353_, _22351_, _04703_);
  and (_22354_, _05414_, _04515_);
  or (_22355_, _22354_, _04694_);
  and (_22356_, _22355_, _22353_);
  nor (_22357_, _22356_, _22325_);
  or (_22358_, _22357_, _03959_);
  nor (_22359_, _22358_, _22350_);
  nor (_22360_, _08710_, _09536_);
  nor (_22361_, _22360_, _22312_);
  and (_22362_, _08709_, _05414_);
  nor (_22364_, _22362_, _22361_);
  nor (_22365_, _22364_, _04701_);
  nor (_22366_, _22365_, _03866_);
  not (_22367_, _22366_);
  nor (_22368_, _22367_, _22359_);
  and (_22369_, _12206_, _05414_);
  or (_22370_, _22369_, _22312_);
  and (_22371_, _22370_, _03866_);
  or (_22372_, _22371_, _22368_);
  and (_22373_, _22372_, _04706_);
  nor (_22375_, _22362_, _22312_);
  nor (_22376_, _22375_, _04706_);
  or (_22377_, _22376_, _22373_);
  and (_22378_, _22377_, _06532_);
  nor (_22379_, _12205_, _09536_);
  or (_22380_, _22379_, _22312_);
  and (_22381_, _22380_, _03835_);
  or (_22382_, _22381_, _22378_);
  and (_22383_, _22382_, _06537_);
  nor (_22384_, _22361_, _06537_);
  or (_22386_, _22384_, _22383_);
  and (_22387_, _22386_, _03704_);
  and (_22388_, _22327_, _03703_);
  or (_22389_, _22388_, _22387_);
  and (_22390_, _22389_, _03702_);
  nor (_22391_, _22326_, _22312_);
  nor (_22392_, _22391_, _03702_);
  nor (_22393_, _22392_, _22390_);
  nand (_22394_, _22393_, _42908_);
  or (_22395_, _42908_, \oc8051_golden_model_1.TMOD [1]);
  and (_22397_, _22395_, _41654_);
  and (_43225_, _22397_, _22394_);
  not (_22398_, \oc8051_golden_model_1.TMOD [2]);
  nor (_22399_, _05414_, _22398_);
  nor (_22400_, _09536_, _05236_);
  nor (_22401_, _22400_, _22399_);
  and (_22402_, _22401_, _07544_);
  and (_22403_, _05414_, \oc8051_golden_model_1.ACC [2]);
  nor (_22404_, _22403_, _22399_);
  nor (_22405_, _22404_, _03751_);
  nor (_22407_, _22404_, _04616_);
  nor (_22408_, _04615_, _22398_);
  or (_22409_, _22408_, _22407_);
  and (_22410_, _22409_, _04630_);
  nor (_22411_, _12427_, _09536_);
  nor (_22412_, _22411_, _22399_);
  nor (_22413_, _22412_, _04630_);
  or (_22414_, _22413_, _22410_);
  and (_22415_, _22414_, _04537_);
  nor (_22416_, _22401_, _04537_);
  nor (_22418_, _22416_, _22415_);
  nor (_22419_, _22418_, _03750_);
  or (_22420_, _22419_, _07544_);
  nor (_22421_, _22420_, _22405_);
  nor (_22422_, _22421_, _22402_);
  nor (_22423_, _22422_, _04678_);
  and (_22424_, _06938_, _05414_);
  nor (_22425_, _22399_, _04679_);
  not (_22426_, _22425_);
  nor (_22427_, _22426_, _22424_);
  nor (_22429_, _22427_, _07559_);
  not (_22430_, _22429_);
  nor (_22431_, _22430_, _22423_);
  nor (_22432_, _12523_, _09536_);
  nor (_22433_, _22432_, _22399_);
  nor (_22434_, _22433_, _03415_);
  or (_22435_, _22434_, _08854_);
  or (_22436_, _22435_, _22431_);
  and (_22437_, _12537_, _05414_);
  or (_22438_, _22399_, _04703_);
  or (_22440_, _22438_, _22437_);
  and (_22441_, _05414_, _06457_);
  nor (_22442_, _22441_, _22399_);
  and (_22443_, _22442_, _03839_);
  nor (_22444_, _22443_, _03959_);
  and (_22445_, _22444_, _22440_);
  and (_22446_, _22445_, _22436_);
  and (_22447_, _08707_, _05414_);
  nor (_22448_, _22447_, _22399_);
  nor (_22449_, _22448_, _04701_);
  nor (_22451_, _22449_, _22446_);
  nor (_22452_, _22451_, _03866_);
  nor (_22453_, _22399_, _05700_);
  not (_22454_, _22453_);
  nor (_22455_, _22442_, _04708_);
  and (_22456_, _22455_, _22454_);
  nor (_22457_, _22456_, _22452_);
  nor (_22458_, _22457_, _03967_);
  nor (_22459_, _22404_, _04706_);
  and (_22460_, _22459_, _22454_);
  or (_22462_, _22460_, _22458_);
  and (_22463_, _22462_, _06532_);
  nor (_22464_, _12536_, _09536_);
  nor (_22465_, _22464_, _22399_);
  nor (_22466_, _22465_, _06532_);
  or (_22467_, _22466_, _22463_);
  and (_22468_, _22467_, _06537_);
  nor (_22469_, _08706_, _09536_);
  nor (_22470_, _22469_, _22399_);
  nor (_22471_, _22470_, _06537_);
  or (_22473_, _22471_, _03703_);
  nor (_22474_, _22473_, _22468_);
  and (_22475_, _22412_, _03703_);
  or (_22476_, _22475_, _03701_);
  nor (_22477_, _22476_, _22474_);
  and (_22478_, _12596_, _05414_);
  nor (_22479_, _22478_, _22399_);
  nor (_22480_, _22479_, _03702_);
  or (_22481_, _22480_, _22477_);
  or (_22482_, _22481_, _42912_);
  or (_22484_, _42908_, \oc8051_golden_model_1.TMOD [2]);
  and (_22485_, _22484_, _41654_);
  and (_43226_, _22485_, _22482_);
  and (_22486_, _09536_, \oc8051_golden_model_1.TMOD [3]);
  nor (_22487_, _12610_, _09536_);
  or (_22488_, _22487_, _22486_);
  or (_22489_, _22488_, _04630_);
  and (_22490_, _05414_, \oc8051_golden_model_1.ACC [3]);
  or (_22491_, _22490_, _22486_);
  and (_22492_, _22491_, _04615_);
  and (_22494_, _04616_, \oc8051_golden_model_1.TMOD [3]);
  or (_22495_, _22494_, _03757_);
  or (_22496_, _22495_, _22492_);
  and (_22497_, _22496_, _04537_);
  and (_22498_, _22497_, _22489_);
  nor (_22499_, _09536_, _05050_);
  or (_22500_, _22499_, _22486_);
  and (_22501_, _22500_, _03755_);
  or (_22502_, _22501_, _22498_);
  and (_22503_, _22502_, _03751_);
  and (_22505_, _22491_, _03750_);
  or (_22506_, _22505_, _07544_);
  or (_22507_, _22506_, _22503_);
  or (_22508_, _22500_, _06994_);
  and (_22509_, _22508_, _22507_);
  or (_22510_, _22509_, _04678_);
  and (_22511_, _06937_, _05414_);
  or (_22512_, _22486_, _04679_);
  or (_22513_, _22512_, _22511_);
  and (_22514_, _22513_, _03415_);
  and (_22516_, _22514_, _22510_);
  nor (_22517_, _12724_, _09536_);
  or (_22518_, _22517_, _22486_);
  and (_22519_, _22518_, _07559_);
  or (_22520_, _22519_, _08854_);
  or (_22521_, _22520_, _22516_);
  and (_22522_, _12738_, _05414_);
  or (_22523_, _22486_, _04703_);
  or (_22524_, _22523_, _22522_);
  and (_22525_, _05414_, _06415_);
  or (_22527_, _22525_, _22486_);
  or (_22528_, _22527_, _04694_);
  and (_22529_, _22528_, _04701_);
  and (_22530_, _22529_, _22524_);
  and (_22531_, _22530_, _22521_);
  and (_22532_, _10455_, _05414_);
  or (_22533_, _22532_, _22486_);
  and (_22534_, _22533_, _03959_);
  or (_22535_, _22534_, _22531_);
  and (_22536_, _22535_, _04708_);
  or (_22538_, _22486_, _05554_);
  and (_22539_, _22527_, _03866_);
  and (_22540_, _22539_, _22538_);
  or (_22541_, _22540_, _22536_);
  and (_22542_, _22541_, _04706_);
  and (_22543_, _22491_, _03967_);
  and (_22544_, _22543_, _22538_);
  or (_22545_, _22544_, _03835_);
  or (_22546_, _22545_, _22542_);
  nor (_22547_, _12737_, _09536_);
  or (_22549_, _22486_, _06532_);
  or (_22550_, _22549_, _22547_);
  and (_22551_, _22550_, _06537_);
  and (_22552_, _22551_, _22546_);
  nor (_22553_, _08701_, _09536_);
  or (_22554_, _22553_, _22486_);
  and (_22555_, _22554_, _03954_);
  or (_22556_, _22555_, _03703_);
  or (_22557_, _22556_, _22552_);
  or (_22558_, _22488_, _03704_);
  and (_22560_, _22558_, _03702_);
  and (_22561_, _22560_, _22557_);
  and (_22562_, _12792_, _05414_);
  or (_22563_, _22562_, _22486_);
  and (_22564_, _22563_, _03701_);
  or (_22565_, _22564_, _22561_);
  or (_22566_, _22565_, _42912_);
  or (_22567_, _42908_, \oc8051_golden_model_1.TMOD [3]);
  and (_22568_, _22567_, _41654_);
  and (_43227_, _22568_, _22566_);
  not (_22570_, \oc8051_golden_model_1.TMOD [4]);
  nor (_22571_, _05414_, _22570_);
  and (_22572_, _06422_, _05414_);
  nor (_22573_, _22572_, _22571_);
  and (_22574_, _22573_, _03839_);
  and (_22575_, _05414_, \oc8051_golden_model_1.ACC [4]);
  nor (_22576_, _22575_, _22571_);
  nor (_22577_, _22576_, _03751_);
  nor (_22578_, _22576_, _04616_);
  nor (_22579_, _04615_, _22570_);
  or (_22581_, _22579_, _22578_);
  and (_22582_, _22581_, _04630_);
  nor (_22583_, _12828_, _09536_);
  nor (_22584_, _22583_, _22571_);
  nor (_22585_, _22584_, _04630_);
  or (_22586_, _22585_, _22582_);
  and (_22587_, _22586_, _04537_);
  nor (_22588_, _05898_, _09536_);
  nor (_22589_, _22588_, _22571_);
  nor (_22590_, _22589_, _04537_);
  nor (_22592_, _22590_, _22587_);
  nor (_22593_, _22592_, _03750_);
  or (_22594_, _22593_, _07544_);
  nor (_22595_, _22594_, _22577_);
  and (_22596_, _22589_, _07544_);
  nor (_22597_, _22596_, _22595_);
  nor (_22598_, _22597_, _04678_);
  and (_22599_, _06942_, _05414_);
  nor (_22600_, _22571_, _04679_);
  not (_22601_, _22600_);
  nor (_22603_, _22601_, _22599_);
  or (_22604_, _22603_, _07559_);
  nor (_22605_, _22604_, _22598_);
  nor (_22606_, _12919_, _09536_);
  nor (_22607_, _22606_, _22571_);
  nor (_22608_, _22607_, _03415_);
  or (_22609_, _22608_, _03839_);
  nor (_22610_, _22609_, _22605_);
  nor (_22611_, _22610_, _22574_);
  or (_22612_, _22611_, _03838_);
  and (_22614_, _12933_, _05414_);
  or (_22615_, _22614_, _22571_);
  or (_22616_, _22615_, _04703_);
  and (_22617_, _22616_, _04701_);
  and (_22618_, _22617_, _22612_);
  and (_22619_, _08700_, _05414_);
  nor (_22620_, _22619_, _22571_);
  nor (_22621_, _22620_, _04701_);
  nor (_22622_, _22621_, _22618_);
  nor (_22623_, _22622_, _03866_);
  nor (_22625_, _22571_, _08303_);
  not (_22626_, _22625_);
  nor (_22627_, _22573_, _04708_);
  and (_22628_, _22627_, _22626_);
  nor (_22629_, _22628_, _22623_);
  nor (_22630_, _22629_, _03967_);
  nor (_22631_, _22576_, _04706_);
  and (_22632_, _22631_, _22626_);
  or (_22633_, _22632_, _22630_);
  and (_22634_, _22633_, _06532_);
  nor (_22636_, _12931_, _09536_);
  nor (_22637_, _22636_, _22571_);
  nor (_22638_, _22637_, _06532_);
  or (_22639_, _22638_, _22634_);
  and (_22640_, _22639_, _06537_);
  nor (_22641_, _08699_, _09536_);
  nor (_22642_, _22641_, _22571_);
  nor (_22643_, _22642_, _06537_);
  or (_22644_, _22643_, _03703_);
  nor (_22645_, _22644_, _22640_);
  and (_22647_, _22584_, _03703_);
  or (_22648_, _22647_, _03701_);
  nor (_22649_, _22648_, _22645_);
  and (_22650_, _12991_, _05414_);
  nor (_22651_, _22650_, _22571_);
  nor (_22652_, _22651_, _03702_);
  or (_22653_, _22652_, _22649_);
  or (_22654_, _22653_, _42912_);
  or (_22655_, _42908_, \oc8051_golden_model_1.TMOD [4]);
  and (_22656_, _22655_, _41654_);
  and (_43228_, _22656_, _22654_);
  not (_22658_, \oc8051_golden_model_1.TMOD [5]);
  nor (_22659_, _05414_, _22658_);
  and (_22660_, _06941_, _05414_);
  or (_22661_, _22660_, _22659_);
  and (_22662_, _22661_, _04678_);
  and (_22663_, _05414_, \oc8051_golden_model_1.ACC [5]);
  nor (_22664_, _22663_, _22659_);
  nor (_22665_, _22664_, _03751_);
  nor (_22666_, _22664_, _04616_);
  nor (_22668_, _04615_, _22658_);
  or (_22669_, _22668_, _22666_);
  and (_22670_, _22669_, _04630_);
  nor (_22671_, _13025_, _09536_);
  nor (_22672_, _22671_, _22659_);
  nor (_22673_, _22672_, _04630_);
  or (_22674_, _22673_, _22670_);
  and (_22675_, _22674_, _04537_);
  nor (_22676_, _05799_, _09536_);
  nor (_22677_, _22676_, _22659_);
  nor (_22679_, _22677_, _04537_);
  nor (_22680_, _22679_, _22675_);
  nor (_22681_, _22680_, _03750_);
  or (_22682_, _22681_, _07544_);
  nor (_22683_, _22682_, _22665_);
  and (_22684_, _22677_, _07544_);
  or (_22685_, _22684_, _04678_);
  nor (_22686_, _22685_, _22683_);
  or (_22687_, _22686_, _22662_);
  and (_22688_, _22687_, _03415_);
  nor (_22690_, _13118_, _09536_);
  nor (_22691_, _22690_, _22659_);
  nor (_22692_, _22691_, _03415_);
  or (_22693_, _22692_, _08854_);
  or (_22694_, _22693_, _22688_);
  and (_22695_, _13133_, _05414_);
  or (_22696_, _22659_, _04703_);
  nor (_22697_, _22696_, _22695_);
  and (_22698_, _06371_, _05414_);
  nor (_22699_, _22698_, _22659_);
  and (_22701_, _22699_, _03839_);
  or (_22702_, _22701_, _03959_);
  nor (_22703_, _22702_, _22697_);
  and (_22704_, _22703_, _22694_);
  and (_22705_, _10451_, _05414_);
  nor (_22706_, _22705_, _22659_);
  nor (_22707_, _22706_, _04701_);
  nor (_22708_, _22707_, _22704_);
  nor (_22709_, _22708_, _03866_);
  nor (_22710_, _22659_, _08302_);
  not (_22712_, _22710_);
  nor (_22713_, _22699_, _04708_);
  and (_22714_, _22713_, _22712_);
  nor (_22715_, _22714_, _22709_);
  nor (_22716_, _22715_, _03967_);
  nor (_22717_, _22664_, _04706_);
  and (_22718_, _22717_, _22712_);
  nor (_22719_, _22718_, _03835_);
  not (_22720_, _22719_);
  nor (_22721_, _22720_, _22716_);
  nor (_22723_, _13131_, _09536_);
  or (_22724_, _22659_, _06532_);
  nor (_22725_, _22724_, _22723_);
  or (_22726_, _22725_, _03954_);
  nor (_22727_, _22726_, _22721_);
  nor (_22728_, _08697_, _09536_);
  nor (_22729_, _22728_, _22659_);
  nor (_22730_, _22729_, _06537_);
  nor (_22731_, _22730_, _22727_);
  nor (_22732_, _22731_, _03703_);
  nor (_22734_, _22672_, _03704_);
  or (_22735_, _22734_, _03701_);
  nor (_22736_, _22735_, _22732_);
  and (_22737_, _13193_, _05414_);
  nor (_22738_, _22737_, _22659_);
  and (_22739_, _22738_, _03701_);
  nor (_22740_, _22739_, _22736_);
  or (_22741_, _22740_, _42912_);
  or (_22742_, _42908_, \oc8051_golden_model_1.TMOD [5]);
  and (_22743_, _22742_, _41654_);
  and (_43229_, _22743_, _22741_);
  not (_22745_, \oc8051_golden_model_1.TMOD [6]);
  nor (_22746_, _05414_, _22745_);
  and (_22747_, _13333_, _05414_);
  nor (_22748_, _22747_, _22746_);
  and (_22749_, _22748_, _03839_);
  nor (_22750_, _06013_, _09536_);
  nor (_22751_, _22750_, _22746_);
  and (_22752_, _22751_, _07544_);
  and (_22753_, _05414_, \oc8051_golden_model_1.ACC [6]);
  nor (_22755_, _22753_, _22746_);
  nor (_22756_, _22755_, _03751_);
  nor (_22757_, _22755_, _04616_);
  nor (_22758_, _04615_, _22745_);
  or (_22759_, _22758_, _22757_);
  and (_22760_, _22759_, _04630_);
  nor (_22761_, _13234_, _09536_);
  nor (_22762_, _22761_, _22746_);
  nor (_22763_, _22762_, _04630_);
  or (_22764_, _22763_, _22760_);
  and (_22766_, _22764_, _04537_);
  nor (_22767_, _22751_, _04537_);
  nor (_22768_, _22767_, _22766_);
  nor (_22769_, _22768_, _03750_);
  or (_22770_, _22769_, _07544_);
  nor (_22771_, _22770_, _22756_);
  nor (_22772_, _22771_, _22752_);
  nor (_22773_, _22772_, _04678_);
  and (_22774_, _06933_, _05414_);
  nor (_22775_, _22746_, _04679_);
  not (_22777_, _22775_);
  nor (_22778_, _22777_, _22774_);
  or (_22779_, _22778_, _07559_);
  nor (_22780_, _22779_, _22773_);
  nor (_22781_, _13326_, _09536_);
  nor (_22782_, _22781_, _22746_);
  nor (_22783_, _22782_, _03415_);
  or (_22784_, _22783_, _03839_);
  nor (_22785_, _22784_, _22780_);
  nor (_22786_, _22785_, _22749_);
  or (_22788_, _22786_, _03838_);
  and (_22789_, _13341_, _05414_);
  or (_22790_, _22789_, _22746_);
  or (_22791_, _22790_, _04703_);
  and (_22792_, _22791_, _04701_);
  and (_22793_, _22792_, _22788_);
  and (_22794_, _08695_, _05414_);
  nor (_22795_, _22794_, _22746_);
  nor (_22796_, _22795_, _04701_);
  nor (_22797_, _22796_, _22793_);
  nor (_22799_, _22797_, _03866_);
  nor (_22800_, _22746_, _08289_);
  not (_22801_, _22800_);
  nor (_22802_, _22748_, _04708_);
  and (_22803_, _22802_, _22801_);
  nor (_22804_, _22803_, _22799_);
  nor (_22805_, _22804_, _03967_);
  nor (_22806_, _22755_, _04706_);
  and (_22807_, _22806_, _22801_);
  or (_22808_, _22807_, _22805_);
  and (_22810_, _22808_, _06532_);
  nor (_22811_, _13340_, _09536_);
  nor (_22812_, _22811_, _22746_);
  nor (_22813_, _22812_, _06532_);
  or (_22814_, _22813_, _22810_);
  and (_22815_, _22814_, _06537_);
  nor (_22816_, _08694_, _09536_);
  nor (_22817_, _22816_, _22746_);
  nor (_22818_, _22817_, _06537_);
  or (_22819_, _22818_, _03703_);
  nor (_22821_, _22819_, _22815_);
  and (_22822_, _22762_, _03703_);
  or (_22823_, _22822_, _03701_);
  nor (_22824_, _22823_, _22821_);
  nor (_22825_, _13399_, _09536_);
  nor (_22826_, _22825_, _22746_);
  nor (_22827_, _22826_, _03702_);
  or (_22828_, _22827_, _22824_);
  or (_22829_, _22828_, _42912_);
  or (_22830_, _42908_, \oc8051_golden_model_1.TMOD [6]);
  and (_22832_, _22830_, _41654_);
  and (_43230_, _22832_, _22829_);
  not (_22833_, \oc8051_golden_model_1.IE [0]);
  nor (_22834_, _05398_, _22833_);
  nor (_22835_, _05652_, _09594_);
  nor (_22836_, _22835_, _22834_);
  nor (_22837_, _22836_, _03702_);
  and (_22838_, _05398_, _06428_);
  nor (_22839_, _22838_, _22834_);
  and (_22840_, _22839_, _03839_);
  and (_22842_, _05398_, _04608_);
  nor (_22843_, _22842_, _22834_);
  and (_22844_, _22843_, _07544_);
  and (_22845_, _05398_, \oc8051_golden_model_1.ACC [0]);
  nor (_22846_, _22845_, _22834_);
  nor (_22847_, _22846_, _04616_);
  nor (_22848_, _04615_, _22833_);
  or (_22849_, _22848_, _22847_);
  and (_22850_, _22849_, _04630_);
  nor (_22851_, _22836_, _04630_);
  or (_22853_, _22851_, _22850_);
  and (_22854_, _22853_, _03697_);
  nor (_22855_, _06101_, _22833_);
  and (_22856_, _12032_, _06101_);
  nor (_22857_, _22856_, _22855_);
  nor (_22858_, _22857_, _03697_);
  nor (_22859_, _22858_, _22854_);
  nor (_22860_, _22859_, _03755_);
  nor (_22861_, _22843_, _04537_);
  or (_22862_, _22861_, _22860_);
  and (_22864_, _22862_, _03751_);
  nor (_22865_, _22846_, _03751_);
  or (_22866_, _22865_, _22864_);
  and (_22867_, _22866_, _03692_);
  and (_22868_, _22834_, _03691_);
  or (_22869_, _22868_, _22867_);
  and (_22870_, _22869_, _03685_);
  nor (_22871_, _22836_, _03685_);
  or (_22872_, _22871_, _22870_);
  and (_22873_, _22872_, _03680_);
  nor (_22875_, _22855_, _14175_);
  or (_22876_, _22875_, _03680_);
  or (_22877_, _22876_, _22857_);
  and (_22878_, _22877_, _06994_);
  not (_22879_, _22878_);
  nor (_22880_, _22879_, _22873_);
  nor (_22881_, _22880_, _22844_);
  nor (_22882_, _22881_, _04678_);
  and (_22883_, _06935_, _05398_);
  nor (_22884_, _22834_, _04679_);
  not (_22885_, _22884_);
  nor (_22886_, _22885_, _22883_);
  or (_22887_, _22886_, _07559_);
  nor (_22888_, _22887_, _22882_);
  nor (_22889_, _12119_, _09594_);
  nor (_22890_, _22889_, _22834_);
  nor (_22891_, _22890_, _03415_);
  or (_22892_, _22891_, _03839_);
  nor (_22893_, _22892_, _22888_);
  nor (_22894_, _22893_, _22840_);
  or (_22897_, _22894_, _03838_);
  and (_22898_, _12133_, _05398_);
  or (_22899_, _22834_, _04703_);
  nor (_22900_, _22899_, _22898_);
  nor (_22901_, _22900_, _03959_);
  and (_22902_, _22901_, _22897_);
  nor (_22903_, _10458_, _09594_);
  nor (_22904_, _22903_, _22834_);
  and (_22905_, _22845_, _05652_);
  or (_22906_, _22905_, _04701_);
  nor (_22908_, _22906_, _22904_);
  nor (_22909_, _22908_, _22902_);
  nor (_22910_, _22909_, _03866_);
  and (_22911_, _12013_, _05398_);
  or (_22912_, _22911_, _22834_);
  and (_22913_, _22912_, _03866_);
  or (_22914_, _22913_, _22910_);
  and (_22915_, _22914_, _04706_);
  nor (_22916_, _22905_, _22834_);
  nor (_22917_, _22916_, _04706_);
  or (_22918_, _22917_, _22915_);
  and (_22919_, _22918_, _06532_);
  nor (_22920_, _12132_, _09594_);
  nor (_22921_, _22920_, _22834_);
  nor (_22922_, _22921_, _06532_);
  or (_22923_, _22922_, _22919_);
  and (_22924_, _22923_, _06537_);
  nor (_22925_, _22904_, _06537_);
  or (_22926_, _22925_, _03703_);
  or (_22927_, _22926_, _22924_);
  nand (_22930_, _22836_, _03703_);
  and (_22931_, _22930_, _22927_);
  nor (_22932_, _22931_, _03384_);
  nor (_22933_, _22834_, _03385_);
  nor (_22934_, _22933_, _22932_);
  and (_22935_, _22934_, _03702_);
  nor (_22936_, _22935_, _22837_);
  nand (_22937_, _22936_, _42908_);
  or (_22938_, _42908_, \oc8051_golden_model_1.IE [0]);
  and (_22939_, _22938_, _41654_);
  and (_43233_, _22939_, _22937_);
  not (_22941_, \oc8051_golden_model_1.IE [1]);
  nor (_22942_, _05398_, _22941_);
  and (_22943_, _06934_, _05398_);
  or (_22944_, _22943_, _22942_);
  and (_22945_, _22944_, _04678_);
  and (_22946_, _05398_, \oc8051_golden_model_1.ACC [1]);
  nor (_22947_, _22946_, _22942_);
  nor (_22948_, _22947_, _04616_);
  nor (_22949_, _04615_, _22941_);
  or (_22950_, _22949_, _22948_);
  and (_22951_, _22950_, _04630_);
  nor (_22952_, _05398_, \oc8051_golden_model_1.IE [1]);
  and (_22953_, _12225_, _05398_);
  nor (_22954_, _22953_, _22952_);
  and (_22955_, _22954_, _03757_);
  or (_22956_, _22955_, _22951_);
  and (_22957_, _22956_, _03697_);
  nor (_22958_, _06101_, _22941_);
  and (_22959_, _12212_, _06101_);
  nor (_22962_, _22959_, _22958_);
  nor (_22963_, _22962_, _03697_);
  or (_22964_, _22963_, _22957_);
  and (_22965_, _22964_, _04537_);
  and (_22966_, _05398_, _04813_);
  nor (_22967_, _22966_, _22942_);
  nor (_22968_, _22967_, _04537_);
  or (_22969_, _22968_, _22965_);
  and (_22970_, _22969_, _03751_);
  nor (_22971_, _22947_, _03751_);
  or (_22973_, _22971_, _22970_);
  and (_22974_, _22973_, _03692_);
  and (_22975_, _12200_, _06101_);
  nor (_22976_, _22975_, _22958_);
  nor (_22977_, _22976_, _03692_);
  or (_22978_, _22977_, _03684_);
  or (_22979_, _22978_, _22974_);
  and (_22980_, _22959_, _12211_);
  or (_22981_, _22958_, _03685_);
  or (_22982_, _22981_, _22980_);
  and (_22983_, _22982_, _22979_);
  and (_22984_, _22983_, _03680_);
  nor (_22985_, _12256_, _09607_);
  nor (_22986_, _22958_, _22985_);
  nor (_22987_, _22986_, _03680_);
  or (_22988_, _22987_, _07544_);
  nor (_22989_, _22988_, _22984_);
  and (_22990_, _22967_, _07544_);
  or (_22991_, _22990_, _04678_);
  nor (_22992_, _22991_, _22989_);
  or (_22995_, _22992_, _22945_);
  and (_22996_, _22995_, _03415_);
  nor (_22997_, _12313_, _09594_);
  nor (_22998_, _22997_, _22942_);
  nor (_22999_, _22998_, _03415_);
  nor (_23000_, _22999_, _22996_);
  nor (_23001_, _23000_, _08854_);
  nor (_23002_, _12207_, _09594_);
  or (_23003_, _23002_, _04703_);
  and (_23004_, _05398_, _04515_);
  or (_23006_, _23004_, _04694_);
  and (_23007_, _23006_, _23003_);
  nor (_23008_, _23007_, _22952_);
  or (_23009_, _23008_, _03959_);
  nor (_23010_, _23009_, _23001_);
  nor (_23011_, _08710_, _09594_);
  nor (_23012_, _23011_, _22942_);
  and (_23013_, _08709_, _05398_);
  nor (_23014_, _23013_, _23012_);
  nor (_23015_, _23014_, _04701_);
  nor (_23016_, _23015_, _03866_);
  not (_23017_, _23016_);
  nor (_23018_, _23017_, _23010_);
  and (_23019_, _12206_, _05398_);
  or (_23020_, _23019_, _22942_);
  and (_23021_, _23020_, _03866_);
  or (_23022_, _23021_, _23018_);
  and (_23023_, _23022_, _04706_);
  nor (_23024_, _23013_, _22942_);
  nor (_23025_, _23024_, _04706_);
  or (_23028_, _23025_, _23023_);
  and (_23029_, _23028_, _06532_);
  and (_23030_, _23004_, _05602_);
  or (_23031_, _23030_, _06532_);
  nor (_23032_, _23031_, _22952_);
  or (_23033_, _23032_, _23029_);
  and (_23034_, _23033_, _06537_);
  nor (_23035_, _23012_, _06537_);
  or (_23036_, _23035_, _23034_);
  and (_23037_, _23036_, _03704_);
  and (_23039_, _22954_, _03703_);
  or (_23040_, _23039_, _23037_);
  and (_23041_, _23040_, _03385_);
  nor (_23042_, _22976_, _03385_);
  nor (_23043_, _23042_, _03701_);
  not (_23044_, _23043_);
  nor (_23045_, _23044_, _23041_);
  nor (_23046_, _22953_, _22942_);
  and (_23047_, _23046_, _03701_);
  nor (_23048_, _23047_, _23045_);
  or (_23049_, _23048_, _42912_);
  or (_23050_, _42908_, \oc8051_golden_model_1.IE [1]);
  and (_23051_, _23050_, _41654_);
  and (_43234_, _23051_, _23049_);
  not (_23052_, \oc8051_golden_model_1.IE [2]);
  nor (_23053_, _05398_, _23052_);
  and (_23054_, _05398_, _06457_);
  nor (_23055_, _23054_, _23053_);
  and (_23056_, _23055_, _03839_);
  nor (_23057_, _09594_, _05236_);
  nor (_23060_, _23057_, _23053_);
  and (_23061_, _23060_, _07544_);
  and (_23062_, _05398_, \oc8051_golden_model_1.ACC [2]);
  nor (_23063_, _23062_, _23053_);
  nor (_23064_, _23063_, _04616_);
  nor (_23065_, _04615_, _23052_);
  or (_23066_, _23065_, _23064_);
  and (_23067_, _23066_, _04630_);
  nor (_23068_, _12427_, _09594_);
  nor (_23069_, _23068_, _23053_);
  nor (_23071_, _23069_, _04630_);
  or (_23072_, _23071_, _23067_);
  and (_23073_, _23072_, _03697_);
  nor (_23074_, _06101_, _23052_);
  and (_23075_, _12419_, _06101_);
  nor (_23076_, _23075_, _23074_);
  nor (_23077_, _23076_, _03697_);
  or (_23078_, _23077_, _23073_);
  and (_23079_, _23078_, _04537_);
  nor (_23080_, _23060_, _04537_);
  or (_23081_, _23080_, _23079_);
  and (_23082_, _23081_, _03751_);
  nor (_23083_, _23063_, _03751_);
  or (_23084_, _23083_, _23082_);
  and (_23085_, _23084_, _03692_);
  and (_23086_, _12422_, _06101_);
  nor (_23087_, _23086_, _23074_);
  nor (_23088_, _23087_, _03692_);
  or (_23089_, _23088_, _03684_);
  or (_23090_, _23089_, _23085_);
  and (_23093_, _23075_, _12418_);
  or (_23094_, _23074_, _03685_);
  or (_23095_, _23094_, _23093_);
  and (_23096_, _23095_, _03680_);
  and (_23097_, _23096_, _23090_);
  nor (_23098_, _12465_, _09607_);
  nor (_23099_, _23098_, _23074_);
  nor (_23100_, _23099_, _03680_);
  nor (_23101_, _23100_, _07544_);
  not (_23102_, _23101_);
  nor (_23104_, _23102_, _23097_);
  nor (_23105_, _23104_, _23061_);
  nor (_23106_, _23105_, _04678_);
  and (_23107_, _06938_, _05398_);
  nor (_23108_, _23053_, _04679_);
  not (_23109_, _23108_);
  nor (_23110_, _23109_, _23107_);
  or (_23111_, _23110_, _07559_);
  nor (_23112_, _23111_, _23106_);
  nor (_23113_, _12523_, _09594_);
  nor (_23115_, _23053_, _23113_);
  nor (_23116_, _23115_, _03415_);
  or (_23117_, _23116_, _03839_);
  nor (_23118_, _23117_, _23112_);
  nor (_23119_, _23118_, _23056_);
  or (_23120_, _23119_, _03838_);
  and (_23121_, _12537_, _05398_);
  or (_23122_, _23053_, _04703_);
  nor (_23123_, _23122_, _23121_);
  nor (_23124_, _23123_, _03959_);
  and (_23126_, _23124_, _23120_);
  and (_23127_, _08707_, _05398_);
  nor (_23128_, _23127_, _23053_);
  nor (_23129_, _23128_, _04701_);
  nor (_23130_, _23129_, _23126_);
  nor (_23131_, _23130_, _03866_);
  nor (_23132_, _23053_, _05700_);
  not (_23133_, _23132_);
  nor (_23134_, _23055_, _04708_);
  and (_23135_, _23134_, _23133_);
  nor (_23137_, _23135_, _23131_);
  nor (_23138_, _23137_, _03967_);
  nor (_23139_, _23063_, _04706_);
  and (_23140_, _23139_, _23133_);
  or (_23141_, _23140_, _23138_);
  and (_23142_, _23141_, _06532_);
  nor (_23143_, _12536_, _09594_);
  nor (_23144_, _23143_, _23053_);
  nor (_23145_, _23144_, _06532_);
  or (_23146_, _23145_, _23142_);
  and (_23148_, _23146_, _06537_);
  nor (_23149_, _08706_, _09594_);
  nor (_23150_, _23149_, _23053_);
  nor (_23151_, _23150_, _06537_);
  or (_23152_, _23151_, _23148_);
  and (_23153_, _23152_, _03704_);
  nor (_23154_, _23069_, _03704_);
  or (_23155_, _23154_, _23153_);
  and (_23156_, _23155_, _03385_);
  nor (_23157_, _23087_, _03385_);
  or (_23159_, _23157_, _23156_);
  and (_23160_, _23159_, _03702_);
  and (_23161_, _12596_, _05398_);
  nor (_23162_, _23161_, _23053_);
  nor (_23163_, _23162_, _03702_);
  or (_23164_, _23163_, _23160_);
  or (_23165_, _23164_, _42912_);
  or (_23166_, _42908_, \oc8051_golden_model_1.IE [2]);
  and (_23167_, _23166_, _41654_);
  and (_43235_, _23167_, _23165_);
  and (_23169_, _09594_, \oc8051_golden_model_1.IE [3]);
  nor (_23170_, _09594_, _05050_);
  or (_23171_, _23170_, _23169_);
  or (_23172_, _23171_, _06994_);
  nor (_23173_, _12610_, _09594_);
  or (_23174_, _23173_, _23169_);
  or (_23175_, _23174_, _04630_);
  and (_23176_, _05398_, \oc8051_golden_model_1.ACC [3]);
  or (_23177_, _23176_, _23169_);
  and (_23178_, _23177_, _04615_);
  and (_23180_, _04616_, \oc8051_golden_model_1.IE [3]);
  or (_23181_, _23180_, _03757_);
  or (_23182_, _23181_, _23178_);
  and (_23183_, _23182_, _03697_);
  and (_23184_, _23183_, _23175_);
  and (_23185_, _09607_, \oc8051_golden_model_1.IE [3]);
  and (_23186_, _12619_, _06101_);
  or (_23187_, _23186_, _23185_);
  and (_23188_, _23187_, _03696_);
  or (_23189_, _23188_, _03755_);
  or (_23191_, _23189_, _23184_);
  or (_23192_, _23171_, _04537_);
  and (_23193_, _23192_, _23191_);
  or (_23194_, _23193_, _03750_);
  or (_23195_, _23177_, _03751_);
  and (_23196_, _23195_, _03692_);
  and (_23197_, _23196_, _23194_);
  and (_23198_, _12622_, _06101_);
  or (_23199_, _23198_, _23185_);
  and (_23200_, _23199_, _03691_);
  or (_23202_, _23200_, _03684_);
  or (_23203_, _23202_, _23197_);
  or (_23204_, _23185_, _12618_);
  and (_23205_, _23204_, _23187_);
  or (_23206_, _23205_, _03685_);
  and (_23207_, _23206_, _03680_);
  and (_23208_, _23207_, _23203_);
  nor (_23209_, _12665_, _09607_);
  or (_23210_, _23209_, _23185_);
  and (_23211_, _23210_, _03679_);
  or (_23213_, _23211_, _07544_);
  or (_23214_, _23213_, _23208_);
  and (_23215_, _23214_, _23172_);
  or (_23216_, _23215_, _04678_);
  and (_23217_, _06937_, _05398_);
  or (_23218_, _23169_, _04679_);
  or (_23219_, _23218_, _23217_);
  and (_23220_, _23219_, _03415_);
  and (_23221_, _23220_, _23216_);
  nor (_23222_, _12724_, _09594_);
  or (_23224_, _23169_, _23222_);
  and (_23225_, _23224_, _07559_);
  or (_23226_, _23225_, _23221_);
  or (_23227_, _23226_, _08854_);
  and (_23228_, _12738_, _05398_);
  or (_23229_, _23169_, _04703_);
  or (_23230_, _23229_, _23228_);
  and (_23231_, _05398_, _06415_);
  or (_23232_, _23231_, _23169_);
  or (_23233_, _23232_, _04694_);
  and (_23235_, _23233_, _04701_);
  and (_23236_, _23235_, _23230_);
  and (_23237_, _23236_, _23227_);
  and (_23238_, _10455_, _05398_);
  or (_23239_, _23238_, _23169_);
  and (_23240_, _23239_, _03959_);
  or (_23241_, _23240_, _23237_);
  and (_23242_, _23241_, _04708_);
  or (_23243_, _23169_, _05554_);
  and (_23244_, _23232_, _03866_);
  and (_23246_, _23244_, _23243_);
  or (_23247_, _23246_, _23242_);
  and (_23248_, _23247_, _04706_);
  and (_23249_, _23177_, _03967_);
  and (_23250_, _23249_, _23243_);
  or (_23251_, _23250_, _03835_);
  or (_23252_, _23251_, _23248_);
  nor (_23253_, _12737_, _09594_);
  or (_23254_, _23169_, _06532_);
  or (_23255_, _23254_, _23253_);
  and (_23257_, _23255_, _06537_);
  and (_23258_, _23257_, _23252_);
  nor (_23259_, _08701_, _09594_);
  or (_23260_, _23259_, _23169_);
  and (_23261_, _23260_, _03954_);
  or (_23262_, _23261_, _03703_);
  or (_23263_, _23262_, _23258_);
  or (_23264_, _23174_, _03704_);
  and (_23265_, _23264_, _03385_);
  and (_23266_, _23265_, _23263_);
  and (_23268_, _23199_, _03384_);
  or (_23269_, _23268_, _03701_);
  or (_23270_, _23269_, _23266_);
  and (_23271_, _12792_, _05398_);
  or (_23272_, _23271_, _23169_);
  or (_23273_, _23272_, _03702_);
  and (_23274_, _23273_, _23270_);
  or (_23275_, _23274_, _42912_);
  or (_23276_, _42908_, \oc8051_golden_model_1.IE [3]);
  and (_23277_, _23276_, _41654_);
  and (_43236_, _23277_, _23275_);
  and (_23279_, _09594_, \oc8051_golden_model_1.IE [4]);
  nor (_23280_, _05898_, _09594_);
  or (_23281_, _23280_, _23279_);
  or (_23282_, _23281_, _06994_);
  and (_23283_, _09607_, \oc8051_golden_model_1.IE [4]);
  and (_23284_, _12808_, _06101_);
  or (_23285_, _23284_, _23283_);
  and (_23286_, _23285_, _03691_);
  nor (_23287_, _12828_, _09594_);
  or (_23289_, _23287_, _23279_);
  or (_23290_, _23289_, _04630_);
  and (_23291_, _05398_, \oc8051_golden_model_1.ACC [4]);
  or (_23292_, _23291_, _23279_);
  and (_23293_, _23292_, _04615_);
  and (_23294_, _04616_, \oc8051_golden_model_1.IE [4]);
  or (_23295_, _23294_, _03757_);
  or (_23296_, _23295_, _23293_);
  and (_23297_, _23296_, _03697_);
  and (_23298_, _23297_, _23290_);
  and (_23300_, _12832_, _06101_);
  or (_23301_, _23300_, _23283_);
  and (_23302_, _23301_, _03696_);
  or (_23303_, _23302_, _03755_);
  or (_23304_, _23303_, _23298_);
  or (_23305_, _23281_, _04537_);
  and (_23306_, _23305_, _23304_);
  or (_23307_, _23306_, _03750_);
  or (_23308_, _23292_, _03751_);
  and (_23309_, _23308_, _03692_);
  and (_23311_, _23309_, _23307_);
  or (_23312_, _23311_, _23286_);
  and (_23313_, _23312_, _03685_);
  and (_23314_, _12848_, _06101_);
  or (_23315_, _23314_, _23283_);
  and (_23316_, _23315_, _03684_);
  or (_23317_, _23316_, _23313_);
  and (_23318_, _23317_, _03680_);
  nor (_23319_, _12810_, _09607_);
  or (_23320_, _23319_, _23283_);
  and (_23322_, _23320_, _03679_);
  or (_23323_, _23322_, _07544_);
  or (_23324_, _23323_, _23318_);
  and (_23325_, _23324_, _23282_);
  or (_23326_, _23325_, _04678_);
  and (_23327_, _06942_, _05398_);
  or (_23328_, _23279_, _04679_);
  or (_23329_, _23328_, _23327_);
  and (_23330_, _23329_, _03415_);
  and (_23331_, _23330_, _23326_);
  nor (_23333_, _12919_, _09594_);
  or (_23334_, _23333_, _23279_);
  and (_23335_, _23334_, _07559_);
  or (_23336_, _23335_, _08854_);
  or (_23337_, _23336_, _23331_);
  and (_23338_, _12933_, _05398_);
  or (_23339_, _23279_, _04703_);
  or (_23340_, _23339_, _23338_);
  and (_23341_, _06422_, _05398_);
  or (_23342_, _23341_, _23279_);
  or (_23344_, _23342_, _04694_);
  and (_23345_, _23344_, _04701_);
  and (_23346_, _23345_, _23340_);
  and (_23347_, _23346_, _23337_);
  and (_23348_, _08700_, _05398_);
  or (_23349_, _23348_, _23279_);
  and (_23350_, _23349_, _03959_);
  or (_23351_, _23350_, _23347_);
  and (_23352_, _23351_, _04708_);
  or (_23353_, _23279_, _08303_);
  and (_23355_, _23342_, _03866_);
  and (_23356_, _23355_, _23353_);
  or (_23357_, _23356_, _23352_);
  and (_23358_, _23357_, _04706_);
  and (_23359_, _23292_, _03967_);
  and (_23360_, _23359_, _23353_);
  or (_23361_, _23360_, _03835_);
  or (_23362_, _23361_, _23358_);
  nor (_23363_, _12931_, _09594_);
  or (_23364_, _23279_, _06532_);
  or (_23366_, _23364_, _23363_);
  and (_23367_, _23366_, _06537_);
  and (_23368_, _23367_, _23362_);
  nor (_23369_, _08699_, _09594_);
  or (_23370_, _23369_, _23279_);
  and (_23371_, _23370_, _03954_);
  or (_23372_, _23371_, _03703_);
  or (_23373_, _23372_, _23368_);
  or (_23374_, _23289_, _03704_);
  and (_23375_, _23374_, _03385_);
  and (_23377_, _23375_, _23373_);
  and (_23378_, _23285_, _03384_);
  or (_23379_, _23378_, _03701_);
  or (_23380_, _23379_, _23377_);
  and (_23381_, _12991_, _05398_);
  or (_23382_, _23381_, _23279_);
  or (_23383_, _23382_, _03702_);
  and (_23384_, _23383_, _23380_);
  or (_23385_, _23384_, _42912_);
  or (_23386_, _42908_, \oc8051_golden_model_1.IE [4]);
  and (_23388_, _23386_, _41654_);
  and (_43237_, _23388_, _23385_);
  and (_23389_, _09594_, \oc8051_golden_model_1.IE [5]);
  nor (_23390_, _13025_, _09594_);
  or (_23391_, _23390_, _23389_);
  or (_23392_, _23391_, _04630_);
  and (_23393_, _05398_, \oc8051_golden_model_1.ACC [5]);
  or (_23394_, _23393_, _23389_);
  and (_23395_, _23394_, _04615_);
  and (_23396_, _04616_, \oc8051_golden_model_1.IE [5]);
  or (_23398_, _23396_, _03757_);
  or (_23399_, _23398_, _23395_);
  and (_23400_, _23399_, _03697_);
  and (_23401_, _23400_, _23392_);
  and (_23402_, _09607_, \oc8051_golden_model_1.IE [5]);
  and (_23403_, _13029_, _06101_);
  or (_23404_, _23403_, _23402_);
  and (_23405_, _23404_, _03696_);
  or (_23406_, _23405_, _03755_);
  or (_23407_, _23406_, _23401_);
  nor (_23409_, _05799_, _09594_);
  or (_23410_, _23409_, _23389_);
  or (_23411_, _23410_, _04537_);
  and (_23412_, _23411_, _23407_);
  or (_23413_, _23412_, _03750_);
  or (_23414_, _23394_, _03751_);
  and (_23415_, _23414_, _03692_);
  and (_23416_, _23415_, _23413_);
  and (_23417_, _13007_, _06101_);
  or (_23418_, _23417_, _23402_);
  and (_23420_, _23418_, _03691_);
  or (_23421_, _23420_, _03684_);
  or (_23422_, _23421_, _23416_);
  or (_23423_, _23402_, _13044_);
  and (_23424_, _23423_, _23404_);
  or (_23425_, _23424_, _03685_);
  and (_23426_, _23425_, _03680_);
  and (_23427_, _23426_, _23422_);
  nor (_23428_, _13009_, _09607_);
  or (_23429_, _23428_, _23402_);
  and (_23431_, _23429_, _03679_);
  or (_23432_, _23431_, _07544_);
  or (_23433_, _23432_, _23427_);
  or (_23434_, _23410_, _06994_);
  and (_23435_, _23434_, _23433_);
  or (_23436_, _23435_, _04678_);
  and (_23437_, _06941_, _05398_);
  or (_23438_, _23389_, _04679_);
  or (_23439_, _23438_, _23437_);
  and (_23440_, _23439_, _03415_);
  and (_23442_, _23440_, _23436_);
  nor (_23443_, _13118_, _09594_);
  or (_23444_, _23443_, _23389_);
  and (_23445_, _23444_, _07559_);
  or (_23446_, _23445_, _08854_);
  or (_23447_, _23446_, _23442_);
  and (_23448_, _13133_, _05398_);
  or (_23449_, _23389_, _04703_);
  or (_23450_, _23449_, _23448_);
  and (_23451_, _06371_, _05398_);
  or (_23453_, _23451_, _23389_);
  or (_23454_, _23453_, _04694_);
  and (_23455_, _23454_, _04701_);
  and (_23456_, _23455_, _23450_);
  and (_23457_, _23456_, _23447_);
  and (_23458_, _10451_, _05398_);
  or (_23459_, _23458_, _23389_);
  and (_23460_, _23459_, _03959_);
  or (_23461_, _23460_, _23457_);
  and (_23462_, _23461_, _04708_);
  or (_23464_, _23389_, _08302_);
  and (_23465_, _23453_, _03866_);
  and (_23466_, _23465_, _23464_);
  or (_23467_, _23466_, _23462_);
  and (_23468_, _23467_, _04706_);
  and (_23469_, _23394_, _03967_);
  and (_23470_, _23469_, _23464_);
  or (_23471_, _23470_, _03835_);
  or (_23472_, _23471_, _23468_);
  nor (_23473_, _13131_, _09594_);
  or (_23475_, _23389_, _06532_);
  or (_23476_, _23475_, _23473_);
  and (_23477_, _23476_, _06537_);
  and (_23478_, _23477_, _23472_);
  nor (_23479_, _08697_, _09594_);
  or (_23480_, _23479_, _23389_);
  and (_23481_, _23480_, _03954_);
  or (_23482_, _23481_, _03703_);
  or (_23483_, _23482_, _23478_);
  or (_23484_, _23391_, _03704_);
  and (_23486_, _23484_, _03385_);
  and (_23487_, _23486_, _23483_);
  and (_23488_, _23418_, _03384_);
  or (_23489_, _23488_, _03701_);
  or (_23490_, _23489_, _23487_);
  and (_23491_, _13193_, _05398_);
  or (_23492_, _23491_, _23389_);
  or (_23493_, _23492_, _03702_);
  and (_23494_, _23493_, _23490_);
  or (_23495_, _23494_, _42912_);
  or (_23497_, _42908_, \oc8051_golden_model_1.IE [5]);
  and (_23498_, _23497_, _41654_);
  and (_43238_, _23498_, _23495_);
  and (_23499_, _09594_, \oc8051_golden_model_1.IE [6]);
  nor (_23500_, _06013_, _09594_);
  or (_23501_, _23500_, _23499_);
  or (_23502_, _23501_, _06994_);
  and (_23503_, _09607_, \oc8051_golden_model_1.IE [6]);
  and (_23504_, _13218_, _06101_);
  or (_23505_, _23504_, _23503_);
  and (_23507_, _23505_, _03691_);
  nor (_23508_, _13234_, _09594_);
  or (_23509_, _23508_, _23499_);
  or (_23510_, _23509_, _04630_);
  and (_23511_, _05398_, \oc8051_golden_model_1.ACC [6]);
  or (_23512_, _23511_, _23499_);
  and (_23513_, _23512_, _04615_);
  and (_23514_, _04616_, \oc8051_golden_model_1.IE [6]);
  or (_23515_, _23514_, _03757_);
  or (_23516_, _23515_, _23513_);
  and (_23518_, _23516_, _03697_);
  and (_23519_, _23518_, _23510_);
  and (_23520_, _13238_, _06101_);
  or (_23521_, _23520_, _23503_);
  and (_23522_, _23521_, _03696_);
  or (_23523_, _23522_, _03755_);
  or (_23524_, _23523_, _23519_);
  or (_23525_, _23501_, _04537_);
  and (_23526_, _23525_, _23524_);
  or (_23527_, _23526_, _03750_);
  or (_23529_, _23512_, _03751_);
  and (_23530_, _23529_, _03692_);
  and (_23531_, _23530_, _23527_);
  or (_23532_, _23531_, _23507_);
  and (_23533_, _23532_, _03685_);
  or (_23534_, _23503_, _13253_);
  and (_23535_, _23534_, _03684_);
  and (_23536_, _23535_, _23521_);
  or (_23537_, _23536_, _23533_);
  and (_23538_, _23537_, _03680_);
  nor (_23540_, _13220_, _09607_);
  or (_23541_, _23540_, _23503_);
  and (_23542_, _23541_, _03679_);
  or (_23543_, _23542_, _07544_);
  or (_23544_, _23543_, _23538_);
  and (_23545_, _23544_, _23502_);
  or (_23546_, _23545_, _04678_);
  and (_23547_, _06933_, _05398_);
  or (_23548_, _23499_, _04679_);
  or (_23549_, _23548_, _23547_);
  and (_23551_, _23549_, _03415_);
  and (_23552_, _23551_, _23546_);
  nor (_23553_, _13326_, _09594_);
  or (_23554_, _23553_, _23499_);
  and (_23555_, _23554_, _07559_);
  or (_23556_, _23555_, _08854_);
  or (_23557_, _23556_, _23552_);
  and (_23558_, _13341_, _05398_);
  or (_23559_, _23499_, _04703_);
  or (_23560_, _23559_, _23558_);
  and (_23562_, _13333_, _05398_);
  or (_23563_, _23562_, _23499_);
  or (_23564_, _23563_, _04694_);
  and (_23565_, _23564_, _04701_);
  and (_23566_, _23565_, _23560_);
  and (_23567_, _23566_, _23557_);
  and (_23568_, _08695_, _05398_);
  or (_23569_, _23568_, _23499_);
  and (_23570_, _23569_, _03959_);
  or (_23571_, _23570_, _23567_);
  and (_23573_, _23571_, _04708_);
  or (_23574_, _23499_, _08289_);
  and (_23575_, _23563_, _03866_);
  and (_23576_, _23575_, _23574_);
  or (_23577_, _23576_, _23573_);
  and (_23578_, _23577_, _04706_);
  and (_23579_, _23512_, _03967_);
  and (_23580_, _23579_, _23574_);
  or (_23581_, _23580_, _03835_);
  or (_23582_, _23581_, _23578_);
  nor (_23584_, _13340_, _09594_);
  or (_23585_, _23499_, _06532_);
  or (_23586_, _23585_, _23584_);
  and (_23587_, _23586_, _06537_);
  and (_23588_, _23587_, _23582_);
  nor (_23589_, _08694_, _09594_);
  or (_23590_, _23589_, _23499_);
  and (_23591_, _23590_, _03954_);
  or (_23592_, _23591_, _03703_);
  or (_23593_, _23592_, _23588_);
  or (_23595_, _23509_, _03704_);
  and (_23596_, _23595_, _03385_);
  and (_23597_, _23596_, _23593_);
  and (_23598_, _23505_, _03384_);
  or (_23599_, _23598_, _03701_);
  or (_23600_, _23599_, _23597_);
  nor (_23601_, _13399_, _09594_);
  or (_23602_, _23601_, _23499_);
  or (_23603_, _23602_, _03702_);
  and (_23604_, _23603_, _23600_);
  or (_23606_, _23604_, _42912_);
  or (_23607_, _42908_, \oc8051_golden_model_1.IE [6]);
  and (_23608_, _23607_, _41654_);
  and (_43239_, _23608_, _23606_);
  not (_23609_, \oc8051_golden_model_1.IP [0]);
  nor (_23610_, _05347_, _23609_);
  nor (_23611_, _05652_, _09696_);
  nor (_23612_, _23611_, _23610_);
  nor (_23613_, _23612_, _03702_);
  and (_23614_, _05347_, _06428_);
  nor (_23616_, _23614_, _23610_);
  and (_23617_, _23616_, _03839_);
  and (_23618_, _05347_, _04608_);
  nor (_23619_, _23618_, _23610_);
  and (_23620_, _23619_, _07544_);
  and (_23621_, _05347_, \oc8051_golden_model_1.ACC [0]);
  nor (_23622_, _23621_, _23610_);
  nor (_23623_, _23622_, _04616_);
  nor (_23624_, _04615_, _23609_);
  or (_23625_, _23624_, _23623_);
  and (_23627_, _23625_, _04630_);
  nor (_23628_, _23612_, _04630_);
  or (_23629_, _23628_, _23627_);
  and (_23630_, _23629_, _03697_);
  nor (_23631_, _06089_, _23609_);
  and (_23632_, _12032_, _06089_);
  nor (_23633_, _23632_, _23631_);
  nor (_23634_, _23633_, _03697_);
  nor (_23635_, _23634_, _23630_);
  nor (_23636_, _23635_, _03755_);
  nor (_23638_, _23619_, _04537_);
  or (_23639_, _23638_, _23636_);
  and (_23640_, _23639_, _03751_);
  nor (_23641_, _23622_, _03751_);
  or (_23642_, _23641_, _23640_);
  and (_23643_, _23642_, _03692_);
  and (_23644_, _23610_, _03691_);
  or (_23645_, _23644_, _23643_);
  and (_23646_, _23645_, _03685_);
  nor (_23647_, _23612_, _03685_);
  or (_23649_, _23647_, _23646_);
  and (_23650_, _23649_, _03680_);
  nor (_23651_, _23631_, _14175_);
  or (_23652_, _23651_, _03680_);
  nor (_23653_, _23652_, _23633_);
  nor (_23654_, _23653_, _07544_);
  not (_23655_, _23654_);
  nor (_23656_, _23655_, _23650_);
  nor (_23657_, _23656_, _23620_);
  nor (_23658_, _23657_, _04678_);
  and (_23660_, _06935_, _05347_);
  nor (_23661_, _23610_, _04679_);
  not (_23662_, _23661_);
  nor (_23663_, _23662_, _23660_);
  or (_23664_, _23663_, _07559_);
  nor (_23665_, _23664_, _23658_);
  nor (_23666_, _12119_, _09696_);
  nor (_23667_, _23666_, _23610_);
  nor (_23668_, _23667_, _03415_);
  or (_23669_, _23668_, _03839_);
  nor (_23671_, _23669_, _23665_);
  nor (_23672_, _23671_, _23617_);
  or (_23673_, _23672_, _03838_);
  and (_23674_, _12133_, _05347_);
  or (_23675_, _23610_, _04703_);
  nor (_23676_, _23675_, _23674_);
  nor (_23677_, _23676_, _03959_);
  and (_23678_, _23677_, _23673_);
  nor (_23679_, _10458_, _09696_);
  nor (_23680_, _23679_, _23610_);
  and (_23682_, _23621_, _05652_);
  or (_23683_, _23682_, _04701_);
  nor (_23684_, _23683_, _23680_);
  nor (_23685_, _23684_, _23678_);
  nor (_23686_, _23685_, _03866_);
  and (_23687_, _12013_, _05347_);
  or (_23688_, _23687_, _23610_);
  and (_23689_, _23688_, _03866_);
  or (_23690_, _23689_, _23686_);
  and (_23691_, _23690_, _04706_);
  nor (_23693_, _23682_, _23610_);
  nor (_23694_, _23693_, _04706_);
  or (_23695_, _23694_, _23691_);
  and (_23696_, _23695_, _06532_);
  nor (_23697_, _12132_, _09696_);
  nor (_23698_, _23697_, _23610_);
  nor (_23699_, _23698_, _06532_);
  or (_23700_, _23699_, _23696_);
  and (_23701_, _23700_, _06537_);
  nor (_23702_, _23680_, _06537_);
  or (_23704_, _23702_, _03703_);
  or (_23705_, _23704_, _23701_);
  nand (_23706_, _23612_, _03703_);
  and (_23707_, _23706_, _23705_);
  nor (_23708_, _23707_, _03384_);
  nor (_23709_, _23610_, _03385_);
  nor (_23710_, _23709_, _23708_);
  and (_23711_, _23710_, _03702_);
  nor (_23712_, _23711_, _23613_);
  nand (_23713_, _23712_, _42908_);
  or (_23715_, _42908_, \oc8051_golden_model_1.IP [0]);
  and (_23716_, _23715_, _41654_);
  and (_43240_, _23716_, _23713_);
  not (_23717_, \oc8051_golden_model_1.IP [1]);
  nor (_23718_, _05347_, _23717_);
  and (_23719_, _06934_, _05347_);
  or (_23720_, _23719_, _23718_);
  and (_23721_, _23720_, _04678_);
  and (_23722_, _05347_, \oc8051_golden_model_1.ACC [1]);
  nor (_23723_, _23722_, _23718_);
  nor (_23725_, _23723_, _04616_);
  nor (_23726_, _04615_, _23717_);
  or (_23727_, _23726_, _23725_);
  and (_23728_, _23727_, _04630_);
  nor (_23729_, _05347_, \oc8051_golden_model_1.IP [1]);
  and (_23730_, _12225_, _05347_);
  nor (_23731_, _23730_, _23729_);
  and (_23732_, _23731_, _03757_);
  or (_23733_, _23732_, _23728_);
  and (_23734_, _23733_, _03697_);
  nor (_23736_, _06089_, _23717_);
  and (_23737_, _12212_, _06089_);
  nor (_23738_, _23737_, _23736_);
  nor (_23739_, _23738_, _03697_);
  or (_23740_, _23739_, _23734_);
  and (_23741_, _23740_, _04537_);
  and (_23742_, _05347_, _04813_);
  nor (_23743_, _23742_, _23718_);
  nor (_23744_, _23743_, _04537_);
  or (_23745_, _23744_, _23741_);
  and (_23747_, _23745_, _03751_);
  nor (_23748_, _23723_, _03751_);
  or (_23749_, _23748_, _23747_);
  and (_23750_, _23749_, _03692_);
  and (_23751_, _12200_, _06089_);
  nor (_23752_, _23751_, _23736_);
  nor (_23753_, _23752_, _03692_);
  or (_23754_, _23753_, _03684_);
  or (_23755_, _23754_, _23750_);
  and (_23756_, _23737_, _12211_);
  or (_23758_, _23736_, _03685_);
  or (_23759_, _23758_, _23756_);
  and (_23760_, _23759_, _23755_);
  and (_23761_, _23760_, _03680_);
  nor (_23762_, _12256_, _09709_);
  nor (_23763_, _23736_, _23762_);
  nor (_23764_, _23763_, _03680_);
  or (_23765_, _23764_, _07544_);
  nor (_23766_, _23765_, _23761_);
  and (_23767_, _23743_, _07544_);
  or (_23769_, _23767_, _04678_);
  nor (_23770_, _23769_, _23766_);
  or (_23771_, _23770_, _23721_);
  and (_23772_, _23771_, _03415_);
  nor (_23773_, _12313_, _09696_);
  nor (_23774_, _23773_, _23718_);
  nor (_23775_, _23774_, _03415_);
  nor (_23776_, _23775_, _23772_);
  nor (_23777_, _23776_, _08854_);
  nor (_23778_, _12207_, _09696_);
  or (_23779_, _23778_, _04703_);
  and (_23780_, _05347_, _04515_);
  or (_23781_, _23780_, _04694_);
  and (_23782_, _23781_, _23779_);
  nor (_23783_, _23782_, _23729_);
  or (_23784_, _23783_, _03959_);
  nor (_23785_, _23784_, _23777_);
  nor (_23786_, _08710_, _09696_);
  nor (_23787_, _23786_, _23718_);
  and (_23788_, _08709_, _05347_);
  nor (_23790_, _23788_, _23787_);
  nor (_23791_, _23790_, _04701_);
  nor (_23792_, _23791_, _03866_);
  not (_23793_, _23792_);
  nor (_23794_, _23793_, _23785_);
  and (_23795_, _12206_, _05347_);
  or (_23796_, _23795_, _23718_);
  and (_23797_, _23796_, _03866_);
  or (_23798_, _23797_, _23794_);
  and (_23799_, _23798_, _04706_);
  nor (_23801_, _23788_, _23718_);
  nor (_23802_, _23801_, _04706_);
  or (_23803_, _23802_, _23799_);
  and (_23804_, _23803_, _06532_);
  nor (_23805_, _12205_, _09696_);
  or (_23806_, _23805_, _23718_);
  and (_23807_, _23806_, _03835_);
  or (_23808_, _23807_, _23804_);
  and (_23809_, _23808_, _06537_);
  nor (_23810_, _23787_, _06537_);
  or (_23811_, _23810_, _23809_);
  and (_23812_, _23811_, _03704_);
  and (_23813_, _23731_, _03703_);
  or (_23814_, _23813_, _23812_);
  and (_23815_, _23814_, _03385_);
  nor (_23816_, _23752_, _03385_);
  nor (_23817_, _23816_, _03701_);
  not (_23818_, _23817_);
  nor (_23819_, _23818_, _23815_);
  nor (_23820_, _23730_, _23718_);
  and (_23821_, _23820_, _03701_);
  nor (_23822_, _23821_, _23819_);
  or (_23823_, _23822_, _42912_);
  or (_23824_, _42908_, \oc8051_golden_model_1.IP [1]);
  and (_23825_, _23824_, _41654_);
  and (_43243_, _23825_, _23823_);
  not (_23826_, \oc8051_golden_model_1.IP [2]);
  nor (_23827_, _05347_, _23826_);
  and (_23828_, _05347_, _06457_);
  nor (_23829_, _23828_, _23827_);
  and (_23830_, _23829_, _03839_);
  nor (_23831_, _09696_, _05236_);
  nor (_23832_, _23831_, _23827_);
  and (_23833_, _23832_, _07544_);
  and (_23834_, _05347_, \oc8051_golden_model_1.ACC [2]);
  nor (_23835_, _23834_, _23827_);
  nor (_23836_, _23835_, _04616_);
  nor (_23837_, _04615_, _23826_);
  or (_23838_, _23837_, _23836_);
  and (_23839_, _23838_, _04630_);
  nor (_23840_, _12427_, _09696_);
  nor (_23841_, _23840_, _23827_);
  nor (_23842_, _23841_, _04630_);
  or (_23843_, _23842_, _23839_);
  and (_23844_, _23843_, _03697_);
  nor (_23845_, _06089_, _23826_);
  and (_23846_, _12419_, _06089_);
  nor (_23847_, _23846_, _23845_);
  nor (_23848_, _23847_, _03697_);
  or (_23849_, _23848_, _23844_);
  and (_23850_, _23849_, _04537_);
  nor (_23851_, _23832_, _04537_);
  or (_23852_, _23851_, _23850_);
  and (_23853_, _23852_, _03751_);
  nor (_23854_, _23835_, _03751_);
  or (_23855_, _23854_, _23853_);
  and (_23856_, _23855_, _03692_);
  and (_23857_, _12422_, _06089_);
  nor (_23858_, _23857_, _23845_);
  nor (_23859_, _23858_, _03692_);
  or (_23861_, _23859_, _03684_);
  or (_23862_, _23861_, _23856_);
  and (_23863_, _23846_, _12418_);
  or (_23864_, _23845_, _03685_);
  or (_23865_, _23864_, _23863_);
  and (_23866_, _23865_, _03680_);
  and (_23867_, _23866_, _23862_);
  nor (_23868_, _12465_, _09709_);
  nor (_23869_, _23868_, _23845_);
  nor (_23870_, _23869_, _03680_);
  nor (_23872_, _23870_, _07544_);
  not (_23873_, _23872_);
  nor (_23874_, _23873_, _23867_);
  nor (_23875_, _23874_, _23833_);
  nor (_23876_, _23875_, _04678_);
  and (_23877_, _06938_, _05347_);
  nor (_23878_, _23827_, _04679_);
  not (_23879_, _23878_);
  nor (_23880_, _23879_, _23877_);
  or (_23881_, _23880_, _07559_);
  nor (_23882_, _23881_, _23876_);
  nor (_23883_, _12523_, _09696_);
  nor (_23884_, _23827_, _23883_);
  nor (_23885_, _23884_, _03415_);
  or (_23886_, _23885_, _03839_);
  nor (_23887_, _23886_, _23882_);
  nor (_23888_, _23887_, _23830_);
  or (_23889_, _23888_, _03838_);
  and (_23890_, _12537_, _05347_);
  or (_23891_, _23827_, _04703_);
  nor (_23893_, _23891_, _23890_);
  nor (_23894_, _23893_, _03959_);
  and (_23895_, _23894_, _23889_);
  and (_23896_, _08707_, _05347_);
  nor (_23897_, _23896_, _23827_);
  nor (_23898_, _23897_, _04701_);
  nor (_23899_, _23898_, _23895_);
  nor (_23900_, _23899_, _03866_);
  nor (_23901_, _23827_, _05700_);
  not (_23902_, _23901_);
  nor (_23904_, _23829_, _04708_);
  and (_23905_, _23904_, _23902_);
  nor (_23906_, _23905_, _23900_);
  nor (_23907_, _23906_, _03967_);
  nor (_23908_, _23835_, _04706_);
  and (_23909_, _23908_, _23902_);
  nor (_23910_, _23909_, _03835_);
  not (_23911_, _23910_);
  nor (_23912_, _23911_, _23907_);
  nor (_23913_, _12536_, _09696_);
  or (_23915_, _23827_, _06532_);
  nor (_23916_, _23915_, _23913_);
  or (_23917_, _23916_, _03954_);
  nor (_23918_, _23917_, _23912_);
  nor (_23919_, _08706_, _09696_);
  nor (_23920_, _23919_, _23827_);
  nor (_23921_, _23920_, _06537_);
  or (_23922_, _23921_, _23918_);
  and (_23923_, _23922_, _03704_);
  nor (_23924_, _23841_, _03704_);
  or (_23926_, _23924_, _23923_);
  and (_23927_, _23926_, _03385_);
  nor (_23928_, _23858_, _03385_);
  or (_23929_, _23928_, _23927_);
  and (_23930_, _23929_, _03702_);
  and (_23931_, _12596_, _05347_);
  nor (_23932_, _23931_, _23827_);
  nor (_23933_, _23932_, _03702_);
  or (_23934_, _23933_, _23930_);
  or (_23935_, _23934_, _42912_);
  or (_23936_, _42908_, \oc8051_golden_model_1.IP [2]);
  and (_23937_, _23936_, _41654_);
  and (_43244_, _23937_, _23935_);
  and (_23938_, _09696_, \oc8051_golden_model_1.IP [3]);
  nor (_23939_, _09696_, _05050_);
  or (_23940_, _23939_, _23938_);
  or (_23941_, _23940_, _06994_);
  nor (_23942_, _12610_, _09696_);
  or (_23943_, _23942_, _23938_);
  or (_23944_, _23943_, _04630_);
  and (_23946_, _05347_, \oc8051_golden_model_1.ACC [3]);
  or (_23947_, _23946_, _23938_);
  and (_23948_, _23947_, _04615_);
  and (_23949_, _04616_, \oc8051_golden_model_1.IP [3]);
  or (_23950_, _23949_, _03757_);
  or (_23951_, _23950_, _23948_);
  and (_23952_, _23951_, _03697_);
  and (_23953_, _23952_, _23944_);
  and (_23954_, _09709_, \oc8051_golden_model_1.IP [3]);
  and (_23955_, _12619_, _06089_);
  or (_23957_, _23955_, _23954_);
  and (_23958_, _23957_, _03696_);
  or (_23959_, _23958_, _03755_);
  or (_23960_, _23959_, _23953_);
  or (_23961_, _23940_, _04537_);
  and (_23962_, _23961_, _23960_);
  or (_23963_, _23962_, _03750_);
  or (_23964_, _23947_, _03751_);
  and (_23965_, _23964_, _03692_);
  and (_23966_, _23965_, _23963_);
  and (_23968_, _12622_, _06089_);
  or (_23969_, _23968_, _23954_);
  and (_23970_, _23969_, _03691_);
  or (_23971_, _23970_, _03684_);
  or (_23972_, _23971_, _23966_);
  or (_23973_, _23954_, _12618_);
  and (_23974_, _23973_, _23957_);
  or (_23975_, _23974_, _03685_);
  and (_23976_, _23975_, _03680_);
  and (_23977_, _23976_, _23972_);
  nor (_23979_, _12665_, _09709_);
  or (_23980_, _23979_, _23954_);
  and (_23981_, _23980_, _03679_);
  or (_23982_, _23981_, _07544_);
  or (_23983_, _23982_, _23977_);
  and (_23984_, _23983_, _23941_);
  or (_23985_, _23984_, _04678_);
  and (_23986_, _06937_, _05347_);
  or (_23987_, _23938_, _04679_);
  or (_23988_, _23987_, _23986_);
  and (_23990_, _23988_, _03415_);
  and (_23991_, _23990_, _23985_);
  nor (_23992_, _12724_, _09696_);
  or (_23993_, _23938_, _23992_);
  and (_23994_, _23993_, _07559_);
  or (_23995_, _23994_, _23991_);
  or (_23996_, _23995_, _08854_);
  and (_23997_, _12738_, _05347_);
  or (_23998_, _23938_, _04703_);
  or (_23999_, _23998_, _23997_);
  and (_24000_, _05347_, _06415_);
  or (_24001_, _24000_, _23938_);
  or (_24002_, _24001_, _04694_);
  and (_24003_, _24002_, _04701_);
  and (_24004_, _24003_, _23999_);
  and (_24005_, _24004_, _23996_);
  and (_24006_, _10455_, _05347_);
  or (_24007_, _24006_, _23938_);
  and (_24008_, _24007_, _03959_);
  or (_24009_, _24008_, _24005_);
  and (_24011_, _24009_, _04708_);
  or (_24012_, _23938_, _05554_);
  and (_24013_, _24001_, _03866_);
  and (_24014_, _24013_, _24012_);
  or (_24015_, _24014_, _24011_);
  and (_24016_, _24015_, _04706_);
  and (_24017_, _23947_, _03967_);
  and (_24018_, _24017_, _24012_);
  or (_24019_, _24018_, _03835_);
  or (_24020_, _24019_, _24016_);
  nor (_24022_, _12737_, _09696_);
  or (_24023_, _23938_, _06532_);
  or (_24024_, _24023_, _24022_);
  and (_24025_, _24024_, _06537_);
  and (_24026_, _24025_, _24020_);
  nor (_24027_, _08701_, _09696_);
  or (_24028_, _24027_, _23938_);
  and (_24029_, _24028_, _03954_);
  or (_24030_, _24029_, _03703_);
  or (_24031_, _24030_, _24026_);
  or (_24033_, _23943_, _03704_);
  and (_24034_, _24033_, _03385_);
  and (_24035_, _24034_, _24031_);
  and (_24036_, _23969_, _03384_);
  or (_24037_, _24036_, _03701_);
  or (_24038_, _24037_, _24035_);
  and (_24039_, _12792_, _05347_);
  or (_24040_, _24039_, _23938_);
  or (_24041_, _24040_, _03702_);
  and (_24042_, _24041_, _24038_);
  or (_24044_, _24042_, _42912_);
  or (_24045_, _42908_, \oc8051_golden_model_1.IP [3]);
  and (_24046_, _24045_, _41654_);
  and (_43245_, _24046_, _24044_);
  and (_24047_, _09696_, \oc8051_golden_model_1.IP [4]);
  nor (_24048_, _05898_, _09696_);
  or (_24049_, _24048_, _24047_);
  or (_24050_, _24049_, _06994_);
  and (_24051_, _09709_, \oc8051_golden_model_1.IP [4]);
  and (_24052_, _12808_, _06089_);
  or (_24054_, _24052_, _24051_);
  and (_24055_, _24054_, _03691_);
  nor (_24056_, _12828_, _09696_);
  or (_24057_, _24056_, _24047_);
  or (_24058_, _24057_, _04630_);
  and (_24059_, _05347_, \oc8051_golden_model_1.ACC [4]);
  or (_24060_, _24059_, _24047_);
  and (_24061_, _24060_, _04615_);
  and (_24062_, _04616_, \oc8051_golden_model_1.IP [4]);
  or (_24063_, _24062_, _03757_);
  or (_24065_, _24063_, _24061_);
  and (_24066_, _24065_, _03697_);
  and (_24067_, _24066_, _24058_);
  and (_24068_, _12832_, _06089_);
  or (_24069_, _24068_, _24051_);
  and (_24070_, _24069_, _03696_);
  or (_24071_, _24070_, _03755_);
  or (_24072_, _24071_, _24067_);
  or (_24073_, _24049_, _04537_);
  and (_24074_, _24073_, _24072_);
  or (_24076_, _24074_, _03750_);
  or (_24077_, _24060_, _03751_);
  and (_24078_, _24077_, _03692_);
  and (_24079_, _24078_, _24076_);
  or (_24080_, _24079_, _24055_);
  and (_24081_, _24080_, _03685_);
  or (_24082_, _24051_, _12847_);
  and (_24083_, _24082_, _03684_);
  and (_24084_, _24083_, _24069_);
  or (_24085_, _24084_, _24081_);
  and (_24088_, _24085_, _03680_);
  nor (_24089_, _12810_, _09709_);
  or (_24090_, _24089_, _24051_);
  and (_24091_, _24090_, _03679_);
  or (_24092_, _24091_, _07544_);
  or (_24093_, _24092_, _24088_);
  and (_24094_, _24093_, _24050_);
  or (_24095_, _24094_, _04678_);
  and (_24096_, _06942_, _05347_);
  or (_24097_, _24047_, _04679_);
  or (_24100_, _24097_, _24096_);
  and (_24101_, _24100_, _03415_);
  and (_24102_, _24101_, _24095_);
  nor (_24103_, _12919_, _09696_);
  or (_24104_, _24103_, _24047_);
  and (_24105_, _24104_, _07559_);
  or (_24106_, _24105_, _08854_);
  or (_24107_, _24106_, _24102_);
  and (_24108_, _12933_, _05347_);
  or (_24109_, _24047_, _04703_);
  or (_24112_, _24109_, _24108_);
  and (_24113_, _06422_, _05347_);
  or (_24114_, _24113_, _24047_);
  or (_24115_, _24114_, _04694_);
  and (_24116_, _24115_, _04701_);
  and (_24117_, _24116_, _24112_);
  and (_24118_, _24117_, _24107_);
  and (_24119_, _08700_, _05347_);
  or (_24120_, _24119_, _24047_);
  and (_24121_, _24120_, _03959_);
  or (_24124_, _24121_, _24118_);
  and (_24125_, _24124_, _04708_);
  or (_24126_, _24047_, _08303_);
  and (_24127_, _24114_, _03866_);
  and (_24128_, _24127_, _24126_);
  or (_24129_, _24128_, _24125_);
  and (_24130_, _24129_, _04706_);
  and (_24131_, _24060_, _03967_);
  and (_24132_, _24131_, _24126_);
  or (_24133_, _24132_, _03835_);
  or (_24136_, _24133_, _24130_);
  nor (_24137_, _12931_, _09696_);
  or (_24138_, _24047_, _06532_);
  or (_24139_, _24138_, _24137_);
  and (_24140_, _24139_, _06537_);
  and (_24141_, _24140_, _24136_);
  nor (_24142_, _08699_, _09696_);
  or (_24143_, _24142_, _24047_);
  and (_24144_, _24143_, _03954_);
  or (_24145_, _24144_, _03703_);
  or (_24147_, _24145_, _24141_);
  or (_24148_, _24057_, _03704_);
  and (_24149_, _24148_, _03385_);
  and (_24150_, _24149_, _24147_);
  and (_24151_, _24054_, _03384_);
  or (_24152_, _24151_, _03701_);
  or (_24153_, _24152_, _24150_);
  and (_24154_, _12991_, _05347_);
  or (_24155_, _24154_, _24047_);
  or (_24156_, _24155_, _03702_);
  and (_24158_, _24156_, _24153_);
  or (_24159_, _24158_, _42912_);
  or (_24160_, _42908_, \oc8051_golden_model_1.IP [4]);
  and (_24161_, _24160_, _41654_);
  and (_43246_, _24161_, _24159_);
  and (_24162_, _09696_, \oc8051_golden_model_1.IP [5]);
  nor (_24163_, _13025_, _09696_);
  or (_24164_, _24163_, _24162_);
  or (_24165_, _24164_, _04630_);
  and (_24166_, _05347_, \oc8051_golden_model_1.ACC [5]);
  or (_24168_, _24166_, _24162_);
  and (_24169_, _24168_, _04615_);
  and (_24170_, _04616_, \oc8051_golden_model_1.IP [5]);
  or (_24171_, _24170_, _03757_);
  or (_24172_, _24171_, _24169_);
  and (_24173_, _24172_, _03697_);
  and (_24174_, _24173_, _24165_);
  and (_24175_, _09709_, \oc8051_golden_model_1.IP [5]);
  and (_24176_, _13029_, _06089_);
  or (_24177_, _24176_, _24175_);
  and (_24179_, _24177_, _03696_);
  or (_24180_, _24179_, _03755_);
  or (_24181_, _24180_, _24174_);
  nor (_24182_, _05799_, _09696_);
  or (_24183_, _24182_, _24162_);
  or (_24184_, _24183_, _04537_);
  and (_24185_, _24184_, _24181_);
  or (_24186_, _24185_, _03750_);
  or (_24187_, _24168_, _03751_);
  and (_24188_, _24187_, _03692_);
  and (_24190_, _24188_, _24186_);
  and (_24191_, _13007_, _06089_);
  or (_24192_, _24191_, _24175_);
  and (_24193_, _24192_, _03691_);
  or (_24194_, _24193_, _03684_);
  or (_24195_, _24194_, _24190_);
  or (_24196_, _24175_, _13044_);
  and (_24197_, _24196_, _24177_);
  or (_24198_, _24197_, _03685_);
  and (_24199_, _24198_, _03680_);
  and (_24200_, _24199_, _24195_);
  nor (_24201_, _13009_, _09709_);
  or (_24202_, _24201_, _24175_);
  and (_24203_, _24202_, _03679_);
  or (_24204_, _24203_, _07544_);
  or (_24205_, _24204_, _24200_);
  or (_24206_, _24183_, _06994_);
  and (_24207_, _24206_, _24205_);
  or (_24208_, _24207_, _04678_);
  and (_24209_, _06941_, _05347_);
  or (_24211_, _24162_, _04679_);
  or (_24212_, _24211_, _24209_);
  and (_24213_, _24212_, _03415_);
  and (_24214_, _24213_, _24208_);
  nor (_24215_, _13118_, _09696_);
  or (_24216_, _24215_, _24162_);
  and (_24217_, _24216_, _07559_);
  or (_24218_, _24217_, _08854_);
  or (_24219_, _24218_, _24214_);
  and (_24220_, _13133_, _05347_);
  or (_24222_, _24162_, _04703_);
  or (_24223_, _24222_, _24220_);
  and (_24224_, _06371_, _05347_);
  or (_24225_, _24224_, _24162_);
  or (_24226_, _24225_, _04694_);
  and (_24227_, _24226_, _04701_);
  and (_24228_, _24227_, _24223_);
  and (_24229_, _24228_, _24219_);
  and (_24230_, _10451_, _05347_);
  or (_24231_, _24230_, _24162_);
  and (_24233_, _24231_, _03959_);
  or (_24234_, _24233_, _24229_);
  and (_24235_, _24234_, _04708_);
  or (_24236_, _24162_, _08302_);
  and (_24237_, _24225_, _03866_);
  and (_24238_, _24237_, _24236_);
  or (_24239_, _24238_, _24235_);
  and (_24240_, _24239_, _04706_);
  and (_24241_, _24168_, _03967_);
  and (_24242_, _24241_, _24236_);
  or (_24244_, _24242_, _03835_);
  or (_24245_, _24244_, _24240_);
  nor (_24246_, _13131_, _09696_);
  or (_24247_, _24162_, _06532_);
  or (_24248_, _24247_, _24246_);
  and (_24249_, _24248_, _06537_);
  and (_24250_, _24249_, _24245_);
  nor (_24251_, _08697_, _09696_);
  or (_24252_, _24251_, _24162_);
  and (_24253_, _24252_, _03954_);
  or (_24255_, _24253_, _03703_);
  or (_24256_, _24255_, _24250_);
  or (_24257_, _24164_, _03704_);
  and (_24258_, _24257_, _03385_);
  and (_24259_, _24258_, _24256_);
  and (_24260_, _24192_, _03384_);
  or (_24261_, _24260_, _03701_);
  or (_24262_, _24261_, _24259_);
  and (_24263_, _13193_, _05347_);
  or (_24264_, _24263_, _24162_);
  or (_24266_, _24264_, _03702_);
  and (_24267_, _24266_, _24262_);
  or (_24268_, _24267_, _42912_);
  or (_24269_, _42908_, \oc8051_golden_model_1.IP [5]);
  and (_24270_, _24269_, _41654_);
  and (_43247_, _24270_, _24268_);
  and (_24271_, _09696_, \oc8051_golden_model_1.IP [6]);
  nor (_24272_, _06013_, _09696_);
  or (_24273_, _24272_, _24271_);
  or (_24274_, _24273_, _06994_);
  and (_24276_, _09709_, \oc8051_golden_model_1.IP [6]);
  and (_24277_, _13218_, _06089_);
  or (_24278_, _24277_, _24276_);
  and (_24279_, _24278_, _03691_);
  nor (_24280_, _13234_, _09696_);
  or (_24281_, _24280_, _24271_);
  or (_24282_, _24281_, _04630_);
  and (_24283_, _05347_, \oc8051_golden_model_1.ACC [6]);
  or (_24284_, _24283_, _24271_);
  and (_24285_, _24284_, _04615_);
  and (_24286_, _04616_, \oc8051_golden_model_1.IP [6]);
  or (_24287_, _24286_, _03757_);
  or (_24288_, _24287_, _24285_);
  and (_24289_, _24288_, _03697_);
  and (_24290_, _24289_, _24282_);
  and (_24291_, _13238_, _06089_);
  or (_24292_, _24291_, _24276_);
  and (_24293_, _24292_, _03696_);
  or (_24294_, _24293_, _03755_);
  or (_24295_, _24294_, _24290_);
  or (_24297_, _24273_, _04537_);
  and (_24298_, _24297_, _24295_);
  or (_24299_, _24298_, _03750_);
  or (_24300_, _24284_, _03751_);
  and (_24301_, _24300_, _03692_);
  and (_24302_, _24301_, _24299_);
  or (_24303_, _24302_, _24279_);
  and (_24304_, _24303_, _03685_);
  or (_24305_, _24276_, _13253_);
  and (_24306_, _24305_, _03684_);
  and (_24308_, _24306_, _24292_);
  or (_24309_, _24308_, _24304_);
  and (_24310_, _24309_, _03680_);
  nor (_24311_, _13220_, _09709_);
  or (_24312_, _24311_, _24276_);
  and (_24313_, _24312_, _03679_);
  or (_24314_, _24313_, _07544_);
  or (_24315_, _24314_, _24310_);
  and (_24316_, _24315_, _24274_);
  or (_24317_, _24316_, _04678_);
  and (_24319_, _06933_, _05347_);
  or (_24320_, _24271_, _04679_);
  or (_24321_, _24320_, _24319_);
  and (_24322_, _24321_, _03415_);
  and (_24323_, _24322_, _24317_);
  nor (_24324_, _13326_, _09696_);
  or (_24325_, _24324_, _24271_);
  and (_24326_, _24325_, _07559_);
  or (_24327_, _24326_, _08854_);
  or (_24328_, _24327_, _24323_);
  and (_24330_, _13341_, _05347_);
  or (_24331_, _24271_, _04703_);
  or (_24332_, _24331_, _24330_);
  and (_24333_, _13333_, _05347_);
  or (_24334_, _24333_, _24271_);
  or (_24335_, _24334_, _04694_);
  and (_24336_, _24335_, _04701_);
  and (_24337_, _24336_, _24332_);
  and (_24338_, _24337_, _24328_);
  and (_24339_, _08695_, _05347_);
  or (_24341_, _24339_, _24271_);
  and (_24342_, _24341_, _03959_);
  or (_24343_, _24342_, _24338_);
  and (_24344_, _24343_, _04708_);
  or (_24345_, _24271_, _08289_);
  and (_24346_, _24334_, _03866_);
  and (_24347_, _24346_, _24345_);
  or (_24348_, _24347_, _24344_);
  and (_24349_, _24348_, _04706_);
  and (_24350_, _24284_, _03967_);
  and (_24351_, _24350_, _24345_);
  or (_24352_, _24351_, _03835_);
  or (_24353_, _24352_, _24349_);
  nor (_24354_, _13340_, _09696_);
  or (_24355_, _24271_, _06532_);
  or (_24356_, _24355_, _24354_);
  and (_24357_, _24356_, _06537_);
  and (_24358_, _24357_, _24353_);
  nor (_24359_, _08694_, _09696_);
  or (_24360_, _24359_, _24271_);
  and (_24362_, _24360_, _03954_);
  or (_24363_, _24362_, _03703_);
  or (_24364_, _24363_, _24358_);
  or (_24365_, _24281_, _03704_);
  and (_24366_, _24365_, _03385_);
  and (_24367_, _24366_, _24364_);
  and (_24368_, _24278_, _03384_);
  or (_24369_, _24368_, _03701_);
  or (_24370_, _24369_, _24367_);
  nor (_24371_, _13399_, _09696_);
  or (_24373_, _24371_, _24271_);
  or (_24374_, _24373_, _03702_);
  and (_24375_, _24374_, _24370_);
  or (_24376_, _24375_, _42912_);
  or (_24377_, _42908_, \oc8051_golden_model_1.IP [6]);
  and (_24378_, _24377_, _41654_);
  and (_43248_, _24378_, _24376_);
  not (_24379_, \oc8051_golden_model_1.DPL [0]);
  nor (_24380_, _42908_, _24379_);
  nor (_24381_, _05545_, _24379_);
  and (_24383_, _05440_, _04608_);
  or (_24384_, _24383_, _24381_);
  or (_24385_, _24384_, _06994_);
  and (_24386_, _05545_, \oc8051_golden_model_1.ACC [0]);
  or (_24387_, _24386_, _24381_);
  or (_24388_, _24387_, _03751_);
  nor (_24389_, _05652_, _09802_);
  or (_24390_, _24389_, _24381_);
  or (_24391_, _24390_, _04630_);
  and (_24392_, _24387_, _04615_);
  nor (_24394_, _04615_, _24379_);
  or (_24395_, _24394_, _03757_);
  or (_24396_, _24395_, _24392_);
  and (_24397_, _24396_, _04537_);
  and (_24398_, _24397_, _24391_);
  and (_24399_, _24384_, _03755_);
  or (_24400_, _24399_, _03750_);
  or (_24401_, _24400_, _24398_);
  and (_24402_, _24401_, _24388_);
  or (_24403_, _24402_, _09821_);
  nand (_24405_, _09821_, \oc8051_golden_model_1.DPL [0]);
  and (_24406_, _24405_, _09806_);
  and (_24407_, _24406_, _24403_);
  nor (_24408_, _04326_, _09806_);
  or (_24409_, _24408_, _07544_);
  or (_24410_, _24409_, _24407_);
  and (_24411_, _24410_, _24385_);
  or (_24412_, _24411_, _04678_);
  or (_24413_, _24381_, _04679_);
  and (_24414_, _06935_, _05545_);
  or (_24416_, _24414_, _24413_);
  and (_24417_, _24416_, _24412_);
  or (_24418_, _24417_, _07559_);
  nor (_24419_, _12119_, _09802_);
  or (_24420_, _24381_, _03415_);
  or (_24421_, _24420_, _24419_);
  and (_24422_, _24421_, _04694_);
  and (_24423_, _24422_, _24418_);
  and (_24424_, _05545_, _06428_);
  or (_24425_, _24424_, _24381_);
  and (_24427_, _24425_, _03839_);
  or (_24428_, _24427_, _03838_);
  or (_24429_, _24428_, _24423_);
  and (_24430_, _12133_, _05545_);
  or (_24431_, _24430_, _24381_);
  or (_24432_, _24431_, _04703_);
  and (_24433_, _24432_, _04701_);
  and (_24434_, _24433_, _24429_);
  nor (_24435_, _10458_, _09802_);
  or (_24436_, _24435_, _24381_);
  and (_24438_, _24386_, _05652_);
  nor (_24439_, _24438_, _04701_);
  and (_24440_, _24439_, _24436_);
  or (_24441_, _24440_, _24434_);
  and (_24442_, _24441_, _04708_);
  nand (_24443_, _24425_, _03866_);
  nor (_24444_, _24443_, _24389_);
  or (_24445_, _24444_, _03967_);
  or (_24446_, _24445_, _24442_);
  or (_24447_, _24438_, _24381_);
  or (_24449_, _24447_, _04706_);
  and (_24450_, _24449_, _24446_);
  or (_24451_, _24450_, _03835_);
  nor (_24452_, _12132_, _09802_);
  or (_24453_, _24381_, _06532_);
  or (_24454_, _24453_, _24452_);
  and (_24455_, _24454_, _06537_);
  and (_24456_, _24455_, _24451_);
  and (_24457_, _24436_, _03954_);
  or (_24458_, _24457_, _17066_);
  or (_24460_, _24458_, _24456_);
  or (_24461_, _24390_, _04170_);
  and (_24462_, _24461_, _42908_);
  and (_24463_, _24462_, _24460_);
  or (_24464_, _24463_, _24380_);
  and (_43251_, _24464_, _41654_);
  and (_24465_, _42912_, \oc8051_golden_model_1.DPL [1]);
  nor (_24466_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_24467_, _24466_, _09826_);
  and (_24468_, _24467_, _09821_);
  or (_24470_, _05545_, \oc8051_golden_model_1.DPL [1]);
  and (_24471_, _12225_, _05440_);
  not (_24472_, _24471_);
  and (_24473_, _24472_, _24470_);
  or (_24474_, _24473_, _04630_);
  and (_24475_, _09848_, \oc8051_golden_model_1.DPL [1]);
  and (_24476_, _05545_, \oc8051_golden_model_1.ACC [1]);
  or (_24477_, _24476_, _24475_);
  and (_24478_, _24477_, _04615_);
  and (_24479_, _04616_, \oc8051_golden_model_1.DPL [1]);
  or (_24481_, _24479_, _03757_);
  or (_24482_, _24481_, _24478_);
  and (_24483_, _24482_, _04537_);
  and (_24484_, _24483_, _24474_);
  and (_24485_, _05440_, _04813_);
  or (_24486_, _24485_, _24475_);
  and (_24487_, _24486_, _03755_);
  or (_24488_, _24487_, _03750_);
  or (_24489_, _24488_, _24484_);
  or (_24490_, _24477_, _03751_);
  and (_24492_, _24490_, _09822_);
  and (_24493_, _24492_, _24489_);
  or (_24494_, _24493_, _24468_);
  and (_24495_, _24494_, _09806_);
  nor (_24496_, _04515_, _09806_);
  or (_24497_, _24496_, _07544_);
  or (_24498_, _24497_, _24495_);
  or (_24499_, _24486_, _06994_);
  and (_24500_, _24499_, _24498_);
  or (_24501_, _24500_, _04678_);
  and (_24504_, _06934_, _05545_);
  or (_24505_, _24475_, _04679_);
  or (_24506_, _24505_, _24504_);
  and (_24507_, _24506_, _03415_);
  and (_24508_, _24507_, _24501_);
  and (_24509_, _24470_, _07559_);
  nand (_24510_, _12313_, _05440_);
  and (_24511_, _24510_, _24509_);
  or (_24512_, _24511_, _24508_);
  and (_24513_, _24512_, _03840_);
  or (_24515_, _12207_, _09802_);
  and (_24516_, _24515_, _03838_);
  nand (_24517_, _05440_, _04515_);
  and (_24518_, _24517_, _03839_);
  or (_24519_, _24518_, _24516_);
  and (_24520_, _24519_, _24470_);
  or (_24521_, _24520_, _03959_);
  or (_24522_, _24521_, _24513_);
  nor (_24523_, _08710_, _09802_);
  or (_24524_, _24523_, _24475_);
  nand (_24526_, _08709_, _05440_);
  and (_24527_, _24526_, _24524_);
  or (_24528_, _24527_, _04701_);
  and (_24529_, _24528_, _04708_);
  and (_24530_, _24529_, _24522_);
  or (_24531_, _12206_, _09802_);
  and (_24532_, _24470_, _03866_);
  and (_24533_, _24532_, _24531_);
  or (_24534_, _24533_, _03967_);
  or (_24535_, _24534_, _24530_);
  nor (_24537_, _24475_, _04706_);
  nand (_24538_, _24537_, _24526_);
  and (_24539_, _24538_, _06532_);
  and (_24540_, _24539_, _24535_);
  or (_24541_, _24517_, _05603_);
  and (_24542_, _24470_, _03835_);
  and (_24543_, _24542_, _24541_);
  or (_24544_, _24543_, _03954_);
  or (_24545_, _24544_, _24540_);
  or (_24546_, _24524_, _06537_);
  and (_24548_, _24546_, _03704_);
  and (_24549_, _24548_, _24545_);
  and (_24550_, _24473_, _03703_);
  or (_24551_, _24550_, _03701_);
  or (_24552_, _24551_, _24549_);
  or (_24553_, _24475_, _03702_);
  or (_24554_, _24553_, _24471_);
  and (_24555_, _24554_, _42908_);
  and (_24556_, _24555_, _24552_);
  or (_24557_, _24556_, _24465_);
  and (_43252_, _24557_, _41654_);
  or (_24559_, _42908_, \oc8051_golden_model_1.DPL [2]);
  and (_24560_, _24559_, _41654_);
  and (_24561_, _09848_, \oc8051_golden_model_1.DPL [2]);
  nor (_24562_, _09802_, _05236_);
  or (_24563_, _24562_, _24561_);
  or (_24564_, _24563_, _06994_);
  nor (_24565_, _09826_, \oc8051_golden_model_1.DPL [2]);
  nor (_24566_, _24565_, _09827_);
  and (_24567_, _24566_, _09821_);
  nor (_24569_, _12427_, _09802_);
  or (_24570_, _24569_, _24561_);
  or (_24571_, _24570_, _04630_);
  and (_24572_, _05545_, \oc8051_golden_model_1.ACC [2]);
  or (_24573_, _24572_, _24561_);
  and (_24574_, _24573_, _04615_);
  and (_24575_, _04616_, \oc8051_golden_model_1.DPL [2]);
  or (_24576_, _24575_, _03757_);
  or (_24577_, _24576_, _24574_);
  and (_24578_, _24577_, _04537_);
  and (_24580_, _24578_, _24571_);
  and (_24581_, _24563_, _03755_);
  or (_24582_, _24581_, _03750_);
  or (_24583_, _24582_, _24580_);
  or (_24584_, _24573_, _03751_);
  and (_24585_, _24584_, _09822_);
  and (_24586_, _24585_, _24583_);
  or (_24587_, _24586_, _24567_);
  and (_24588_, _24587_, _09806_);
  nor (_24589_, _04077_, _09806_);
  or (_24591_, _24589_, _07544_);
  or (_24592_, _24591_, _24588_);
  and (_24593_, _24592_, _24564_);
  or (_24594_, _24593_, _04678_);
  or (_24595_, _24561_, _04679_);
  and (_24596_, _06938_, _05545_);
  or (_24597_, _24596_, _24595_);
  and (_24598_, _24597_, _03415_);
  and (_24599_, _24598_, _24594_);
  nor (_24600_, _12523_, _09848_);
  or (_24602_, _24600_, _24561_);
  and (_24603_, _24602_, _07559_);
  or (_24604_, _24603_, _24599_);
  or (_24605_, _24604_, _08854_);
  and (_24606_, _12537_, _05440_);
  or (_24607_, _24561_, _04703_);
  or (_24608_, _24607_, _24606_);
  and (_24609_, _05545_, _06457_);
  or (_24610_, _24609_, _24561_);
  or (_24611_, _24610_, _04694_);
  and (_24613_, _24611_, _04701_);
  and (_24614_, _24613_, _24608_);
  and (_24615_, _24614_, _24605_);
  and (_24616_, _08707_, _05545_);
  or (_24617_, _24616_, _24561_);
  and (_24618_, _24617_, _03959_);
  or (_24619_, _24618_, _24615_);
  and (_24620_, _24619_, _04708_);
  or (_24621_, _24561_, _05700_);
  and (_24622_, _24610_, _03866_);
  and (_24624_, _24622_, _24621_);
  or (_24625_, _24624_, _24620_);
  and (_24626_, _24625_, _04706_);
  and (_24627_, _24573_, _03967_);
  and (_24628_, _24627_, _24621_);
  or (_24629_, _24628_, _03835_);
  or (_24630_, _24629_, _24626_);
  nor (_24631_, _12536_, _09802_);
  or (_24632_, _24561_, _06532_);
  or (_24633_, _24632_, _24631_);
  and (_24635_, _24633_, _06537_);
  and (_24636_, _24635_, _24630_);
  nor (_24637_, _08706_, _09802_);
  or (_24638_, _24637_, _24561_);
  and (_24639_, _24638_, _03954_);
  or (_24640_, _24639_, _03703_);
  or (_24641_, _24640_, _24636_);
  or (_24642_, _24570_, _03704_);
  and (_24643_, _24642_, _03702_);
  and (_24644_, _24643_, _24641_);
  and (_24646_, _12596_, _05440_);
  or (_24647_, _24646_, _24561_);
  and (_24648_, _24647_, _03701_);
  or (_24649_, _24648_, _42912_);
  or (_24650_, _24649_, _24644_);
  and (_43253_, _24650_, _24560_);
  or (_24651_, _42908_, \oc8051_golden_model_1.DPL [3]);
  and (_24652_, _24651_, _41654_);
  nor (_24653_, _09827_, \oc8051_golden_model_1.DPL [3]);
  nor (_24654_, _24653_, _09828_);
  and (_24656_, _24654_, _09821_);
  and (_24657_, _09848_, \oc8051_golden_model_1.DPL [3]);
  nor (_24658_, _12610_, _09802_);
  or (_24659_, _24658_, _24657_);
  or (_24660_, _24659_, _04630_);
  and (_24661_, _05545_, \oc8051_golden_model_1.ACC [3]);
  or (_24662_, _24661_, _24657_);
  and (_24663_, _24662_, _04615_);
  and (_24664_, _04616_, \oc8051_golden_model_1.DPL [3]);
  or (_24665_, _24664_, _03757_);
  or (_24667_, _24665_, _24663_);
  and (_24668_, _24667_, _04537_);
  and (_24669_, _24668_, _24660_);
  nor (_24670_, _09802_, _05050_);
  or (_24671_, _24670_, _24657_);
  and (_24672_, _24671_, _03755_);
  or (_24673_, _24672_, _03750_);
  or (_24674_, _24673_, _24669_);
  or (_24675_, _24662_, _03751_);
  and (_24676_, _24675_, _09822_);
  and (_24678_, _24676_, _24674_);
  or (_24679_, _24678_, _24656_);
  and (_24680_, _24679_, _09806_);
  nor (_24681_, _03946_, _09806_);
  or (_24682_, _24681_, _07544_);
  or (_24683_, _24682_, _24680_);
  or (_24684_, _24671_, _06994_);
  and (_24685_, _24684_, _24683_);
  or (_24686_, _24685_, _04678_);
  and (_24687_, _06937_, _05545_);
  or (_24689_, _24657_, _04679_);
  or (_24690_, _24689_, _24687_);
  and (_24691_, _24690_, _03415_);
  and (_24692_, _24691_, _24686_);
  nor (_24693_, _12724_, _09802_);
  or (_24694_, _24693_, _24657_);
  and (_24695_, _24694_, _07559_);
  or (_24696_, _24695_, _08854_);
  or (_24697_, _24696_, _24692_);
  and (_24698_, _12738_, _05440_);
  or (_24700_, _24657_, _04703_);
  or (_24701_, _24700_, _24698_);
  and (_24702_, _05545_, _06415_);
  or (_24703_, _24702_, _24657_);
  or (_24704_, _24703_, _04694_);
  and (_24705_, _24704_, _04701_);
  and (_24706_, _24705_, _24701_);
  and (_24707_, _24706_, _24697_);
  and (_24708_, _10455_, _05545_);
  or (_24709_, _24708_, _24657_);
  and (_24711_, _24709_, _03959_);
  or (_24712_, _24711_, _24707_);
  and (_24713_, _24712_, _04708_);
  or (_24714_, _24657_, _05554_);
  and (_24715_, _24703_, _03866_);
  and (_24716_, _24715_, _24714_);
  or (_24717_, _24716_, _24713_);
  and (_24718_, _24717_, _04706_);
  and (_24719_, _24662_, _03967_);
  and (_24720_, _24719_, _24714_);
  or (_24722_, _24720_, _03835_);
  or (_24723_, _24722_, _24718_);
  nor (_24724_, _12737_, _09802_);
  or (_24725_, _24657_, _06532_);
  or (_24726_, _24725_, _24724_);
  and (_24727_, _24726_, _06537_);
  and (_24728_, _24727_, _24723_);
  nor (_24729_, _08701_, _09802_);
  or (_24730_, _24729_, _24657_);
  and (_24731_, _24730_, _03954_);
  or (_24733_, _24731_, _03703_);
  or (_24734_, _24733_, _24728_);
  or (_24735_, _24659_, _03704_);
  and (_24736_, _24735_, _03702_);
  and (_24737_, _24736_, _24734_);
  and (_24738_, _12792_, _05440_);
  or (_24739_, _24738_, _24657_);
  and (_24740_, _24739_, _03701_);
  or (_24741_, _24740_, _42912_);
  or (_24742_, _24741_, _24737_);
  and (_43254_, _24742_, _24652_);
  or (_24744_, _42908_, \oc8051_golden_model_1.DPL [4]);
  and (_24745_, _24744_, _41654_);
  and (_24746_, _09848_, \oc8051_golden_model_1.DPL [4]);
  nor (_24747_, _05898_, _09802_);
  or (_24748_, _24747_, _24746_);
  or (_24749_, _24748_, _06994_);
  nor (_24750_, _12828_, _09802_);
  or (_24751_, _24750_, _24746_);
  or (_24752_, _24751_, _04630_);
  and (_24754_, _05545_, \oc8051_golden_model_1.ACC [4]);
  or (_24755_, _24754_, _24746_);
  and (_24756_, _24755_, _04615_);
  and (_24757_, _04616_, \oc8051_golden_model_1.DPL [4]);
  or (_24758_, _24757_, _03757_);
  or (_24759_, _24758_, _24756_);
  and (_24760_, _24759_, _04537_);
  and (_24761_, _24760_, _24752_);
  and (_24762_, _24748_, _03755_);
  or (_24763_, _24762_, _03750_);
  or (_24765_, _24763_, _24761_);
  or (_24766_, _24755_, _03751_);
  and (_24767_, _24766_, _09822_);
  and (_24768_, _24767_, _24765_);
  nor (_24769_, _09828_, \oc8051_golden_model_1.DPL [4]);
  nor (_24770_, _24769_, _09829_);
  and (_24771_, _24770_, _09821_);
  or (_24772_, _24771_, _24768_);
  and (_24773_, _24772_, _09806_);
  nor (_24774_, _06339_, _09806_);
  or (_24776_, _24774_, _07544_);
  or (_24777_, _24776_, _24773_);
  and (_24778_, _24777_, _24749_);
  or (_24779_, _24778_, _04678_);
  or (_24780_, _24746_, _04679_);
  and (_24781_, _06942_, _05545_);
  or (_24782_, _24781_, _24780_);
  and (_24783_, _24782_, _03415_);
  and (_24784_, _24783_, _24779_);
  nor (_24785_, _12919_, _09848_);
  or (_24787_, _24785_, _24746_);
  and (_24788_, _24787_, _07559_);
  or (_24789_, _24788_, _24784_);
  or (_24790_, _24789_, _08854_);
  and (_24791_, _12933_, _05440_);
  or (_24792_, _24746_, _04703_);
  or (_24793_, _24792_, _24791_);
  and (_24794_, _06422_, _05545_);
  or (_24795_, _24794_, _24746_);
  or (_24796_, _24795_, _04694_);
  and (_24798_, _24796_, _04701_);
  and (_24799_, _24798_, _24793_);
  and (_24800_, _24799_, _24790_);
  and (_24801_, _08700_, _05545_);
  or (_24802_, _24801_, _24746_);
  and (_24803_, _24802_, _03959_);
  or (_24804_, _24803_, _24800_);
  and (_24805_, _24804_, _04708_);
  or (_24806_, _24746_, _08303_);
  and (_24807_, _24795_, _03866_);
  and (_24809_, _24807_, _24806_);
  or (_24810_, _24809_, _24805_);
  and (_24811_, _24810_, _04706_);
  and (_24812_, _24755_, _03967_);
  and (_24813_, _24812_, _24806_);
  or (_24814_, _24813_, _03835_);
  or (_24815_, _24814_, _24811_);
  nor (_24816_, _12931_, _09802_);
  or (_24817_, _24746_, _06532_);
  or (_24818_, _24817_, _24816_);
  and (_24820_, _24818_, _06537_);
  and (_24821_, _24820_, _24815_);
  nor (_24822_, _08699_, _09802_);
  or (_24823_, _24822_, _24746_);
  and (_24824_, _24823_, _03954_);
  or (_24825_, _24824_, _03703_);
  or (_24826_, _24825_, _24821_);
  or (_24827_, _24751_, _03704_);
  and (_24828_, _24827_, _03702_);
  and (_24829_, _24828_, _24826_);
  and (_24831_, _12991_, _05440_);
  or (_24832_, _24831_, _24746_);
  and (_24833_, _24832_, _03701_);
  or (_24834_, _24833_, _42912_);
  or (_24835_, _24834_, _24829_);
  and (_43255_, _24835_, _24745_);
  and (_24836_, _42912_, \oc8051_golden_model_1.DPL [5]);
  and (_24837_, _09848_, \oc8051_golden_model_1.DPL [5]);
  nor (_24838_, _05799_, _09802_);
  or (_24839_, _24838_, _24837_);
  or (_24841_, _24839_, _06994_);
  nor (_24842_, _13025_, _09802_);
  or (_24843_, _24842_, _24837_);
  or (_24844_, _24843_, _04630_);
  and (_24845_, _05545_, \oc8051_golden_model_1.ACC [5]);
  or (_24846_, _24845_, _24837_);
  and (_24847_, _24846_, _04615_);
  and (_24848_, _04616_, \oc8051_golden_model_1.DPL [5]);
  or (_24849_, _24848_, _03757_);
  or (_24850_, _24849_, _24847_);
  and (_24852_, _24850_, _04537_);
  and (_24853_, _24852_, _24844_);
  and (_24854_, _24839_, _03755_);
  or (_24855_, _24854_, _03750_);
  or (_24856_, _24855_, _24853_);
  or (_24857_, _24846_, _03751_);
  and (_24858_, _24857_, _09822_);
  and (_24859_, _24858_, _24856_);
  nor (_24860_, _09829_, \oc8051_golden_model_1.DPL [5]);
  nor (_24861_, _24860_, _09830_);
  and (_24863_, _24861_, _09821_);
  or (_24864_, _24863_, _24859_);
  and (_24865_, _24864_, _09806_);
  nor (_24866_, _06370_, _09806_);
  or (_24867_, _24866_, _07544_);
  or (_24868_, _24867_, _24865_);
  and (_24869_, _24868_, _24841_);
  or (_24870_, _24869_, _04678_);
  or (_24871_, _24837_, _04679_);
  and (_24872_, _06941_, _05545_);
  or (_24874_, _24872_, _24871_);
  and (_24875_, _24874_, _03415_);
  and (_24876_, _24875_, _24870_);
  nor (_24877_, _13118_, _09848_);
  or (_24878_, _24877_, _24837_);
  and (_24879_, _24878_, _07559_);
  or (_24880_, _24879_, _24876_);
  or (_24881_, _24880_, _08854_);
  and (_24882_, _13133_, _05440_);
  or (_24883_, _24837_, _04703_);
  or (_24885_, _24883_, _24882_);
  and (_24886_, _06371_, _05545_);
  or (_24887_, _24886_, _24837_);
  or (_24888_, _24887_, _04694_);
  and (_24889_, _24888_, _04701_);
  and (_24890_, _24889_, _24885_);
  and (_24891_, _24890_, _24881_);
  and (_24892_, _10451_, _05545_);
  or (_24893_, _24892_, _24837_);
  and (_24894_, _24893_, _03959_);
  or (_24896_, _24894_, _24891_);
  and (_24897_, _24896_, _04708_);
  or (_24898_, _24837_, _08302_);
  and (_24899_, _24887_, _03866_);
  and (_24900_, _24899_, _24898_);
  or (_24901_, _24900_, _24897_);
  and (_24902_, _24901_, _04706_);
  and (_24903_, _24846_, _03967_);
  and (_24904_, _24903_, _24898_);
  or (_24905_, _24904_, _03835_);
  or (_24907_, _24905_, _24902_);
  nor (_24908_, _13131_, _09802_);
  or (_24909_, _24837_, _06532_);
  or (_24910_, _24909_, _24908_);
  and (_24911_, _24910_, _06537_);
  and (_24912_, _24911_, _24907_);
  nor (_24913_, _08697_, _09802_);
  or (_24914_, _24913_, _24837_);
  and (_24915_, _24914_, _03954_);
  or (_24916_, _24915_, _24912_);
  and (_24918_, _24916_, _03704_);
  and (_24919_, _24843_, _03703_);
  or (_24920_, _24919_, _03701_);
  or (_24921_, _24920_, _24918_);
  and (_24922_, _13193_, _05440_);
  or (_24923_, _24837_, _03702_);
  or (_24924_, _24923_, _24922_);
  and (_24925_, _24924_, _42908_);
  and (_24926_, _24925_, _24921_);
  or (_24927_, _24926_, _24836_);
  and (_43256_, _24927_, _41654_);
  or (_24929_, _42908_, \oc8051_golden_model_1.DPL [6]);
  and (_24930_, _24929_, _41654_);
  and (_24931_, _09848_, \oc8051_golden_model_1.DPL [6]);
  nor (_24932_, _06013_, _09802_);
  or (_24933_, _24932_, _24931_);
  or (_24934_, _24933_, _06994_);
  nor (_24935_, _13234_, _09802_);
  or (_24936_, _24935_, _24931_);
  or (_24937_, _24936_, _04630_);
  and (_24939_, _05545_, \oc8051_golden_model_1.ACC [6]);
  or (_24940_, _24939_, _24931_);
  and (_24941_, _24940_, _04615_);
  and (_24942_, _04616_, \oc8051_golden_model_1.DPL [6]);
  or (_24943_, _24942_, _03757_);
  or (_24944_, _24943_, _24941_);
  and (_24945_, _24944_, _04537_);
  and (_24946_, _24945_, _24937_);
  and (_24947_, _24933_, _03755_);
  or (_24948_, _24947_, _03750_);
  or (_24950_, _24948_, _24946_);
  or (_24951_, _24940_, _03751_);
  and (_24952_, _24951_, _09822_);
  and (_24953_, _24952_, _24950_);
  nor (_24954_, _09830_, \oc8051_golden_model_1.DPL [6]);
  nor (_24955_, _24954_, _09831_);
  and (_24956_, _24955_, _09821_);
  or (_24957_, _24956_, _24953_);
  and (_24958_, _24957_, _09806_);
  nor (_24959_, _06406_, _09806_);
  or (_24961_, _24959_, _07544_);
  or (_24962_, _24961_, _24958_);
  and (_24963_, _24962_, _24934_);
  or (_24964_, _24963_, _04678_);
  or (_24965_, _24931_, _04679_);
  and (_24966_, _06933_, _05545_);
  or (_24967_, _24966_, _24965_);
  and (_24968_, _24967_, _03415_);
  and (_24969_, _24968_, _24964_);
  nor (_24970_, _13326_, _09848_);
  or (_24972_, _24970_, _24931_);
  and (_24973_, _24972_, _07559_);
  or (_24974_, _24973_, _24969_);
  or (_24975_, _24974_, _08854_);
  and (_24976_, _13341_, _05440_);
  or (_24977_, _24931_, _04703_);
  or (_24978_, _24977_, _24976_);
  and (_24979_, _13333_, _05545_);
  or (_24980_, _24979_, _24931_);
  or (_24981_, _24980_, _04694_);
  and (_24982_, _24981_, _04701_);
  and (_24983_, _24982_, _24978_);
  and (_24984_, _24983_, _24975_);
  and (_24985_, _08695_, _05545_);
  or (_24986_, _24985_, _24931_);
  and (_24987_, _24986_, _03959_);
  or (_24988_, _24987_, _24984_);
  and (_24989_, _24988_, _04708_);
  or (_24990_, _24931_, _08289_);
  and (_24991_, _24980_, _03866_);
  and (_24994_, _24991_, _24990_);
  or (_24995_, _24994_, _24989_);
  and (_24996_, _24995_, _04706_);
  and (_24997_, _24940_, _03967_);
  and (_24998_, _24997_, _24990_);
  or (_24999_, _24998_, _03835_);
  or (_25000_, _24999_, _24996_);
  nor (_25001_, _13340_, _09802_);
  or (_25002_, _24931_, _06532_);
  or (_25003_, _25002_, _25001_);
  and (_25005_, _25003_, _06537_);
  and (_25006_, _25005_, _25000_);
  nor (_25007_, _08694_, _09802_);
  or (_25008_, _25007_, _24931_);
  and (_25009_, _25008_, _03954_);
  or (_25010_, _25009_, _03703_);
  or (_25011_, _25010_, _25006_);
  or (_25012_, _24936_, _03704_);
  and (_25013_, _25012_, _03702_);
  and (_25014_, _25013_, _25011_);
  nor (_25016_, _13399_, _09802_);
  or (_25017_, _25016_, _24931_);
  and (_25018_, _25017_, _03701_);
  or (_25019_, _25018_, _42912_);
  or (_25020_, _25019_, _25014_);
  and (_43257_, _25020_, _24930_);
  nor (_25021_, _42908_, _10545_);
  nand (_25022_, _08712_, _05422_);
  nor (_25023_, _05422_, _10545_);
  nor (_25024_, _25023_, _04706_);
  nand (_25025_, _25024_, _25022_);
  nor (_25026_, _09833_, \oc8051_golden_model_1.DPH [0]);
  nor (_25027_, _25026_, _09920_);
  and (_25028_, _25027_, _09821_);
  nor (_25029_, _05652_, _09899_);
  or (_25030_, _25029_, _25023_);
  or (_25031_, _25030_, _04630_);
  and (_25032_, _05422_, \oc8051_golden_model_1.ACC [0]);
  or (_25033_, _25032_, _25023_);
  and (_25034_, _25033_, _04615_);
  nor (_25037_, _04615_, _10545_);
  or (_25038_, _25037_, _03757_);
  or (_25039_, _25038_, _25034_);
  and (_25040_, _25039_, _04537_);
  and (_25041_, _25040_, _25031_);
  and (_25042_, _05422_, _04608_);
  or (_25043_, _25042_, _25023_);
  and (_25044_, _25043_, _03755_);
  or (_25045_, _25044_, _03750_);
  or (_25046_, _25045_, _25041_);
  or (_25048_, _25033_, _03751_);
  and (_25049_, _25048_, _09822_);
  and (_25050_, _25049_, _25046_);
  or (_25051_, _25050_, _25028_);
  and (_25052_, _25051_, _09806_);
  nor (_25053_, _04211_, _09806_);
  or (_25054_, _25053_, _07544_);
  or (_25055_, _25054_, _25052_);
  or (_25056_, _25043_, _06994_);
  and (_25057_, _25056_, _25055_);
  or (_25058_, _25057_, _04678_);
  and (_25059_, _06935_, _05422_);
  or (_25060_, _25023_, _04679_);
  or (_25061_, _25060_, _25059_);
  and (_25062_, _25061_, _25058_);
  or (_25063_, _25062_, _07559_);
  nor (_25064_, _12119_, _09899_);
  or (_25065_, _25023_, _03415_);
  or (_25066_, _25065_, _25064_);
  and (_25067_, _25066_, _04694_);
  and (_25070_, _25067_, _25063_);
  and (_25071_, _05422_, _06428_);
  or (_25072_, _25071_, _25023_);
  and (_25073_, _25072_, _03839_);
  or (_25074_, _25073_, _03838_);
  or (_25075_, _25074_, _25070_);
  and (_25076_, _12133_, _05422_);
  or (_25077_, _25076_, _25023_);
  or (_25078_, _25077_, _04703_);
  and (_25079_, _25078_, _04701_);
  and (_25081_, _25079_, _25075_);
  nor (_25082_, _10458_, _09899_);
  or (_25083_, _25082_, _25023_);
  and (_25084_, _25022_, _03959_);
  and (_25085_, _25084_, _25083_);
  or (_25086_, _25085_, _25081_);
  and (_25087_, _25086_, _04708_);
  nand (_25088_, _25072_, _03866_);
  nor (_25089_, _25088_, _25029_);
  or (_25090_, _25089_, _03967_);
  or (_25092_, _25090_, _25087_);
  and (_25093_, _25092_, _25025_);
  or (_25094_, _25093_, _03835_);
  nor (_25095_, _12132_, _09899_);
  or (_25096_, _25023_, _06532_);
  or (_25097_, _25096_, _25095_);
  and (_25098_, _25097_, _06537_);
  and (_25099_, _25098_, _25094_);
  and (_25100_, _25083_, _03954_);
  or (_25101_, _25100_, _17066_);
  or (_25103_, _25101_, _25099_);
  or (_25104_, _25030_, _04170_);
  and (_25105_, _25104_, _42908_);
  and (_25106_, _25105_, _25103_);
  or (_25107_, _25106_, _25021_);
  and (_43258_, _25107_, _41654_);
  or (_25108_, _42908_, \oc8051_golden_model_1.DPH [1]);
  and (_25109_, _25108_, _41654_);
  nor (_25110_, _09920_, \oc8051_golden_model_1.DPH [1]);
  nor (_25111_, _25110_, _09921_);
  and (_25112_, _25111_, _09821_);
  or (_25113_, _05422_, \oc8051_golden_model_1.DPH [1]);
  and (_25114_, _12225_, _05422_);
  not (_25115_, _25114_);
  and (_25116_, _25115_, _25113_);
  or (_25117_, _25116_, _04630_);
  not (_25118_, \oc8051_golden_model_1.DPH [1]);
  nor (_25119_, _05422_, _25118_);
  and (_25120_, _05422_, \oc8051_golden_model_1.ACC [1]);
  or (_25121_, _25120_, _25119_);
  and (_25124_, _25121_, _04615_);
  nor (_25125_, _04615_, _25118_);
  or (_25126_, _25125_, _03757_);
  or (_25127_, _25126_, _25124_);
  and (_25128_, _25127_, _04537_);
  and (_25129_, _25128_, _25117_);
  and (_25130_, _05422_, _04813_);
  or (_25131_, _25130_, _25119_);
  and (_25132_, _25131_, _03755_);
  or (_25133_, _25132_, _03750_);
  or (_25135_, _25133_, _25129_);
  or (_25136_, _25121_, _03751_);
  and (_25137_, _25136_, _09822_);
  and (_25138_, _25137_, _25135_);
  or (_25139_, _25138_, _25112_);
  and (_25140_, _25139_, _09806_);
  nor (_25141_, _04482_, _09806_);
  or (_25142_, _25141_, _07544_);
  or (_25143_, _25142_, _25140_);
  or (_25144_, _25131_, _06994_);
  and (_25146_, _25144_, _25143_);
  or (_25147_, _25146_, _04678_);
  and (_25148_, _06934_, _05422_);
  or (_25149_, _25119_, _04679_);
  or (_25150_, _25149_, _25148_);
  and (_25151_, _25150_, _03415_);
  and (_25152_, _25151_, _25147_);
  nor (_25153_, _12313_, _09899_);
  or (_25154_, _25153_, _25119_);
  and (_25155_, _25154_, _07559_);
  or (_25157_, _25155_, _25152_);
  and (_25158_, _25157_, _03840_);
  or (_25159_, _12207_, _09899_);
  and (_25160_, _25113_, _03838_);
  and (_25161_, _25160_, _25159_);
  nand (_25162_, _05422_, _04515_);
  and (_25163_, _25162_, _03839_);
  and (_25164_, _25163_, _25113_);
  or (_25165_, _25164_, _03959_);
  or (_25166_, _25165_, _25161_);
  or (_25168_, _25166_, _25158_);
  and (_25169_, _08711_, _05422_);
  or (_25170_, _25169_, _25119_);
  or (_25171_, _25170_, _04701_);
  and (_25172_, _25171_, _04708_);
  and (_25173_, _25172_, _25168_);
  or (_25174_, _12206_, _09899_);
  and (_25175_, _25113_, _03866_);
  and (_25176_, _25175_, _25174_);
  or (_25177_, _25176_, _03967_);
  or (_25179_, _25177_, _25173_);
  and (_25180_, _25120_, _05603_);
  or (_25181_, _25119_, _04706_);
  or (_25182_, _25181_, _25180_);
  and (_25183_, _25182_, _06532_);
  and (_25184_, _25183_, _25179_);
  or (_25185_, _25162_, _05603_);
  and (_25186_, _25185_, _03835_);
  and (_25187_, _25186_, _25113_);
  or (_25188_, _25187_, _03954_);
  or (_25190_, _25188_, _25184_);
  nor (_25191_, _08710_, _09899_);
  or (_25192_, _25191_, _25119_);
  or (_25193_, _25192_, _06537_);
  and (_25194_, _25193_, _25190_);
  or (_25195_, _25194_, _03703_);
  or (_25196_, _25116_, _03704_);
  and (_25197_, _25196_, _03702_);
  and (_25198_, _25197_, _25195_);
  or (_25199_, _25114_, _25119_);
  and (_25201_, _25199_, _03701_);
  or (_25202_, _25201_, _42912_);
  or (_25203_, _25202_, _25198_);
  and (_43259_, _25203_, _25109_);
  or (_25204_, _42908_, \oc8051_golden_model_1.DPH [2]);
  and (_25205_, _25204_, _41654_);
  not (_25206_, \oc8051_golden_model_1.DPH [2]);
  nor (_25207_, _05422_, _25206_);
  nor (_25208_, _09899_, _05236_);
  or (_25209_, _25208_, _25207_);
  or (_25211_, _25209_, _06994_);
  or (_25212_, _09921_, \oc8051_golden_model_1.DPH [2]);
  nor (_25213_, _09922_, _09822_);
  and (_25214_, _25213_, _25212_);
  nor (_25215_, _12427_, _09899_);
  or (_25216_, _25215_, _25207_);
  or (_25217_, _25216_, _04630_);
  and (_25218_, _05422_, \oc8051_golden_model_1.ACC [2]);
  or (_25219_, _25218_, _25207_);
  and (_25220_, _25219_, _04615_);
  nor (_25222_, _04615_, _25206_);
  or (_25223_, _25222_, _03757_);
  or (_25224_, _25223_, _25220_);
  and (_25225_, _25224_, _04537_);
  and (_25226_, _25225_, _25217_);
  and (_25227_, _25209_, _03755_);
  or (_25228_, _25227_, _03750_);
  or (_25229_, _25228_, _25226_);
  or (_25230_, _25219_, _03751_);
  and (_25231_, _25230_, _09822_);
  and (_25233_, _25231_, _25229_);
  or (_25234_, _25233_, _25214_);
  and (_25235_, _25234_, _09806_);
  nor (_25236_, _04165_, _09806_);
  or (_25237_, _25236_, _07544_);
  or (_25238_, _25237_, _25235_);
  and (_25239_, _25238_, _25211_);
  or (_25240_, _25239_, _04678_);
  and (_25241_, _06938_, _05422_);
  or (_25242_, _25207_, _04679_);
  or (_25243_, _25242_, _25241_);
  and (_25244_, _25243_, _03415_);
  and (_25245_, _25244_, _25240_);
  nor (_25246_, _12523_, _09899_);
  or (_25247_, _25246_, _25207_);
  and (_25248_, _25247_, _07559_);
  or (_25249_, _25248_, _25245_);
  or (_25250_, _25249_, _08854_);
  and (_25251_, _12537_, _05422_);
  or (_25252_, _25207_, _04703_);
  or (_25255_, _25252_, _25251_);
  and (_25256_, _05422_, _06457_);
  or (_25257_, _25256_, _25207_);
  or (_25258_, _25257_, _04694_);
  and (_25259_, _25258_, _04701_);
  and (_25260_, _25259_, _25255_);
  and (_25261_, _25260_, _25250_);
  and (_25262_, _08707_, _05422_);
  or (_25263_, _25262_, _25207_);
  and (_25264_, _25263_, _03959_);
  or (_25266_, _25264_, _25261_);
  and (_25267_, _25266_, _04708_);
  or (_25268_, _25207_, _05700_);
  and (_25269_, _25257_, _03866_);
  and (_25270_, _25269_, _25268_);
  or (_25271_, _25270_, _25267_);
  and (_25272_, _25271_, _04706_);
  and (_25273_, _25219_, _03967_);
  and (_25274_, _25273_, _25268_);
  or (_25275_, _25274_, _03835_);
  or (_25277_, _25275_, _25272_);
  nor (_25278_, _12536_, _09899_);
  or (_25279_, _25207_, _06532_);
  or (_25280_, _25279_, _25278_);
  and (_25281_, _25280_, _06537_);
  and (_25282_, _25281_, _25277_);
  nor (_25283_, _08706_, _09899_);
  or (_25284_, _25283_, _25207_);
  and (_25285_, _25284_, _03954_);
  or (_25286_, _25285_, _03703_);
  or (_25288_, _25286_, _25282_);
  or (_25289_, _25216_, _03704_);
  and (_25290_, _25289_, _03702_);
  and (_25291_, _25290_, _25288_);
  and (_25292_, _12596_, _05422_);
  or (_25293_, _25292_, _25207_);
  and (_25294_, _25293_, _03701_);
  or (_25295_, _25294_, _42912_);
  or (_25296_, _25295_, _25291_);
  and (_43260_, _25296_, _25205_);
  or (_25298_, _42908_, \oc8051_golden_model_1.DPH [3]);
  and (_25299_, _25298_, _41654_);
  and (_25300_, _09899_, \oc8051_golden_model_1.DPH [3]);
  nor (_25301_, _12610_, _09899_);
  or (_25302_, _25301_, _25300_);
  or (_25303_, _25302_, _04630_);
  and (_25304_, _05422_, \oc8051_golden_model_1.ACC [3]);
  or (_25305_, _25304_, _25300_);
  and (_25306_, _25305_, _04615_);
  and (_25307_, _04616_, \oc8051_golden_model_1.DPH [3]);
  or (_25309_, _25307_, _03757_);
  or (_25310_, _25309_, _25306_);
  and (_25311_, _25310_, _04537_);
  and (_25312_, _25311_, _25303_);
  nor (_25313_, _09899_, _05050_);
  or (_25314_, _25313_, _25300_);
  and (_25315_, _25314_, _03755_);
  or (_25316_, _25315_, _03750_);
  or (_25317_, _25316_, _25312_);
  or (_25318_, _25305_, _03751_);
  and (_25320_, _25318_, _09822_);
  and (_25321_, _25320_, _25317_);
  or (_25322_, _09922_, \oc8051_golden_model_1.DPH [3]);
  nor (_25323_, _09923_, _09822_);
  and (_25324_, _25323_, _25322_);
  or (_25325_, _25324_, _25321_);
  and (_25326_, _25325_, _09806_);
  nor (_25327_, _09806_, _03669_);
  or (_25328_, _25327_, _07544_);
  or (_25329_, _25328_, _25326_);
  or (_25331_, _25314_, _06994_);
  and (_25332_, _25331_, _25329_);
  or (_25333_, _25332_, _04678_);
  and (_25334_, _06937_, _05422_);
  or (_25335_, _25300_, _04679_);
  or (_25336_, _25335_, _25334_);
  and (_25337_, _25336_, _03415_);
  and (_25338_, _25337_, _25333_);
  nor (_25339_, _12724_, _09899_);
  or (_25340_, _25339_, _25300_);
  and (_25342_, _25340_, _07559_);
  or (_25343_, _25342_, _08854_);
  or (_25344_, _25343_, _25338_);
  and (_25345_, _12738_, _05422_);
  or (_25346_, _25300_, _04703_);
  or (_25347_, _25346_, _25345_);
  and (_25348_, _05422_, _06415_);
  or (_25349_, _25348_, _25300_);
  or (_25350_, _25349_, _04694_);
  and (_25351_, _25350_, _04701_);
  and (_25353_, _25351_, _25347_);
  and (_25354_, _25353_, _25344_);
  and (_25355_, _10455_, _05422_);
  or (_25356_, _25355_, _25300_);
  and (_25357_, _25356_, _03959_);
  or (_25358_, _25357_, _25354_);
  and (_25359_, _25358_, _04708_);
  or (_25360_, _25300_, _05554_);
  and (_25361_, _25349_, _03866_);
  and (_25362_, _25361_, _25360_);
  or (_25364_, _25362_, _25359_);
  and (_25365_, _25364_, _04706_);
  and (_25366_, _25305_, _03967_);
  and (_25367_, _25366_, _25360_);
  or (_25368_, _25367_, _03835_);
  or (_25369_, _25368_, _25365_);
  nor (_25370_, _12737_, _09899_);
  or (_25371_, _25300_, _06532_);
  or (_25372_, _25371_, _25370_);
  and (_25373_, _25372_, _06537_);
  and (_25375_, _25373_, _25369_);
  nor (_25376_, _08701_, _09899_);
  or (_25377_, _25376_, _25300_);
  and (_25378_, _25377_, _03954_);
  or (_25379_, _25378_, _03703_);
  or (_25380_, _25379_, _25375_);
  or (_25381_, _25302_, _03704_);
  and (_25382_, _25381_, _03702_);
  and (_25383_, _25382_, _25380_);
  and (_25384_, _12792_, _05422_);
  or (_25386_, _25384_, _25300_);
  and (_25387_, _25386_, _03701_);
  or (_25388_, _25387_, _42912_);
  or (_25389_, _25388_, _25383_);
  and (_43263_, _25389_, _25299_);
  or (_25390_, _42908_, \oc8051_golden_model_1.DPH [4]);
  and (_25391_, _25390_, _41654_);
  not (_25392_, \oc8051_golden_model_1.DPH [4]);
  nor (_25393_, _05422_, _25392_);
  nor (_25394_, _05898_, _09899_);
  or (_25396_, _25394_, _25393_);
  or (_25397_, _25396_, _06994_);
  nor (_25398_, _12828_, _09899_);
  or (_25399_, _25398_, _25393_);
  or (_25400_, _25399_, _04630_);
  and (_25401_, _05422_, \oc8051_golden_model_1.ACC [4]);
  or (_25402_, _25401_, _25393_);
  and (_25403_, _25402_, _04615_);
  nor (_25404_, _04615_, _25392_);
  or (_25405_, _25404_, _03757_);
  or (_25407_, _25405_, _25403_);
  and (_25408_, _25407_, _04537_);
  and (_25409_, _25408_, _25400_);
  and (_25410_, _25396_, _03755_);
  or (_25411_, _25410_, _03750_);
  or (_25412_, _25411_, _25409_);
  or (_25413_, _25402_, _03751_);
  and (_25414_, _25413_, _09822_);
  and (_25415_, _25414_, _25412_);
  or (_25416_, _09923_, \oc8051_golden_model_1.DPH [4]);
  nor (_25417_, _09924_, _09822_);
  and (_25418_, _25417_, _25416_);
  or (_25419_, _25418_, _25415_);
  and (_25420_, _25419_, _09806_);
  nor (_25421_, _04446_, _09806_);
  or (_25422_, _25421_, _07544_);
  or (_25423_, _25422_, _25420_);
  and (_25424_, _25423_, _25397_);
  or (_25425_, _25424_, _04678_);
  and (_25426_, _06942_, _05422_);
  or (_25429_, _25393_, _04679_);
  or (_25430_, _25429_, _25426_);
  and (_25431_, _25430_, _03415_);
  and (_25432_, _25431_, _25425_);
  nor (_25433_, _12919_, _09899_);
  or (_25434_, _25433_, _25393_);
  and (_25435_, _25434_, _07559_);
  or (_25436_, _25435_, _25432_);
  or (_25437_, _25436_, _08854_);
  and (_25438_, _12933_, _05422_);
  or (_25440_, _25393_, _04703_);
  or (_25441_, _25440_, _25438_);
  and (_25442_, _06422_, _05422_);
  or (_25443_, _25442_, _25393_);
  or (_25444_, _25443_, _04694_);
  and (_25445_, _25444_, _04701_);
  and (_25446_, _25445_, _25441_);
  and (_25447_, _25446_, _25437_);
  and (_25448_, _08700_, _05422_);
  or (_25449_, _25448_, _25393_);
  and (_25451_, _25449_, _03959_);
  or (_25452_, _25451_, _25447_);
  and (_25453_, _25452_, _04708_);
  or (_25454_, _25393_, _08303_);
  and (_25455_, _25443_, _03866_);
  and (_25456_, _25455_, _25454_);
  or (_25457_, _25456_, _25453_);
  and (_25458_, _25457_, _04706_);
  and (_25459_, _25402_, _03967_);
  and (_25460_, _25459_, _25454_);
  or (_25462_, _25460_, _03835_);
  or (_25463_, _25462_, _25458_);
  nor (_25464_, _12931_, _09899_);
  or (_25465_, _25393_, _06532_);
  or (_25466_, _25465_, _25464_);
  and (_25467_, _25466_, _06537_);
  and (_25468_, _25467_, _25463_);
  nor (_25469_, _08699_, _09899_);
  or (_25470_, _25469_, _25393_);
  and (_25471_, _25470_, _03954_);
  or (_25473_, _25471_, _03703_);
  or (_25474_, _25473_, _25468_);
  or (_25475_, _25399_, _03704_);
  and (_25476_, _25475_, _03702_);
  and (_25477_, _25476_, _25474_);
  and (_25478_, _12991_, _05422_);
  or (_25479_, _25478_, _25393_);
  and (_25480_, _25479_, _03701_);
  or (_25481_, _25480_, _42912_);
  or (_25482_, _25481_, _25477_);
  and (_43264_, _25482_, _25391_);
  not (_25484_, \oc8051_golden_model_1.DPH [5]);
  nor (_25485_, _42908_, _25484_);
  nor (_25486_, _05422_, _25484_);
  nor (_25487_, _05799_, _09899_);
  or (_25488_, _25487_, _25486_);
  or (_25489_, _25488_, _06994_);
  nor (_25490_, _13025_, _09899_);
  or (_25491_, _25490_, _25486_);
  or (_25492_, _25491_, _04630_);
  and (_25494_, _05422_, \oc8051_golden_model_1.ACC [5]);
  or (_25495_, _25494_, _25486_);
  and (_25496_, _25495_, _04615_);
  nor (_25497_, _04615_, _25484_);
  or (_25498_, _25497_, _03757_);
  or (_25499_, _25498_, _25496_);
  and (_25500_, _25499_, _04537_);
  and (_25501_, _25500_, _25492_);
  and (_25502_, _25488_, _03755_);
  or (_25503_, _25502_, _03750_);
  or (_25505_, _25503_, _25501_);
  or (_25506_, _25495_, _03751_);
  and (_25507_, _25506_, _09822_);
  and (_25508_, _25507_, _25505_);
  or (_25509_, _09924_, \oc8051_golden_model_1.DPH [5]);
  nor (_25510_, _09925_, _09822_);
  and (_25511_, _25510_, _25509_);
  or (_25512_, _25511_, _25508_);
  and (_25513_, _25512_, _09806_);
  nor (_25514_, _04034_, _09806_);
  or (_25516_, _25514_, _07544_);
  or (_25517_, _25516_, _25513_);
  and (_25518_, _25517_, _25489_);
  or (_25519_, _25518_, _04678_);
  and (_25520_, _06941_, _05422_);
  or (_25521_, _25486_, _04679_);
  or (_25522_, _25521_, _25520_);
  and (_25523_, _25522_, _03415_);
  and (_25524_, _25523_, _25519_);
  nor (_25525_, _13118_, _09899_);
  or (_25527_, _25525_, _25486_);
  and (_25528_, _25527_, _07559_);
  or (_25529_, _25528_, _25524_);
  or (_25530_, _25529_, _08854_);
  and (_25531_, _13133_, _05422_);
  or (_25532_, _25486_, _04703_);
  or (_25533_, _25532_, _25531_);
  and (_25534_, _06371_, _05422_);
  or (_25535_, _25534_, _25486_);
  or (_25536_, _25535_, _04694_);
  and (_25538_, _25536_, _04701_);
  and (_25539_, _25538_, _25533_);
  and (_25540_, _25539_, _25530_);
  and (_25541_, _10451_, _05422_);
  or (_25542_, _25541_, _25486_);
  and (_25543_, _25542_, _03959_);
  or (_25544_, _25543_, _25540_);
  and (_25545_, _25544_, _04708_);
  or (_25546_, _25486_, _08302_);
  and (_25547_, _25535_, _03866_);
  and (_25549_, _25547_, _25546_);
  or (_25550_, _25549_, _25545_);
  and (_25551_, _25550_, _04706_);
  and (_25552_, _25495_, _03967_);
  and (_25553_, _25552_, _25546_);
  or (_25554_, _25553_, _03835_);
  or (_25555_, _25554_, _25551_);
  nor (_25556_, _13131_, _09899_);
  or (_25557_, _25486_, _06532_);
  or (_25558_, _25557_, _25556_);
  and (_25560_, _25558_, _06537_);
  and (_25561_, _25560_, _25555_);
  nor (_25562_, _08697_, _09899_);
  or (_25563_, _25562_, _25486_);
  and (_25564_, _25563_, _03954_);
  or (_25565_, _25564_, _25561_);
  and (_25566_, _25565_, _03704_);
  and (_25567_, _25491_, _03703_);
  or (_25568_, _25567_, _03701_);
  or (_25569_, _25568_, _25566_);
  and (_25571_, _13193_, _05422_);
  or (_25572_, _25486_, _03702_);
  or (_25573_, _25572_, _25571_);
  and (_25574_, _25573_, _42908_);
  and (_25575_, _25574_, _25569_);
  or (_25576_, _25575_, _25485_);
  and (_43265_, _25576_, _41654_);
  or (_25577_, _42908_, \oc8051_golden_model_1.DPH [6]);
  and (_25578_, _25577_, _41654_);
  not (_25579_, \oc8051_golden_model_1.DPH [6]);
  nor (_25581_, _05422_, _25579_);
  nor (_25582_, _06013_, _09899_);
  or (_25583_, _25582_, _25581_);
  or (_25584_, _25583_, _06994_);
  nor (_25585_, _13234_, _09899_);
  or (_25586_, _25585_, _25581_);
  or (_25587_, _25586_, _04630_);
  and (_25588_, _05422_, \oc8051_golden_model_1.ACC [6]);
  or (_25589_, _25588_, _25581_);
  and (_25590_, _25589_, _04615_);
  nor (_25592_, _04615_, _25579_);
  or (_25593_, _25592_, _03757_);
  or (_25594_, _25593_, _25590_);
  and (_25595_, _25594_, _04537_);
  and (_25596_, _25595_, _25587_);
  and (_25597_, _25583_, _03755_);
  or (_25598_, _25597_, _03750_);
  or (_25599_, _25598_, _25596_);
  or (_25600_, _25589_, _03751_);
  and (_25601_, _25600_, _09822_);
  and (_25603_, _25601_, _25599_);
  or (_25604_, _09925_, \oc8051_golden_model_1.DPH [6]);
  and (_25605_, _09926_, _09821_);
  and (_25606_, _25605_, _25604_);
  or (_25607_, _25606_, _25603_);
  and (_25608_, _25607_, _09806_);
  nor (_25609_, _09806_, _03740_);
  or (_25610_, _25609_, _07544_);
  or (_25611_, _25610_, _25608_);
  and (_25612_, _25611_, _25584_);
  or (_25613_, _25612_, _04678_);
  and (_25614_, _06933_, _05422_);
  or (_25615_, _25581_, _04679_);
  or (_25616_, _25615_, _25614_);
  and (_25617_, _25616_, _03415_);
  and (_25618_, _25617_, _25613_);
  nor (_25619_, _13326_, _09899_);
  or (_25620_, _25619_, _25581_);
  and (_25621_, _25620_, _07559_);
  or (_25622_, _25621_, _25618_);
  or (_25625_, _25622_, _08854_);
  and (_25626_, _13341_, _05422_);
  or (_25627_, _25581_, _04703_);
  or (_25628_, _25627_, _25626_);
  and (_25629_, _13333_, _05422_);
  or (_25630_, _25629_, _25581_);
  or (_25631_, _25630_, _04694_);
  and (_25632_, _25631_, _04701_);
  and (_25633_, _25632_, _25628_);
  and (_25634_, _25633_, _25625_);
  and (_25636_, _08695_, _05422_);
  or (_25637_, _25636_, _25581_);
  and (_25638_, _25637_, _03959_);
  or (_25639_, _25638_, _25634_);
  and (_25640_, _25639_, _04708_);
  or (_25641_, _25581_, _08289_);
  and (_25642_, _25630_, _03866_);
  and (_25643_, _25642_, _25641_);
  or (_25644_, _25643_, _25640_);
  and (_25645_, _25644_, _04706_);
  and (_25647_, _25589_, _03967_);
  and (_25648_, _25647_, _25641_);
  or (_25649_, _25648_, _03835_);
  or (_25650_, _25649_, _25645_);
  nor (_25651_, _13340_, _09899_);
  or (_25652_, _25581_, _06532_);
  or (_25653_, _25652_, _25651_);
  and (_25654_, _25653_, _06537_);
  and (_25655_, _25654_, _25650_);
  nor (_25656_, _08694_, _09899_);
  or (_25658_, _25656_, _25581_);
  and (_25659_, _25658_, _03954_);
  or (_25660_, _25659_, _03703_);
  or (_25661_, _25660_, _25655_);
  or (_25662_, _25586_, _03704_);
  and (_25663_, _25662_, _03702_);
  and (_25664_, _25663_, _25661_);
  nor (_25665_, _13399_, _09899_);
  or (_25666_, _25665_, _25581_);
  and (_25667_, _25666_, _03701_);
  or (_25669_, _25667_, _42912_);
  or (_25670_, _25669_, _25664_);
  and (_43266_, _25670_, _25578_);
  nor (_25671_, _03841_, _03399_);
  not (_25672_, _25671_);
  and (_25673_, _25672_, _04326_);
  and (_25674_, _10910_, _10917_);
  nor (_25675_, _25674_, _03129_);
  and (_25676_, _10008_, _10870_);
  nor (_25677_, _25676_, _03129_);
  nor (_25679_, _08399_, _03129_);
  and (_25680_, _08399_, _03129_);
  nor (_25681_, _25680_, _25679_);
  nor (_25682_, _25681_, _10015_);
  not (_25683_, _03481_);
  and (_25684_, _10027_, _06532_);
  nor (_25685_, _25684_, _03129_);
  not (_25686_, _03477_);
  and (_25687_, _10612_, _04708_);
  nor (_25688_, _25687_, _03129_);
  not (_25690_, _03486_);
  and (_25691_, _10585_, _04703_);
  nor (_25692_, _25691_, _03129_);
  and (_25693_, _03839_, _03129_);
  nor (_25694_, _03861_, _07559_);
  and (_25695_, _25694_, _10517_);
  nor (_25696_, _25695_, _03129_);
  nor (_25697_, _04326_, _03442_);
  and (_25698_, _10423_, _03129_);
  and (_25699_, _04326_, \oc8051_golden_model_1.PC [0]);
  nor (_25701_, _25699_, _10253_);
  not (_25702_, _25701_);
  nor (_25703_, _25702_, _10423_);
  nor (_25704_, _25703_, _25698_);
  nor (_25705_, _25704_, _10388_);
  nor (_25706_, _04326_, _03448_);
  nor (_25707_, _10344_, _03129_);
  and (_25708_, _04944_, _04235_);
  nor (_25709_, _25708_, _03129_);
  and (_25710_, _25708_, _03129_);
  nor (_25712_, _25710_, _25709_);
  and (_25713_, _25712_, _04948_);
  not (_25714_, _25713_);
  not (_25715_, _10344_);
  nor (_25716_, _04326_, _04948_);
  nor (_25717_, _25716_, _25715_);
  and (_25718_, _25717_, _25714_);
  nor (_25719_, _25718_, _25707_);
  nor (_25720_, _25719_, _10320_);
  and (_25721_, _10326_, \oc8051_golden_model_1.PC [0]);
  not (_25723_, _25721_);
  and (_25724_, _04211_, _03129_);
  nor (_25725_, _25724_, _10092_);
  and (_25726_, _25725_, _10324_);
  nor (_25727_, _25726_, _06140_);
  and (_25728_, _25727_, _25723_);
  or (_25729_, _25728_, _25720_);
  nor (_25730_, _25729_, _04624_);
  and (_25731_, _04624_, _03129_);
  nor (_25732_, _25731_, _25730_);
  nor (_25734_, _25732_, _03757_);
  and (_25735_, _25701_, _10316_);
  and (_25736_, _10314_, _03129_);
  nor (_25737_, _25736_, _25735_);
  nor (_25738_, _25737_, _04630_);
  nor (_25739_, _25738_, _10355_);
  not (_25740_, _25739_);
  nor (_25741_, _25740_, _25734_);
  nor (_25742_, _10354_, _03129_);
  nor (_25743_, _25742_, _04933_);
  not (_25745_, _25743_);
  nor (_25746_, _25745_, _25741_);
  nor (_25747_, _04326_, _03445_);
  and (_25748_, _10375_, _10364_);
  not (_25749_, _25748_);
  nor (_25750_, _25749_, _25747_);
  not (_25751_, _25750_);
  nor (_25752_, _25751_, _25746_);
  nor (_25753_, _25748_, _03129_);
  nor (_25754_, _25753_, _10379_);
  not (_25756_, _25754_);
  nor (_25757_, _25756_, _25752_);
  nor (_25758_, _25757_, _25706_);
  nor (_25759_, _25758_, _10425_);
  nor (_25760_, _25759_, _25705_);
  nor (_25761_, _25760_, _03854_);
  nand (_25762_, _10181_, \oc8051_golden_model_1.PC [0]);
  or (_25763_, _25701_, _10181_);
  and (_25764_, _25763_, _03854_);
  and (_25765_, _25764_, _25762_);
  or (_25767_, _25765_, _25761_);
  and (_25768_, _25767_, _04216_);
  and (_25769_, _10462_, _03129_);
  nor (_25770_, _25702_, _10462_);
  nor (_25771_, _25770_, _25769_);
  nor (_25772_, _25771_, _04216_);
  nor (_25773_, _25772_, _25768_);
  nor (_25774_, _25773_, _03847_);
  and (_25775_, _10446_, \oc8051_golden_model_1.PC [0]);
  nor (_25776_, _25701_, _10446_);
  or (_25778_, _25776_, _11721_);
  nor (_25779_, _25778_, _25775_);
  or (_25780_, _25779_, _25774_);
  and (_25781_, _25780_, _10432_);
  and (_25782_, _10431_, _03129_);
  or (_25783_, _25782_, _25781_);
  and (_25784_, _25783_, _03442_);
  or (_25785_, _25784_, _10481_);
  nor (_25786_, _25785_, _25697_);
  not (_25787_, _03453_);
  nor (_25789_, _10477_, _03129_);
  nor (_25790_, _25789_, _25787_);
  not (_25791_, _25790_);
  nor (_25792_, _25791_, _25786_);
  nor (_25793_, _04326_, _03453_);
  and (_25794_, _10488_, _03422_);
  not (_25795_, _25794_);
  nor (_25796_, _25795_, _25793_);
  not (_25797_, _25796_);
  nor (_25798_, _25797_, _25792_);
  nor (_25800_, _25794_, _03129_);
  nor (_25801_, _25800_, _03676_);
  not (_25802_, _25801_);
  nor (_25803_, _25802_, _25798_);
  nor (_25804_, _04326_, _03418_);
  not (_25805_, _25695_);
  nor (_25806_, _25805_, _25804_);
  not (_25807_, _25806_);
  nor (_25808_, _25807_, _25803_);
  or (_25809_, _25808_, _03487_);
  nor (_25811_, _25809_, _25696_);
  nor (_25812_, _10525_, _03487_);
  not (_25813_, _25812_);
  nand (_25814_, _10526_, _04326_);
  and (_25815_, _25814_, _25813_);
  nor (_25816_, _25815_, _25811_);
  nor (_25817_, _25725_, _10526_);
  nor (_25818_, _25817_, _25816_);
  and (_25819_, _25818_, _04694_);
  or (_25820_, _25819_, _25693_);
  and (_25822_, _25820_, _10541_);
  and (_25823_, _10540_, _03549_);
  or (_25824_, _25823_, _25822_);
  and (_25825_, _25824_, _11594_);
  nor (_25826_, _04326_, _11594_);
  or (_25827_, _25826_, _25825_);
  and (_25828_, _25827_, _10580_);
  not (_25829_, _25691_);
  and (_25830_, _08783_, \oc8051_golden_model_1.PC [0]);
  and (_25831_, _25725_, _10146_);
  or (_25833_, _25831_, _25830_);
  and (_25834_, _25833_, _10145_);
  nor (_25835_, _25834_, _25829_);
  not (_25836_, _25835_);
  nor (_25837_, _25836_, _25828_);
  nor (_25838_, _25837_, _25692_);
  and (_25839_, _25838_, _25690_);
  nor (_25840_, _04326_, _25690_);
  or (_25841_, _25840_, _25839_);
  and (_25842_, _25841_, _10602_);
  not (_25844_, _25687_);
  nor (_25845_, _25725_, _10146_);
  nor (_25846_, _08783_, \oc8051_golden_model_1.PC [0]);
  nor (_25847_, _25846_, _10602_);
  not (_25848_, _25847_);
  nor (_25849_, _25848_, _25845_);
  nor (_25850_, _25849_, _25844_);
  not (_25851_, _25850_);
  nor (_25852_, _25851_, _25842_);
  nor (_25853_, _25852_, _25688_);
  and (_25855_, _25853_, _25686_);
  nor (_25856_, _04326_, _25686_);
  or (_25857_, _25856_, _25855_);
  and (_25858_, _25857_, _10030_);
  not (_25859_, _25684_);
  nor (_25860_, _25725_, \oc8051_golden_model_1.PSW [7]);
  and (_25861_, \oc8051_golden_model_1.PSW [7], _03129_);
  nor (_25862_, _25861_, _10030_);
  not (_25863_, _25862_);
  nor (_25864_, _25863_, _25860_);
  nor (_25866_, _25864_, _25859_);
  not (_25867_, _25866_);
  nor (_25868_, _25867_, _25858_);
  nor (_25869_, _25868_, _25685_);
  and (_25870_, _25869_, _25683_);
  nor (_25871_, _04326_, _25683_);
  or (_25872_, _25871_, _25870_);
  and (_25873_, _25872_, _10015_);
  and (_25874_, _10012_, _08007_);
  not (_25875_, _25874_);
  or (_25877_, _25875_, _25873_);
  nor (_25878_, _25877_, _25682_);
  nor (_25879_, _25874_, _03129_);
  nor (_25880_, _25879_, _03974_);
  not (_25881_, _25880_);
  nor (_25882_, _25881_, _25878_);
  and (_25883_, _06935_, _03974_);
  or (_25884_, _25883_, _25882_);
  and (_25885_, _25884_, _06543_);
  nor (_25886_, _04326_, _06543_);
  or (_25888_, _25886_, _25885_);
  and (_25889_, _25888_, _04386_);
  and (_25890_, _25702_, _10860_);
  nor (_25891_, _10860_, _03129_);
  or (_25892_, _25891_, _04386_);
  or (_25893_, _25892_, _25890_);
  and (_25894_, _25893_, _25676_);
  not (_25895_, _25894_);
  nor (_25896_, _25895_, _25889_);
  nor (_25897_, _25896_, _25677_);
  and (_25899_, _25897_, _03708_);
  and (_25900_, _06935_, _03707_);
  or (_25901_, _25900_, _25899_);
  and (_25902_, _25901_, _03395_);
  nor (_25903_, _04326_, _03395_);
  nor (_25904_, _25903_, _25902_);
  nor (_25905_, _25904_, _03705_);
  and (_25906_, _10860_, \oc8051_golden_model_1.PC [0]);
  nor (_25907_, _25701_, _10860_);
  nor (_25908_, _25907_, _25906_);
  and (_25910_, _25908_, _03705_);
  or (_25911_, _25910_, _25905_);
  and (_25912_, _10887_, _10894_);
  and (_25913_, _25912_, _25911_);
  nor (_25914_, _25912_, \oc8051_golden_model_1.PC [0]);
  or (_25915_, _25914_, _05156_);
  nor (_25916_, _25915_, _25913_);
  and (_25917_, _05156_, _04326_);
  nor (_25918_, _25917_, _03384_);
  not (_25919_, _25918_);
  nor (_25921_, _25919_, _25916_);
  not (_25922_, _25674_);
  and (_25923_, _25908_, _03384_);
  nor (_25924_, _25923_, _25922_);
  not (_25925_, _25924_);
  nor (_25926_, _25925_, _25921_);
  nor (_25927_, _25926_, _25675_);
  nor (_25928_, _25927_, _25672_);
  or (_25929_, _25928_, _10928_);
  nor (_25930_, _25929_, _25673_);
  and (_25932_, _10928_, _03129_);
  nor (_25933_, _25932_, _25930_);
  nand (_25934_, _25933_, _42908_);
  or (_25935_, _42908_, \oc8051_golden_model_1.PC [0]);
  and (_25936_, _25935_, _41654_);
  and (_43269_, _25936_, _25934_);
  nor (_25937_, _10917_, _10251_);
  and (_25938_, _12195_, _10251_);
  nor (_25939_, _04947_, _10251_);
  or (_25940_, _06992_, _04079_);
  and (_25942_, _10860_, _10251_);
  nor (_25943_, _10255_, _10253_);
  nor (_25944_, _25943_, _10256_);
  nor (_25945_, _25944_, _10860_);
  nor (_25946_, _25945_, _25942_);
  and (_25947_, _25946_, _03384_);
  and (_25948_, _03703_, _03100_);
  nor (_25949_, _13156_, _10251_);
  nor (_25950_, _08643_, _10251_);
  nor (_25951_, _10012_, _10251_);
  nor (_25953_, _10027_, _10251_);
  nor (_25954_, _10614_, _03100_);
  and (_25955_, _04671_, _03476_);
  and (_25956_, _25955_, _03492_);
  nor (_25957_, _10585_, _10251_);
  nor (_25958_, _06305_, _03100_);
  and (_25959_, _03679_, \oc8051_golden_model_1.PC [1]);
  nor (_25960_, _10488_, _10251_);
  and (_25961_, _10181_, _03492_);
  not (_25962_, _25961_);
  not (_25963_, _25944_);
  nor (_25964_, _25963_, _10181_);
  nor (_25965_, _25964_, _03855_);
  and (_25966_, _25965_, _25962_);
  and (_25967_, _06241_, _05553_);
  and (_25968_, _05699_, _05602_);
  and (_25969_, _25968_, _05652_);
  and (_25970_, _25969_, _06016_);
  nand (_25971_, _25970_, _25967_);
  or (_25972_, _25971_, _10251_);
  and (_25975_, _25944_, _10316_);
  nor (_25976_, _25975_, _04630_);
  and (_25977_, _25976_, _25972_);
  or (_25978_, _10324_, \oc8051_golden_model_1.PC [1]);
  nor (_25979_, _10094_, _10092_);
  nor (_25980_, _25979_, _10095_);
  nand (_25981_, _25980_, _10324_);
  and (_25982_, _25981_, _10320_);
  and (_25983_, _25982_, _25978_);
  nor (_25984_, _10344_, _10251_);
  nor (_25986_, _04615_, \oc8051_golden_model_1.PC [0]);
  and (_25987_, _04944_, _10331_);
  nor (_25988_, _25987_, _25986_);
  and (_25989_, _25988_, \oc8051_golden_model_1.PC [1]);
  nor (_25990_, _25988_, \oc8051_golden_model_1.PC [1]);
  nor (_25991_, _25990_, _25989_);
  and (_25992_, _25991_, _04948_);
  not (_25993_, _25992_);
  nor (_25994_, _04515_, _04948_);
  nor (_25995_, _25994_, _25715_);
  and (_25997_, _25995_, _25993_);
  nor (_25998_, _25997_, _25984_);
  nor (_25999_, _25998_, _10320_);
  or (_26000_, _25999_, _25983_);
  or (_26001_, _26000_, _04624_);
  nand (_26002_, _04624_, _10251_);
  and (_26003_, _26002_, _04630_);
  and (_26004_, _26003_, _26001_);
  or (_26005_, _26004_, _25977_);
  nand (_26006_, _26005_, _10354_);
  nor (_26008_, _10354_, _10251_);
  nor (_26009_, _26008_, _03696_);
  nand (_26010_, _26009_, _26006_);
  and (_26011_, _03696_, _03100_);
  nor (_26012_, _26011_, _04933_);
  nand (_26013_, _26012_, _26010_);
  and (_26014_, _04515_, _04933_);
  nor (_26015_, _26014_, _03755_);
  nand (_26016_, _26015_, _26013_);
  and (_26017_, _03755_, _03100_);
  nor (_26019_, _26017_, _10365_);
  nand (_26020_, _26019_, _26016_);
  nor (_26021_, _10364_, _10251_);
  nor (_26022_, _26021_, _03750_);
  nand (_26023_, _26022_, _26020_);
  and (_26024_, _03750_, _03100_);
  nor (_26025_, _26024_, _10377_);
  nand (_26026_, _26025_, _26023_);
  nor (_26027_, _10375_, _10251_);
  nor (_26028_, _26027_, _03691_);
  nand (_26030_, _26028_, _26026_);
  and (_26031_, _03691_, _03100_);
  nor (_26032_, _26031_, _10379_);
  nand (_26033_, _26032_, _26030_);
  and (_26034_, _04515_, _10379_);
  nor (_26035_, _26034_, _03690_);
  nand (_26036_, _26035_, _26033_);
  and (_26037_, _03690_, _03100_);
  nor (_26038_, _26037_, _10387_);
  nand (_26039_, _26038_, _26036_);
  not (_26041_, _10386_);
  nor (_26042_, _25944_, _10423_);
  and (_26043_, _10423_, _10251_);
  nor (_26044_, _26043_, _26042_);
  and (_26045_, _26044_, _26041_);
  or (_26046_, _26045_, _10388_);
  nand (_26047_, _26046_, _26039_);
  and (_26048_, _26044_, _10386_);
  nor (_26049_, _26048_, _03854_);
  and (_26050_, _26049_, _26047_);
  nor (_26052_, _26050_, _25966_);
  nand (_26053_, _26052_, _10433_);
  nor (_26054_, _25963_, _10446_);
  and (_26055_, _10446_, _03492_);
  nor (_26056_, _26055_, _26054_);
  nor (_26057_, _26056_, _11721_);
  and (_26058_, _10462_, _03492_);
  nor (_26059_, _25963_, _10462_);
  nor (_26060_, _26059_, _26058_);
  nor (_26061_, _26060_, _04216_);
  nor (_26063_, _26061_, _26057_);
  and (_26064_, _10431_, _10251_);
  nor (_26065_, _26064_, _03684_);
  and (_26066_, _26065_, _26063_);
  nand (_26067_, _26066_, _26053_);
  and (_26068_, _03684_, \oc8051_golden_model_1.PC [1]);
  nor (_26069_, _26068_, _05105_);
  nand (_26070_, _26069_, _26067_);
  nor (_26071_, _04515_, _03442_);
  and (_26072_, _03802_, _03795_);
  nor (_26073_, _03804_, _03777_);
  and (_26074_, _26073_, _04663_);
  and (_26075_, _26074_, _26072_);
  not (_26076_, _26075_);
  nor (_26077_, _26076_, _26071_);
  nand (_26078_, _26077_, _26070_);
  nor (_26079_, _26075_, _03100_);
  nor (_26080_, _26079_, _10474_);
  nand (_26081_, _26080_, _26078_);
  and (_26082_, _10476_, _03492_);
  or (_26085_, _26082_, _10477_);
  nand (_26086_, _26085_, _26081_);
  nor (_26087_, _10476_, _10251_);
  nor (_26088_, _26087_, _03811_);
  nand (_26089_, _26088_, _26086_);
  and (_26090_, _03811_, _03100_);
  nor (_26091_, _26090_, _25787_);
  nand (_26092_, _26091_, _26089_);
  and (_26093_, _04515_, _25787_);
  nor (_26094_, _26093_, _03810_);
  nand (_26096_, _26094_, _26092_);
  and (_26097_, _03810_, _03100_);
  nor (_26098_, _26097_, _10494_);
  and (_26099_, _26098_, _26096_);
  or (_26100_, _26099_, _25960_);
  nand (_26101_, _26100_, _10492_);
  nor (_26102_, _10492_, _03100_);
  nor (_26103_, _26102_, _03547_);
  nand (_26104_, _26103_, _26101_);
  nor (_26105_, _03492_, _03422_);
  nor (_26107_, _26105_, _03679_);
  and (_26108_, _26107_, _26104_);
  or (_26109_, _26108_, _25959_);
  nand (_26110_, _26109_, _03418_);
  and (_26111_, _04515_, _03676_);
  nor (_26112_, _26111_, _03861_);
  nand (_26113_, _26112_, _26110_);
  and (_26114_, _03861_, _03492_);
  nor (_26115_, _26114_, _11528_);
  nand (_26116_, _26115_, _26113_);
  nor (_26118_, _10510_, _03100_);
  nor (_26119_, _26118_, _07559_);
  nand (_26120_, _26119_, _26116_);
  nor (_26121_, _10251_, _03415_);
  nor (_26122_, _26121_, _10521_);
  nand (_26123_, _26122_, _26120_);
  nor (_26124_, _10517_, _10251_);
  nor (_26125_, _26124_, _03746_);
  nand (_26126_, _26125_, _26123_);
  and (_26127_, _03746_, _03100_);
  nor (_26129_, _26127_, _03487_);
  nand (_26130_, _26129_, _26126_);
  and (_26131_, _04515_, _03487_);
  nor (_26132_, _26131_, _10525_);
  nand (_26133_, _26132_, _26130_);
  and (_26134_, _25980_, _10525_);
  nor (_26135_, _26134_, _06306_);
  and (_26136_, _26135_, _26133_);
  or (_26137_, _26136_, _25958_);
  nand (_26138_, _26137_, _04694_);
  and (_26140_, _03839_, _10251_);
  nor (_26141_, _26140_, _08456_);
  nand (_26142_, _26141_, _26138_);
  and (_26143_, _08456_, _03100_);
  nor (_26144_, _26143_, _10540_);
  nand (_26145_, _26144_, _26142_);
  nor (_26146_, _10541_, _03568_);
  nor (_26147_, _26146_, _03745_);
  and (_26148_, _26147_, _26145_);
  and (_26149_, _03745_, _03100_);
  or (_26151_, _26149_, _03483_);
  or (_26152_, _26151_, _26148_);
  and (_26153_, _04515_, _03483_);
  nor (_26154_, _26153_, _10145_);
  nand (_26155_, _26154_, _26152_);
  nor (_26156_, _25980_, _08783_);
  and (_26157_, _08783_, \oc8051_golden_model_1.PC [1]);
  nor (_26158_, _26157_, _10580_);
  not (_26159_, _26158_);
  nor (_26160_, _26159_, _26156_);
  nor (_26162_, _26160_, _10587_);
  and (_26163_, _26162_, _26155_);
  or (_26164_, _26163_, _25957_);
  nand (_26165_, _26164_, _10589_);
  nor (_26166_, _10589_, _03100_);
  nor (_26167_, _26166_, _03838_);
  and (_26168_, _26167_, _26165_);
  and (_26169_, _03838_, _03492_);
  or (_26170_, _26169_, _03959_);
  nor (_26171_, _26170_, _26168_);
  and (_26173_, _03959_, \oc8051_golden_model_1.PC [1]);
  or (_26174_, _26173_, _26171_);
  nand (_26175_, _26174_, _25690_);
  and (_26176_, _04515_, _03486_);
  nor (_26177_, _26176_, _10601_);
  nand (_26178_, _26177_, _26175_);
  nor (_26179_, _25980_, _10146_);
  nor (_26180_, _08783_, _03100_);
  nor (_26181_, _26180_, _10602_);
  not (_26182_, _26181_);
  nor (_26184_, _26182_, _26179_);
  nor (_26185_, _26184_, _25955_);
  and (_26186_, _26185_, _26178_);
  nor (_26187_, _26186_, _25956_);
  nor (_26188_, _04220_, _03789_);
  nor (_26189_, _04957_, _12353_);
  and (_26190_, _26189_, _26188_);
  nor (_26191_, _26190_, _04346_);
  or (_26192_, _26191_, _26187_);
  and (_26193_, _04223_, _03476_);
  and (_26195_, _26191_, _03492_);
  nor (_26196_, _26195_, _26193_);
  nand (_26197_, _26196_, _26192_);
  and (_26198_, _26193_, _10251_);
  nor (_26199_, _26198_, _10615_);
  and (_26200_, _26199_, _26197_);
  or (_26201_, _26200_, _25954_);
  nand (_26202_, _26201_, _04708_);
  and (_26203_, _03866_, _10251_);
  nor (_26204_, _26203_, _03967_);
  nand (_26206_, _26204_, _26202_);
  and (_26207_, _03967_, _03100_);
  nor (_26208_, _26207_, _03477_);
  nand (_26209_, _26208_, _26206_);
  and (_26210_, _04515_, _03477_);
  nor (_26211_, _26210_, _10029_);
  nand (_26212_, _26211_, _26209_);
  nor (_26213_, _25980_, \oc8051_golden_model_1.PSW [7]);
  and (_26214_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor (_26215_, _26214_, _10030_);
  not (_26217_, _26215_);
  nor (_26218_, _26217_, _26213_);
  nor (_26219_, _26218_, _10628_);
  and (_26220_, _26219_, _26212_);
  or (_26221_, _26220_, _25953_);
  nand (_26222_, _26221_, _08527_);
  nor (_26223_, _08527_, _03100_);
  nor (_26224_, _26223_, _03835_);
  and (_26225_, _26224_, _26222_);
  and (_26226_, _03835_, _03492_);
  or (_26228_, _26226_, _03954_);
  nor (_26229_, _26228_, _26225_);
  and (_26230_, _03954_, \oc8051_golden_model_1.PC [1]);
  or (_26231_, _26230_, _26229_);
  nand (_26232_, _26231_, _25683_);
  and (_26233_, _04515_, _03481_);
  nor (_26234_, _26233_, _10014_);
  nand (_26235_, _26234_, _26232_);
  nor (_26236_, _25980_, _08059_);
  and (_26237_, _08059_, \oc8051_golden_model_1.PC [1]);
  nor (_26239_, _26237_, _10015_);
  not (_26240_, _26239_);
  nor (_26241_, _26240_, _26236_);
  nor (_26242_, _26241_, _10646_);
  and (_26243_, _26242_, _26235_);
  or (_26244_, _26243_, _25951_);
  nand (_26245_, _26244_, _10010_);
  nor (_26246_, _10010_, _03100_);
  nor (_26247_, _26246_, _08006_);
  nand (_26248_, _26247_, _26245_);
  and (_26250_, _08006_, _10251_);
  nor (_26251_, _26250_, _03974_);
  and (_26252_, _26251_, _26248_);
  and (_26253_, _06653_, _03974_);
  or (_26254_, _26253_, _26252_);
  nand (_26255_, _26254_, _06543_);
  and (_26256_, _04515_, _03474_);
  nor (_26257_, _26256_, _03831_);
  nand (_26258_, _26257_, _26255_);
  not (_26259_, _08643_);
  and (_26261_, _25963_, _10860_);
  nor (_26262_, _10860_, _03492_);
  or (_26263_, _26262_, _04386_);
  nor (_26264_, _26263_, _26261_);
  nor (_26265_, _26264_, _26259_);
  and (_26266_, _26265_, _26258_);
  or (_26267_, _26266_, _25950_);
  and (_26268_, _12353_, _03393_);
  nor (_26269_, _10005_, _26268_);
  nand (_26270_, _26269_, _26267_);
  and (_26272_, _04223_, _03393_);
  nor (_26273_, _26269_, _10251_);
  nor (_26274_, _26273_, _26272_);
  nand (_26275_, _26274_, _26270_);
  and (_26276_, _26272_, _10251_);
  nor (_26277_, _26276_, _09990_);
  nand (_26278_, _26277_, _26275_);
  nor (_26279_, _09989_, _03100_);
  nor (_26280_, _26279_, _07964_);
  and (_26281_, _26280_, _26278_);
  and (_26283_, _07964_, _10251_);
  or (_26284_, _26283_, _03707_);
  or (_26285_, _26284_, _26281_);
  and (_26286_, _06653_, _03707_);
  nor (_26287_, _26286_, _03394_);
  and (_26288_, _26287_, _26285_);
  nor (_26289_, _04515_, _03395_);
  or (_26290_, _26289_, _26288_);
  nand (_26291_, _26290_, _03706_);
  not (_26292_, _13156_);
  and (_26294_, _25946_, _03705_);
  nor (_26295_, _26294_, _26292_);
  and (_26296_, _26295_, _26291_);
  or (_26297_, _26296_, _25949_);
  nor (_26298_, _04727_, _13157_);
  nand (_26299_, _26298_, _26297_);
  nor (_26300_, _26298_, _10251_);
  nor (_26301_, _26300_, _03703_);
  and (_26302_, _26301_, _26299_);
  or (_26303_, _26302_, _25948_);
  nand (_26305_, _26303_, _10894_);
  nor (_26306_, _10894_, _03492_);
  nor (_26307_, _26306_, _05156_);
  nand (_26308_, _26307_, _26305_);
  and (_26309_, _05156_, _04515_);
  nor (_26310_, _26309_, _03384_);
  and (_26311_, _26310_, _26308_);
  or (_26312_, _26311_, _25947_);
  nand (_26313_, _26312_, _25940_);
  nor (_26314_, _25940_, _03492_);
  nor (_26316_, _12384_, _04905_);
  not (_26317_, _26316_);
  nor (_26318_, _26317_, _26314_);
  and (_26319_, _26318_, _26313_);
  nor (_26320_, _26319_, _25939_);
  nor (_26321_, _26320_, _25938_);
  or (_26322_, _26321_, _03701_);
  not (_26323_, _10917_);
  and (_26324_, _03701_, _03100_);
  nor (_26325_, _26324_, _26323_);
  and (_26327_, _26325_, _26322_);
  or (_26328_, _26327_, _25937_);
  nand (_26329_, _26328_, _25671_);
  and (_26330_, _25672_, _04515_);
  nor (_26331_, _26330_, _10928_);
  and (_26332_, _26331_, _26329_);
  and (_26333_, _10928_, _10251_);
  or (_26334_, _26333_, _26332_);
  or (_26335_, _26334_, _42912_);
  or (_26336_, _42908_, \oc8051_golden_model_1.PC [1]);
  and (_26338_, _26336_, _41654_);
  and (_43270_, _26338_, _26335_);
  and (_26339_, _10928_, _03461_);
  and (_26340_, _03701_, _03405_);
  and (_26341_, _03703_, _03405_);
  nor (_26342_, _10008_, _03461_);
  nor (_26343_, _10012_, _03461_);
  nor (_26344_, _10027_, _03461_);
  nor (_26345_, _10612_, _03461_);
  nor (_26346_, _10585_, _03461_);
  and (_26348_, _10248_, _03861_);
  not (_26349_, _26348_);
  and (_26350_, _03810_, _03405_);
  and (_26351_, _10431_, _03462_);
  and (_26352_, _04624_, _03462_);
  nor (_26353_, _10344_, _03461_);
  nand (_26354_, _04109_, _10089_);
  and (_26355_, _04944_, \oc8051_golden_model_1.PC [2]);
  or (_26356_, _26355_, _04615_);
  and (_26357_, _26356_, _04235_);
  nor (_26359_, _04944_, _03462_);
  or (_26360_, _26359_, _26357_);
  and (_26361_, _26360_, _26354_);
  and (_26362_, _04234_, _03461_);
  nor (_26363_, _26362_, _26361_);
  nor (_26364_, _26363_, _04111_);
  not (_26365_, _26364_);
  nor (_26366_, _04948_, _04077_);
  nor (_26367_, _26366_, _25715_);
  and (_26368_, _26367_, _26365_);
  nor (_26370_, _26368_, _26353_);
  nor (_26371_, _26370_, _10320_);
  or (_26372_, _10324_, _10089_);
  and (_26373_, _10099_, _10096_);
  nor (_26374_, _26373_, _10100_);
  nand (_26375_, _26374_, _10324_);
  and (_26376_, _26375_, _10320_);
  and (_26377_, _26376_, _26372_);
  or (_26378_, _26377_, _26371_);
  and (_26379_, _26378_, _04625_);
  nor (_26381_, _26379_, _26352_);
  and (_26382_, _26381_, _04630_);
  and (_26383_, _06241_, _05699_);
  and (_26384_, _26383_, _05553_);
  and (_26385_, _06016_, _05652_);
  and (_26386_, _26385_, _05602_);
  and (_26387_, _26386_, _26384_);
  and (_26388_, _10260_, _10257_);
  nor (_26389_, _26388_, _10261_);
  or (_26390_, _26389_, _26387_);
  nand (_26392_, _26387_, _10249_);
  and (_26393_, _26392_, _03757_);
  and (_26394_, _26393_, _26390_);
  or (_26395_, _26394_, _10355_);
  or (_26396_, _26395_, _26382_);
  nor (_26397_, _10354_, _03461_);
  nor (_26398_, _26397_, _03696_);
  nand (_26399_, _26398_, _26396_);
  and (_26400_, _03696_, _03405_);
  nor (_26401_, _26400_, _04933_);
  nand (_26403_, _26401_, _26399_);
  and (_26404_, _04077_, _04933_);
  nor (_26405_, _26404_, _03755_);
  nand (_26406_, _26405_, _26403_);
  and (_26407_, _03755_, _03405_);
  nor (_26408_, _26407_, _10365_);
  nand (_26409_, _26408_, _26406_);
  nor (_26410_, _10364_, _03461_);
  nor (_26411_, _26410_, _03750_);
  nand (_26412_, _26411_, _26409_);
  and (_26414_, _03750_, _03405_);
  nor (_26415_, _26414_, _10377_);
  nand (_26416_, _26415_, _26412_);
  nor (_26417_, _10375_, _03461_);
  nor (_26418_, _26417_, _03691_);
  nand (_26419_, _26418_, _26416_);
  and (_26420_, _03691_, _03405_);
  nor (_26421_, _26420_, _10379_);
  nand (_26422_, _26421_, _26419_);
  and (_26423_, _04077_, _10379_);
  nor (_26425_, _26423_, _03690_);
  nand (_26426_, _26425_, _26422_);
  and (_26427_, _03690_, _03405_);
  nor (_26428_, _26427_, _10425_);
  and (_26429_, _26428_, _26426_);
  nor (_26430_, _26389_, _10423_);
  and (_26431_, _10423_, _10249_);
  nor (_26432_, _26431_, _26430_);
  nor (_26433_, _26432_, _10388_);
  or (_26434_, _26433_, _26429_);
  nand (_26436_, _26434_, _03855_);
  not (_26437_, _26389_);
  nor (_26438_, _26437_, _10181_);
  nand (_26439_, _10248_, _10181_);
  nand (_26440_, _26439_, _03854_);
  or (_26441_, _26440_, _26438_);
  and (_26442_, _26441_, _04216_);
  nand (_26443_, _26442_, _26436_);
  and (_26444_, _10462_, _10249_);
  nor (_26445_, _26389_, _10462_);
  or (_26447_, _26445_, _04216_);
  or (_26448_, _26447_, _26444_);
  nand (_26449_, _26448_, _26443_);
  nand (_26450_, _26449_, _11721_);
  and (_26451_, _10446_, _10249_);
  nor (_26452_, _26389_, _10446_);
  or (_26453_, _26452_, _11721_);
  nor (_26454_, _26453_, _26451_);
  nor (_26455_, _26454_, _10431_);
  and (_26456_, _26455_, _26450_);
  or (_26458_, _26456_, _26351_);
  nand (_26459_, _26458_, _03685_);
  and (_26460_, _03684_, _10089_);
  nor (_26461_, _26460_, _05105_);
  nand (_26462_, _26461_, _26459_);
  nor (_26463_, _04077_, _03442_);
  nor (_26464_, _26463_, _26076_);
  and (_26465_, _26464_, _26462_);
  nor (_26466_, _26075_, _03405_);
  or (_26467_, _26466_, _26465_);
  nand (_26469_, _26467_, _10477_);
  nor (_26470_, _10477_, _03461_);
  nor (_26471_, _26470_, _03811_);
  nand (_26472_, _26471_, _26469_);
  and (_26473_, _03811_, _03405_);
  nor (_26474_, _26473_, _25787_);
  nand (_26475_, _26474_, _26472_);
  and (_26476_, _04077_, _25787_);
  nor (_26477_, _26476_, _03810_);
  nand (_26478_, _26477_, _26475_);
  nand (_26480_, _26478_, _10488_);
  nor (_26481_, _26480_, _26350_);
  nor (_26482_, _10488_, _03461_);
  or (_26483_, _26482_, _26481_);
  nand (_26484_, _26483_, _10492_);
  nor (_26485_, _10492_, _03405_);
  nor (_26486_, _26485_, _03547_);
  and (_26487_, _26486_, _26484_);
  nor (_26488_, _03462_, _03422_);
  or (_26489_, _26488_, _03679_);
  nor (_26491_, _26489_, _26487_);
  and (_26492_, _03679_, _10089_);
  or (_26493_, _26492_, _26491_);
  nand (_26494_, _26493_, _03418_);
  and (_26495_, _04077_, _03676_);
  nor (_26496_, _26495_, _03861_);
  nand (_26497_, _26496_, _26494_);
  and (_26498_, _26497_, _26349_);
  or (_26499_, _26498_, _06993_);
  nor (_26500_, _04678_, _04287_);
  nand (_26502_, _06993_, _03405_);
  and (_26503_, _26502_, _26500_);
  nand (_26504_, _26503_, _26499_);
  nor (_26505_, _26500_, _03405_);
  nor (_26506_, _26505_, _07559_);
  nand (_26507_, _26506_, _26504_);
  nor (_26508_, _10249_, _03415_);
  nor (_26509_, _26508_, _10521_);
  nand (_26510_, _26509_, _26507_);
  nor (_26511_, _10517_, _03461_);
  nor (_26513_, _26511_, _03746_);
  and (_26514_, _26513_, _26510_);
  and (_26515_, _03746_, _03405_);
  or (_26516_, _26515_, _03487_);
  nor (_26517_, _26516_, _26514_);
  and (_26518_, _04077_, _03487_);
  or (_26519_, _26518_, _26517_);
  nand (_26520_, _26519_, _10526_);
  nor (_26521_, _26374_, _10526_);
  and (_26522_, _03786_, _03482_);
  not (_26523_, _26522_);
  and (_26524_, _06301_, _26523_);
  and (_26525_, _26524_, _06302_);
  not (_26526_, _26525_);
  nor (_26527_, _26526_, _26521_);
  nand (_26528_, _26527_, _26520_);
  nor (_26529_, _26525_, _10089_);
  and (_26530_, _03789_, _03482_);
  or (_26531_, _04689_, _26530_);
  nor (_26532_, _26531_, _26529_);
  nand (_26535_, _26532_, _26528_);
  nand (_26536_, _26531_, _10089_);
  and (_26537_, _26536_, _04694_);
  and (_26538_, _26537_, _26535_);
  and (_26539_, _10248_, _03839_);
  or (_26540_, _26539_, _08456_);
  nor (_26541_, _26540_, _26538_);
  and (_26542_, _08456_, _10089_);
  or (_26543_, _26542_, _26541_);
  nand (_26544_, _26543_, _10541_);
  and (_26546_, _10540_, _03437_);
  nor (_26547_, _26546_, _03745_);
  nand (_26548_, _26547_, _26544_);
  and (_26549_, _03745_, _03405_);
  nor (_26550_, _26549_, _03483_);
  nand (_26551_, _26550_, _26548_);
  and (_26552_, _04077_, _03483_);
  nor (_26553_, _26552_, _10145_);
  nand (_26554_, _26553_, _26551_);
  and (_26555_, _08783_, _03405_);
  and (_26557_, _26374_, _10146_);
  or (_26558_, _26557_, _26555_);
  and (_26559_, _26558_, _10145_);
  nor (_26560_, _26559_, _10587_);
  and (_26561_, _26560_, _26554_);
  or (_26562_, _26561_, _26346_);
  nand (_26563_, _26562_, _10589_);
  nor (_26564_, _10589_, _03405_);
  nor (_26565_, _26564_, _03838_);
  and (_26566_, _26565_, _26563_);
  and (_26568_, _10248_, _03838_);
  or (_26569_, _26568_, _03959_);
  nor (_26570_, _26569_, _26566_);
  and (_26571_, _03959_, _10089_);
  or (_26572_, _26571_, _26570_);
  nand (_26573_, _26572_, _25690_);
  and (_26574_, _04077_, _03486_);
  nor (_26575_, _26574_, _10601_);
  nand (_26576_, _26575_, _26573_);
  nor (_26577_, _26374_, _10146_);
  nor (_26579_, _08783_, _03405_);
  nor (_26580_, _26579_, _10602_);
  not (_26581_, _26580_);
  nor (_26582_, _26581_, _26577_);
  nor (_26583_, _26582_, _10616_);
  and (_26584_, _26583_, _26576_);
  or (_26585_, _26584_, _26345_);
  nand (_26586_, _26585_, _10614_);
  nor (_26587_, _10614_, _03405_);
  nor (_26588_, _26587_, _03866_);
  and (_26590_, _26588_, _26586_);
  and (_26591_, _10248_, _03866_);
  or (_26592_, _26591_, _03967_);
  nor (_26593_, _26592_, _26590_);
  and (_26594_, _03967_, _10089_);
  or (_26595_, _26594_, _26593_);
  nand (_26596_, _26595_, _25686_);
  and (_26597_, _04077_, _03477_);
  nor (_26598_, _26597_, _10029_);
  nand (_26599_, _26598_, _26596_);
  nor (_26601_, _26374_, \oc8051_golden_model_1.PSW [7]);
  nor (_26602_, _03405_, _08059_);
  nor (_26603_, _26602_, _10030_);
  not (_26604_, _26603_);
  nor (_26605_, _26604_, _26601_);
  nor (_26606_, _26605_, _10628_);
  and (_26607_, _26606_, _26599_);
  or (_26608_, _26607_, _26344_);
  nand (_26609_, _26608_, _08527_);
  nor (_26610_, _08527_, _03405_);
  nor (_26612_, _26610_, _03835_);
  and (_26613_, _26612_, _26609_);
  and (_26614_, _10248_, _03835_);
  or (_26615_, _26614_, _03954_);
  nor (_26616_, _26615_, _26613_);
  and (_26617_, _03954_, _10089_);
  or (_26618_, _26617_, _26616_);
  nand (_26619_, _26618_, _25683_);
  and (_26620_, _04077_, _03481_);
  nor (_26621_, _26620_, _10014_);
  nand (_26623_, _26621_, _26619_);
  nor (_26624_, _26374_, _08059_);
  nor (_26625_, _03405_, \oc8051_golden_model_1.PSW [7]);
  nor (_26626_, _26625_, _10015_);
  not (_26627_, _26626_);
  nor (_26628_, _26627_, _26624_);
  nor (_26629_, _26628_, _10646_);
  and (_26630_, _26629_, _26623_);
  or (_26631_, _26630_, _26343_);
  nand (_26632_, _26631_, _10010_);
  nor (_26634_, _10010_, _03405_);
  nor (_26635_, _26634_, _08006_);
  nand (_26636_, _26635_, _26632_);
  and (_26637_, _08006_, _03461_);
  nor (_26638_, _26637_, _03974_);
  and (_26639_, _26638_, _26636_);
  and (_26640_, _06789_, _03974_);
  or (_26641_, _26640_, _26639_);
  nand (_26642_, _26641_, _06543_);
  and (_26643_, _04077_, _03474_);
  nor (_26645_, _26643_, _03831_);
  nand (_26646_, _26645_, _26642_);
  nor (_26647_, _10248_, _10860_);
  and (_26648_, _26437_, _10860_);
  or (_26649_, _26648_, _04386_);
  nor (_26650_, _26649_, _26647_);
  nor (_26651_, _26650_, _10669_);
  and (_26652_, _26651_, _26646_);
  or (_26653_, _26652_, _26342_);
  nand (_26654_, _26653_, _09989_);
  nor (_26656_, _09989_, _03405_);
  nor (_26657_, _26656_, _07964_);
  nand (_26658_, _26657_, _26654_);
  and (_26659_, _07964_, _03461_);
  nor (_26660_, _26659_, _03707_);
  and (_26661_, _26660_, _26658_);
  and (_26662_, _06789_, _03707_);
  or (_26663_, _26662_, _26661_);
  nand (_26664_, _26663_, _03395_);
  and (_26665_, _04077_, _03394_);
  nor (_26667_, _26665_, _03705_);
  nand (_26668_, _26667_, _26664_);
  nor (_26669_, _26389_, _10860_);
  and (_26670_, _10249_, _10860_);
  nor (_26671_, _26670_, _26669_);
  and (_26672_, _26671_, _03705_);
  nor (_26673_, _26672_, _10888_);
  nand (_26674_, _26673_, _26668_);
  nor (_26675_, _10887_, _03461_);
  nor (_26676_, _26675_, _03703_);
  and (_26678_, _26676_, _26674_);
  or (_26679_, _26678_, _26341_);
  nand (_26680_, _26679_, _10894_);
  nor (_26681_, _10894_, _03462_);
  nor (_26682_, _26681_, _05156_);
  nand (_26683_, _26682_, _26680_);
  and (_26684_, _05156_, _04077_);
  nor (_26685_, _26684_, _03384_);
  nand (_26686_, _26685_, _26683_);
  and (_26687_, _26671_, _03384_);
  nor (_26689_, _26687_, _10911_);
  nand (_26690_, _26689_, _26686_);
  nor (_26691_, _10910_, _03461_);
  nor (_26692_, _26691_, _03701_);
  and (_26693_, _26692_, _26690_);
  or (_26694_, _26693_, _26340_);
  nand (_26695_, _26694_, _10917_);
  nor (_26696_, _10917_, _03462_);
  nor (_26697_, _26696_, _25672_);
  nand (_26698_, _26697_, _26695_);
  and (_26700_, _25672_, _04077_);
  nor (_26701_, _26700_, _10928_);
  and (_26702_, _26701_, _26698_);
  or (_26703_, _26702_, _26339_);
  or (_26704_, _26703_, _42912_);
  or (_26705_, _42908_, \oc8051_golden_model_1.PC [2]);
  and (_26706_, _26705_, _41654_);
  and (_43271_, _26706_, _26704_);
  and (_26707_, _03701_, _03516_);
  and (_26708_, _03703_, _03516_);
  nor (_26710_, _10008_, _03881_);
  and (_26711_, _06744_, _03974_);
  nor (_26712_, _10012_, _03881_);
  nor (_26713_, _10027_, _03881_);
  nor (_26714_, _10612_, _03881_);
  nor (_26715_, _10585_, _03881_);
  nor (_26716_, _06305_, _03516_);
  nor (_26717_, _10488_, _03881_);
  nor (_26718_, _26075_, _03516_);
  or (_26719_, _10246_, _10245_);
  and (_26721_, _26719_, _10262_);
  nor (_26722_, _26719_, _10262_);
  nor (_26723_, _26722_, _26721_);
  and (_26724_, _26723_, _10316_);
  and (_26725_, _10314_, _10243_);
  or (_26726_, _26725_, _26724_);
  and (_26727_, _26726_, _03757_);
  or (_26728_, _10344_, _03881_);
  nand (_26729_, _04944_, _03095_);
  or (_26730_, _04944_, _03881_);
  and (_26732_, _26730_, _26729_);
  or (_26733_, _26732_, _04615_);
  nand (_26734_, _04615_, _03879_);
  and (_26735_, _26734_, _04235_);
  and (_26736_, _26735_, _26733_);
  and (_26737_, _04234_, _03881_);
  or (_26738_, _26737_, _26736_);
  and (_26739_, _26738_, _04948_);
  nor (_26740_, _04948_, _03946_);
  or (_26741_, _26740_, _25715_);
  or (_26743_, _26741_, _26739_);
  and (_26744_, _26743_, _26728_);
  or (_26745_, _26744_, _10320_);
  and (_26746_, _10326_, _03516_);
  or (_26747_, _10088_, _10087_);
  and (_26748_, _26747_, _10101_);
  nor (_26749_, _26747_, _10101_);
  nor (_26750_, _26749_, _26748_);
  and (_26751_, _26750_, _10324_);
  or (_26752_, _26751_, _06140_);
  or (_26754_, _26752_, _26746_);
  and (_26755_, _26754_, _26745_);
  or (_26756_, _26755_, _04624_);
  nand (_26757_, _04624_, _03530_);
  and (_26758_, _26757_, _04630_);
  and (_26759_, _26758_, _26756_);
  or (_26760_, _26759_, _10355_);
  or (_26761_, _26760_, _26727_);
  or (_26762_, _10354_, _03881_);
  and (_26763_, _26762_, _03697_);
  and (_26765_, _26763_, _26761_);
  and (_26766_, _03696_, _03516_);
  or (_26767_, _26766_, _04933_);
  or (_26768_, _26767_, _26765_);
  nand (_26769_, _03946_, _04933_);
  and (_26770_, _26769_, _04537_);
  and (_26771_, _26770_, _26768_);
  nand (_26772_, _03755_, _03516_);
  nand (_26773_, _26772_, _10364_);
  or (_26774_, _26773_, _26771_);
  or (_26776_, _10364_, _03881_);
  and (_26777_, _26776_, _03751_);
  and (_26778_, _26777_, _26774_);
  nand (_26779_, _03750_, _03516_);
  nand (_26780_, _26779_, _10375_);
  or (_26781_, _26780_, _26778_);
  or (_26782_, _10375_, _03881_);
  and (_26783_, _26782_, _03692_);
  and (_26784_, _26783_, _26781_);
  and (_26785_, _03691_, _03516_);
  or (_26787_, _26785_, _10379_);
  or (_26788_, _26787_, _26784_);
  nand (_26789_, _03946_, _10379_);
  and (_26790_, _26789_, _04759_);
  and (_26791_, _26790_, _26788_);
  nand (_26792_, _10423_, _10244_);
  or (_26793_, _26723_, _10423_);
  and (_26794_, _26793_, _26792_);
  and (_26795_, _26794_, _10386_);
  and (_26796_, _03690_, _03516_);
  or (_26798_, _26796_, _10387_);
  or (_26799_, _26798_, _26795_);
  or (_26800_, _26799_, _26791_);
  or (_26801_, _26794_, _10388_);
  and (_26802_, _26801_, _26800_);
  nor (_26803_, _26802_, _03854_);
  and (_26804_, _10243_, _10181_);
  not (_26805_, _26723_);
  nor (_26806_, _26805_, _10181_);
  or (_26807_, _26806_, _03855_);
  or (_26809_, _26807_, _26804_);
  nand (_26810_, _26809_, _10433_);
  or (_26811_, _26810_, _26803_);
  or (_26812_, _26723_, _10446_);
  nand (_26813_, _10446_, _10244_);
  and (_26814_, _26813_, _03847_);
  and (_26815_, _26814_, _26812_);
  and (_26816_, _10462_, _10243_);
  nor (_26817_, _26805_, _10462_);
  nor (_26818_, _26817_, _26816_);
  nor (_26819_, _26818_, _04216_);
  nor (_26820_, _26819_, _26815_);
  and (_26821_, _10431_, _03881_);
  nor (_26822_, _26821_, _03684_);
  and (_26823_, _26822_, _26820_);
  nand (_26824_, _26823_, _26811_);
  and (_26825_, _03684_, _03879_);
  nor (_26826_, _26825_, _05105_);
  nand (_26827_, _26826_, _26824_);
  nor (_26828_, _03946_, _03442_);
  nor (_26831_, _26828_, _26076_);
  and (_26832_, _26831_, _26827_);
  or (_26833_, _26832_, _26718_);
  nand (_26834_, _26833_, _10477_);
  nor (_26835_, _10477_, _03881_);
  nor (_26836_, _26835_, _03811_);
  nand (_26837_, _26836_, _26834_);
  and (_26838_, _03811_, _03516_);
  nor (_26839_, _26838_, _25787_);
  nand (_26840_, _26839_, _26837_);
  and (_26842_, _03946_, _25787_);
  nor (_26843_, _26842_, _03810_);
  nand (_26844_, _26843_, _26840_);
  and (_26845_, _03810_, _03516_);
  nor (_26846_, _26845_, _10494_);
  and (_26847_, _26846_, _26844_);
  or (_26848_, _26847_, _26717_);
  nand (_26849_, _26848_, _10492_);
  nor (_26850_, _10492_, _03516_);
  nor (_26851_, _26850_, _03547_);
  and (_26853_, _26851_, _26849_);
  nor (_26854_, _03422_, _03530_);
  or (_26855_, _26854_, _03679_);
  nor (_26856_, _26855_, _26853_);
  and (_26857_, _03679_, _03879_);
  or (_26858_, _26857_, _26856_);
  nand (_26859_, _26858_, _03418_);
  and (_26860_, _03946_, _03676_);
  nor (_26861_, _26860_, _03861_);
  nand (_26862_, _26861_, _26859_);
  and (_26864_, _10243_, _03861_);
  nor (_26865_, _26864_, _11528_);
  nand (_26866_, _26865_, _26862_);
  nor (_26867_, _10510_, _03516_);
  nor (_26868_, _26867_, _07559_);
  nand (_26869_, _26868_, _26866_);
  nor (_26870_, _10244_, _03415_);
  nor (_26871_, _26870_, _10521_);
  nand (_26872_, _26871_, _26869_);
  nor (_26873_, _10517_, _03881_);
  nor (_26875_, _26873_, _03746_);
  and (_26876_, _26875_, _26872_);
  and (_26877_, _03746_, _03516_);
  or (_26878_, _26877_, _03487_);
  or (_26879_, _26878_, _26876_);
  and (_26880_, _03946_, _03487_);
  nor (_26881_, _26880_, _10525_);
  nand (_26882_, _26881_, _26879_);
  and (_26883_, _26750_, _10525_);
  nor (_26884_, _26883_, _06306_);
  and (_26886_, _26884_, _26882_);
  or (_26887_, _26886_, _26716_);
  nand (_26888_, _26887_, _04694_);
  and (_26889_, _10244_, _03839_);
  nor (_26890_, _26889_, _08456_);
  nand (_26891_, _26890_, _26888_);
  and (_26892_, _08456_, _03516_);
  nor (_26893_, _26892_, _10540_);
  nand (_26894_, _26893_, _26891_);
  nor (_26895_, _10541_, _03526_);
  nor (_26897_, _26895_, _03745_);
  and (_26898_, _26897_, _26894_);
  and (_26899_, _03745_, _03516_);
  or (_26900_, _26899_, _03483_);
  or (_26901_, _26900_, _26898_);
  and (_26902_, _03946_, _03483_);
  nor (_26903_, _26902_, _10145_);
  nand (_26904_, _26903_, _26901_);
  nor (_26905_, _26750_, _08783_);
  nand (_26906_, _08783_, _03879_);
  nand (_26908_, _26906_, _10145_);
  or (_26909_, _26908_, _26905_);
  and (_26910_, _26909_, _10585_);
  and (_26911_, _26910_, _26904_);
  or (_26912_, _26911_, _26715_);
  nand (_26913_, _26912_, _10589_);
  nor (_26914_, _10589_, _03516_);
  nor (_26915_, _26914_, _03838_);
  and (_26916_, _26915_, _26913_);
  and (_26917_, _10243_, _03838_);
  or (_26919_, _26917_, _03959_);
  nor (_26920_, _26919_, _26916_);
  and (_26921_, _03959_, _03879_);
  or (_26922_, _26921_, _26920_);
  nand (_26923_, _26922_, _25690_);
  and (_26924_, _03946_, _03486_);
  nor (_26925_, _26924_, _10601_);
  nand (_26926_, _26925_, _26923_);
  nor (_26927_, _26750_, _10146_);
  nor (_26928_, _08783_, _03516_);
  nor (_26929_, _26928_, _10602_);
  not (_26930_, _26929_);
  nor (_26931_, _26930_, _26927_);
  nor (_26932_, _26931_, _10616_);
  and (_26933_, _26932_, _26926_);
  or (_26934_, _26933_, _26714_);
  nand (_26935_, _26934_, _10614_);
  nor (_26936_, _10614_, _03516_);
  nor (_26937_, _26936_, _03866_);
  and (_26938_, _26937_, _26935_);
  and (_26941_, _10243_, _03866_);
  or (_26942_, _26941_, _03967_);
  nor (_26943_, _26942_, _26938_);
  and (_26944_, _03967_, _03879_);
  or (_26945_, _26944_, _26943_);
  nand (_26946_, _26945_, _25686_);
  and (_26947_, _03946_, _03477_);
  nor (_26948_, _26947_, _10029_);
  nand (_26949_, _26948_, _26946_);
  nor (_26950_, _26750_, \oc8051_golden_model_1.PSW [7]);
  nor (_26952_, _03516_, _08059_);
  nor (_26953_, _26952_, _10030_);
  not (_26954_, _26953_);
  nor (_26955_, _26954_, _26950_);
  nor (_26956_, _26955_, _10628_);
  and (_26957_, _26956_, _26949_);
  or (_26958_, _26957_, _26713_);
  nand (_26959_, _26958_, _08527_);
  nor (_26960_, _08527_, _03516_);
  nor (_26961_, _26960_, _03835_);
  and (_26963_, _26961_, _26959_);
  and (_26964_, _10243_, _03835_);
  or (_26965_, _26964_, _03954_);
  nor (_26966_, _26965_, _26963_);
  and (_26967_, _03954_, _03879_);
  or (_26968_, _26967_, _26966_);
  nand (_26969_, _26968_, _25683_);
  and (_26970_, _03946_, _03481_);
  nor (_26971_, _26970_, _10014_);
  nand (_26972_, _26971_, _26969_);
  nor (_26974_, _26750_, _08059_);
  nor (_26975_, _03516_, \oc8051_golden_model_1.PSW [7]);
  nor (_26976_, _26975_, _10015_);
  not (_26977_, _26976_);
  nor (_26978_, _26977_, _26974_);
  nor (_26979_, _26978_, _10646_);
  and (_26980_, _26979_, _26972_);
  or (_26981_, _26980_, _26712_);
  nand (_26982_, _26981_, _10010_);
  nor (_26983_, _10010_, _03516_);
  nor (_26985_, _26983_, _08006_);
  nand (_26986_, _26985_, _26982_);
  and (_26987_, _08006_, _03881_);
  nor (_26988_, _26987_, _03974_);
  and (_26989_, _26988_, _26986_);
  or (_26990_, _26989_, _26711_);
  nand (_26991_, _26990_, _06543_);
  and (_26992_, _03946_, _03474_);
  nor (_26993_, _26992_, _03831_);
  nand (_26994_, _26993_, _26991_);
  and (_26996_, _26805_, _10860_);
  nor (_26997_, _10243_, _10860_);
  or (_26998_, _26997_, _04386_);
  nor (_26999_, _26998_, _26996_);
  nor (_27000_, _26999_, _10669_);
  and (_27001_, _27000_, _26994_);
  or (_27002_, _27001_, _26710_);
  nand (_27003_, _27002_, _09989_);
  nor (_27004_, _09989_, _03516_);
  nor (_27005_, _27004_, _07964_);
  and (_27007_, _27005_, _27003_);
  and (_27008_, _07964_, _03881_);
  or (_27009_, _27008_, _03707_);
  nor (_27010_, _27009_, _27007_);
  and (_27011_, _06744_, _03707_);
  or (_27012_, _27011_, _27010_);
  nand (_27013_, _27012_, _03395_);
  and (_27014_, _03946_, _03394_);
  nor (_27015_, _27014_, _03705_);
  nand (_27016_, _27015_, _27013_);
  nor (_27018_, _26723_, _10860_);
  and (_27019_, _10244_, _10860_);
  nor (_27020_, _27019_, _27018_);
  and (_27021_, _27020_, _03705_);
  nor (_27022_, _27021_, _10888_);
  nand (_27023_, _27022_, _27016_);
  nor (_27024_, _10887_, _03881_);
  nor (_27025_, _27024_, _03703_);
  and (_27026_, _27025_, _27023_);
  or (_27027_, _27026_, _26708_);
  nand (_27029_, _27027_, _10894_);
  nor (_27030_, _10894_, _03530_);
  nor (_27031_, _27030_, _05156_);
  nand (_27032_, _27031_, _27029_);
  and (_27033_, _05156_, _03946_);
  nor (_27034_, _27033_, _03384_);
  nand (_27035_, _27034_, _27032_);
  and (_27036_, _27020_, _03384_);
  nor (_27037_, _27036_, _10911_);
  nand (_27038_, _27037_, _27035_);
  nor (_27040_, _10910_, _03881_);
  nor (_27041_, _27040_, _03701_);
  and (_27042_, _27041_, _27038_);
  or (_27043_, _27042_, _26707_);
  nand (_27044_, _27043_, _10917_);
  nor (_27045_, _10917_, _03530_);
  nor (_27046_, _27045_, _25672_);
  nand (_27047_, _27046_, _27044_);
  and (_27048_, _25672_, _03946_);
  nor (_27049_, _27048_, _10928_);
  and (_27051_, _27049_, _27047_);
  and (_27052_, _10928_, _03881_);
  or (_27053_, _27052_, _27051_);
  or (_27054_, _27053_, _42912_);
  or (_27055_, _42908_, \oc8051_golden_model_1.PC [3]);
  and (_27056_, _27055_, _41654_);
  and (_43272_, _27056_, _27054_);
  and (_27057_, _09991_, \oc8051_golden_model_1.PC [4]);
  nor (_27058_, _09991_, \oc8051_golden_model_1.PC [4]);
  nor (_27059_, _27058_, _27057_);
  nor (_27061_, _27059_, _10910_);
  and (_27062_, _06339_, _03394_);
  and (_27063_, _10084_, _08783_);
  and (_27064_, _10106_, _10103_);
  nor (_27065_, _27064_, _10107_);
  and (_27066_, _27065_, _10146_);
  or (_27067_, _27066_, _27063_);
  and (_27068_, _27067_, _10145_);
  nor (_27069_, _10084_, _06305_);
  and (_27070_, _10084_, _03810_);
  nor (_27072_, _26075_, _10084_);
  and (_27073_, _10239_, _10181_);
  and (_27074_, _10267_, _10264_);
  nor (_27075_, _27074_, _10268_);
  not (_27076_, _27075_);
  nor (_27077_, _27076_, _10181_);
  or (_27078_, _27077_, _03855_);
  or (_27079_, _27078_, _27073_);
  nand (_27080_, _10085_, _03691_);
  or (_27081_, _27059_, _10360_);
  or (_27083_, _25971_, _10239_);
  or (_27084_, _27075_, _26387_);
  and (_27085_, _27084_, _03757_);
  and (_27086_, _27085_, _27083_);
  nand (_27087_, _06339_, _04111_);
  nand (_27088_, _10085_, _04109_);
  and (_27089_, _04944_, \oc8051_golden_model_1.PC [4]);
  or (_27090_, _27089_, _04615_);
  and (_27091_, _27090_, _04235_);
  not (_27092_, _27059_);
  nor (_27094_, _27092_, _04944_);
  or (_27095_, _27094_, _27091_);
  and (_27096_, _27095_, _27088_);
  and (_27097_, _27059_, _04234_);
  or (_27098_, _27097_, _04111_);
  or (_27099_, _27098_, _27096_);
  and (_27100_, _27099_, _10344_);
  and (_27101_, _27100_, _27087_);
  nor (_27102_, _27092_, _10344_);
  or (_27103_, _27102_, _10320_);
  or (_27105_, _27103_, _27101_);
  and (_27106_, _27065_, _10324_);
  and (_27107_, _10326_, _10084_);
  or (_27108_, _27107_, _27106_);
  or (_27109_, _27108_, _06140_);
  and (_27110_, _27109_, _27105_);
  or (_27111_, _27110_, _04624_);
  and (_27112_, _27111_, _04630_);
  or (_27113_, _27112_, _10355_);
  or (_27114_, _27113_, _27086_);
  and (_27116_, _27114_, _27081_);
  or (_27117_, _27116_, _03696_);
  nand (_27118_, _10085_, _03696_);
  and (_27119_, _27118_, _03445_);
  and (_27120_, _27119_, _27117_);
  nor (_27121_, _06339_, _03445_);
  or (_27122_, _27121_, _03755_);
  or (_27123_, _27122_, _27120_);
  nand (_27124_, _10085_, _03755_);
  and (_27125_, _27124_, _10364_);
  and (_27127_, _27125_, _27123_);
  nor (_27128_, _27092_, _10364_);
  or (_27129_, _27128_, _03750_);
  or (_27130_, _27129_, _27127_);
  nand (_27131_, _10085_, _03750_);
  and (_27132_, _27131_, _10375_);
  and (_27133_, _27132_, _27130_);
  nor (_27134_, _27092_, _10375_);
  or (_27135_, _27134_, _03691_);
  or (_27136_, _27135_, _27133_);
  and (_27138_, _27136_, _27080_);
  or (_27139_, _27138_, _10379_);
  nand (_27140_, _06339_, _10379_);
  and (_27141_, _27140_, _04759_);
  and (_27142_, _27141_, _27139_);
  and (_27143_, _10084_, _03690_);
  or (_27144_, _27143_, _10387_);
  or (_27145_, _27144_, _27142_);
  nand (_27146_, _10423_, _10240_);
  or (_27147_, _27075_, _10423_);
  and (_27148_, _27147_, _27146_);
  and (_27149_, _27148_, _26041_);
  or (_27150_, _27149_, _10388_);
  and (_27151_, _27150_, _27145_);
  and (_27152_, _27148_, _10386_);
  or (_27153_, _27152_, _03854_);
  or (_27154_, _27153_, _27151_);
  and (_27155_, _27154_, _27079_);
  nand (_27156_, _27155_, _10433_);
  and (_27157_, _10446_, _10239_);
  not (_27160_, _10446_);
  and (_27161_, _27075_, _27160_);
  or (_27162_, _27161_, _27157_);
  and (_27163_, _27162_, _03847_);
  and (_27164_, _10462_, _10239_);
  nor (_27165_, _27076_, _10462_);
  nor (_27166_, _27165_, _27164_);
  nor (_27167_, _27166_, _04216_);
  nor (_27168_, _27167_, _27163_);
  and (_27169_, _27059_, _10431_);
  nor (_27171_, _27169_, _03684_);
  and (_27172_, _27171_, _27168_);
  nand (_27173_, _27172_, _27156_);
  and (_27174_, _10085_, _03684_);
  nor (_27175_, _27174_, _05105_);
  nand (_27176_, _27175_, _27173_);
  nor (_27177_, _06339_, _03442_);
  nor (_27178_, _27177_, _26076_);
  and (_27179_, _27178_, _27176_);
  or (_27180_, _27179_, _27072_);
  nand (_27182_, _27180_, _10477_);
  nor (_27183_, _27059_, _10477_);
  nor (_27184_, _27183_, _03811_);
  nand (_27185_, _27184_, _27182_);
  and (_27186_, _10084_, _03811_);
  nor (_27187_, _27186_, _25787_);
  nand (_27188_, _27187_, _27185_);
  and (_27189_, _06339_, _25787_);
  nor (_27190_, _27189_, _03810_);
  and (_27191_, _27190_, _27188_);
  or (_27193_, _27191_, _27070_);
  nand (_27194_, _27193_, _10488_);
  nor (_27195_, _27092_, _10488_);
  nor (_27196_, _27195_, _10493_);
  nand (_27197_, _27196_, _27194_);
  nor (_27198_, _10084_, _10492_);
  nor (_27199_, _27198_, _03547_);
  and (_27200_, _27199_, _27197_);
  nor (_27201_, _27092_, _03422_);
  or (_27202_, _27201_, _03679_);
  nor (_27204_, _27202_, _27200_);
  and (_27205_, _10085_, _03679_);
  or (_27206_, _27205_, _27204_);
  nand (_27207_, _27206_, _03418_);
  and (_27208_, _06339_, _03676_);
  nor (_27209_, _27208_, _03861_);
  nand (_27210_, _27209_, _27207_);
  and (_27211_, _10239_, _03861_);
  nor (_27212_, _27211_, _11528_);
  nand (_27213_, _27212_, _27210_);
  nor (_27215_, _10510_, _10084_);
  nor (_27216_, _27215_, _07559_);
  and (_27217_, _27216_, _27213_);
  nor (_27218_, _10240_, _03415_);
  nor (_27219_, _27218_, _27217_);
  nand (_27220_, _27219_, _10517_);
  nor (_27221_, _27059_, _10517_);
  nor (_27222_, _27221_, _03746_);
  nand (_27223_, _27222_, _27220_);
  nor (_27224_, _10084_, _03487_);
  or (_27226_, _27224_, _10519_);
  nand (_27227_, _27226_, _27223_);
  and (_27228_, _06339_, _03487_);
  nor (_27229_, _27228_, _10525_);
  nand (_27230_, _27229_, _27227_);
  and (_27231_, _27065_, _10525_);
  nor (_27232_, _27231_, _06306_);
  and (_27233_, _27232_, _27230_);
  or (_27234_, _27233_, _27069_);
  nand (_27235_, _27234_, _04694_);
  and (_27237_, _10240_, _03839_);
  nor (_27238_, _27237_, _08456_);
  nand (_27239_, _27238_, _27235_);
  and (_27240_, _10084_, _08456_);
  nor (_27241_, _27240_, _10540_);
  nand (_27242_, _27241_, _27239_);
  and (_27243_, _10558_, _10555_);
  nor (_27244_, _27243_, _10559_);
  nor (_27245_, _27244_, _10541_);
  nor (_27246_, _27245_, _03745_);
  nand (_27248_, _27246_, _27242_);
  and (_27249_, _10084_, _03745_);
  nor (_27250_, _27249_, _03483_);
  nand (_27251_, _27250_, _27248_);
  and (_27252_, _06339_, _03483_);
  nor (_27253_, _27252_, _10145_);
  and (_27254_, _27253_, _27251_);
  or (_27255_, _27254_, _27068_);
  nand (_27256_, _27255_, _10585_);
  nor (_27257_, _27092_, _10585_);
  nor (_27259_, _27257_, _10590_);
  nand (_27260_, _27259_, _27256_);
  nor (_27261_, _10589_, _10084_);
  nor (_27262_, _27261_, _03838_);
  and (_27263_, _27262_, _27260_);
  and (_27264_, _10239_, _03838_);
  or (_27265_, _27264_, _03959_);
  nor (_27266_, _27265_, _27263_);
  and (_27267_, _10085_, _03959_);
  or (_27268_, _27267_, _27266_);
  nand (_27270_, _27268_, _25690_);
  and (_27271_, _06339_, _03486_);
  nor (_27272_, _27271_, _10601_);
  nand (_27273_, _27272_, _27270_);
  or (_27274_, _10085_, _08783_);
  nand (_27275_, _27065_, _08783_);
  and (_27276_, _27275_, _27274_);
  or (_27277_, _27276_, _10602_);
  nand (_27278_, _27277_, _27273_);
  nand (_27279_, _27278_, _10612_);
  nor (_27281_, _27092_, _10612_);
  nor (_27282_, _27281_, _10615_);
  nand (_27283_, _27282_, _27279_);
  nor (_27284_, _10084_, _10614_);
  nor (_27285_, _27284_, _03866_);
  nand (_27286_, _27285_, _27283_);
  and (_27287_, _10239_, _03866_);
  nor (_27288_, _27287_, _03967_);
  and (_27289_, _27288_, _27286_);
  and (_27290_, _10085_, _03967_);
  or (_27292_, _27290_, _27289_);
  nand (_27293_, _27292_, _25686_);
  and (_27294_, _06339_, _03477_);
  nor (_27295_, _27294_, _10029_);
  nand (_27296_, _27295_, _27293_);
  nand (_27297_, _10084_, \oc8051_golden_model_1.PSW [7]);
  nand (_27298_, _27065_, _08059_);
  and (_27299_, _27298_, _27297_);
  or (_27300_, _27299_, _10030_);
  nand (_27301_, _27300_, _27296_);
  nand (_27303_, _27301_, _10027_);
  nor (_27304_, _27092_, _10027_);
  nor (_27305_, _27304_, _08528_);
  nand (_27306_, _27305_, _27303_);
  nor (_27307_, _10084_, _08527_);
  nor (_27308_, _27307_, _03835_);
  nand (_27309_, _27308_, _27306_);
  and (_27310_, _10239_, _03835_);
  nor (_27311_, _27310_, _03954_);
  and (_27312_, _27311_, _27309_);
  and (_27314_, _10085_, _03954_);
  or (_27315_, _27314_, _27312_);
  nand (_27316_, _27315_, _25683_);
  and (_27317_, _06339_, _03481_);
  nor (_27318_, _27317_, _10014_);
  nand (_27319_, _27318_, _27316_);
  nand (_27320_, _10084_, _08059_);
  nand (_27321_, _27065_, \oc8051_golden_model_1.PSW [7]);
  and (_27322_, _27321_, _27320_);
  or (_27323_, _27322_, _10015_);
  nand (_27325_, _27323_, _27319_);
  nand (_27326_, _27325_, _10012_);
  nor (_27327_, _27092_, _10012_);
  nor (_27328_, _27327_, _10011_);
  nand (_27329_, _27328_, _27326_);
  nor (_27330_, _10084_, _10010_);
  nor (_27331_, _27330_, _08006_);
  nand (_27332_, _27331_, _27329_);
  and (_27333_, _27059_, _08006_);
  nor (_27334_, _27333_, _03974_);
  and (_27336_, _27334_, _27332_);
  and (_27337_, _06881_, _03974_);
  or (_27338_, _27337_, _27336_);
  nand (_27339_, _27338_, _06543_);
  and (_27340_, _06339_, _03474_);
  nor (_27341_, _27340_, _03831_);
  and (_27342_, _27341_, _27339_);
  nor (_27343_, _10240_, _10860_);
  and (_27344_, _27075_, _10860_);
  nor (_27345_, _27344_, _27343_);
  nor (_27347_, _27345_, _04386_);
  or (_27348_, _27347_, _27342_);
  nand (_27349_, _27348_, _10008_);
  nor (_27350_, _27092_, _10008_);
  nor (_27351_, _27350_, _09990_);
  nand (_27352_, _27351_, _27349_);
  nor (_27353_, _10084_, _09989_);
  nor (_27354_, _27353_, _07964_);
  nand (_27355_, _27354_, _27352_);
  and (_27356_, _27059_, _07964_);
  nor (_27358_, _27356_, _03707_);
  and (_27359_, _27358_, _27355_);
  and (_27360_, _06881_, _03707_);
  or (_27361_, _27360_, _27359_);
  and (_27362_, _27361_, _03395_);
  or (_27363_, _27362_, _27062_);
  nand (_27364_, _27363_, _03706_);
  and (_27365_, _10240_, _10860_);
  nor (_27366_, _27075_, _10860_);
  nor (_27367_, _27366_, _27365_);
  nor (_27369_, _27367_, _03706_);
  nor (_27370_, _27369_, _10888_);
  nand (_27371_, _27370_, _27364_);
  nor (_27372_, _27092_, _10887_);
  nor (_27373_, _27372_, _03703_);
  nand (_27374_, _27373_, _27371_);
  not (_27375_, _10894_);
  and (_27376_, _10085_, _03703_);
  nor (_27377_, _27376_, _27375_);
  nand (_27378_, _27377_, _27374_);
  nor (_27380_, _27092_, _10894_);
  nor (_27381_, _27380_, _05156_);
  nand (_27382_, _27381_, _27378_);
  and (_27383_, _06339_, _05156_);
  nor (_27384_, _27383_, _03384_);
  nand (_27385_, _27384_, _27382_);
  and (_27386_, _27367_, _03384_);
  nor (_27387_, _27386_, _10911_);
  and (_27388_, _27387_, _27385_);
  or (_27389_, _27388_, _27061_);
  nand (_27391_, _27389_, _03702_);
  and (_27392_, _10085_, _03701_);
  nor (_27393_, _27392_, _26323_);
  nand (_27394_, _27393_, _27391_);
  nor (_27395_, _27092_, _10917_);
  nor (_27396_, _27395_, _25672_);
  nand (_27397_, _27396_, _27394_);
  and (_27398_, _25672_, _06339_);
  nor (_27399_, _27398_, _10928_);
  and (_27400_, _27399_, _27397_);
  and (_27402_, _27059_, _10928_);
  or (_27403_, _27402_, _27400_);
  or (_27404_, _27403_, _42912_);
  or (_27405_, _42908_, \oc8051_golden_model_1.PC [4]);
  and (_27406_, _27405_, _41654_);
  and (_43273_, _27406_, _27404_);
  nor (_27407_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_27408_, _10079_, _03129_);
  nor (_27409_, _27408_, _27407_);
  and (_27410_, _27409_, _10928_);
  and (_27411_, _10079_, _03701_);
  nor (_27412_, _27409_, _10894_);
  or (_27413_, _27409_, _10008_);
  or (_27414_, _06941_, _11621_);
  or (_27415_, _27409_, _10012_);
  or (_27416_, _27409_, _10027_);
  or (_27417_, _27409_, _10612_);
  or (_27418_, _27409_, _10585_);
  nand (_27419_, _10080_, _03745_);
  or (_27420_, _10079_, _06305_);
  or (_27423_, _26075_, _10079_);
  nand (_27424_, _10235_, _10181_);
  or (_27425_, _10237_, _10236_);
  not (_27426_, _27425_);
  nor (_27427_, _27426_, _10269_);
  and (_27428_, _27426_, _10269_);
  nor (_27429_, _27428_, _27427_);
  not (_27430_, _27429_);
  or (_27431_, _27430_, _10181_);
  and (_27432_, _27431_, _03854_);
  and (_27434_, _27432_, _27424_);
  nand (_27435_, _10080_, _03696_);
  or (_27436_, _27409_, _10360_);
  and (_27437_, _10314_, _10234_);
  and (_27438_, _27430_, _10316_);
  or (_27439_, _27438_, _27437_);
  and (_27440_, _27439_, _03757_);
  or (_27441_, _10082_, _10081_);
  nand (_27442_, _27441_, _10108_);
  or (_27443_, _27441_, _10108_);
  and (_27445_, _27443_, _27442_);
  and (_27446_, _27445_, _10324_);
  and (_27447_, _10326_, _10079_);
  or (_27448_, _27447_, _27446_);
  and (_27449_, _27448_, _10320_);
  nand (_27450_, _06370_, _04111_);
  and (_27451_, _10344_, _04948_);
  not (_27452_, _27451_);
  or (_27453_, _27409_, _25708_);
  nand (_27454_, _10080_, _04109_);
  nor (_27456_, _04615_, \oc8051_golden_model_1.PC [5]);
  nand (_27457_, _27456_, _04944_);
  and (_27458_, _27457_, _27454_);
  or (_27459_, _27458_, _04234_);
  and (_27460_, _27459_, _27453_);
  or (_27461_, _27460_, _27452_);
  or (_27462_, _27409_, _10344_);
  and (_27463_, _27462_, _06140_);
  and (_27464_, _27463_, _27461_);
  and (_27465_, _27464_, _27450_);
  or (_27467_, _27465_, _04624_);
  or (_27468_, _27467_, _27449_);
  and (_27469_, _27468_, _04630_);
  or (_27470_, _27469_, _10355_);
  or (_27471_, _27470_, _27440_);
  and (_27472_, _27471_, _27436_);
  or (_27473_, _27472_, _03696_);
  and (_27474_, _27473_, _27435_);
  or (_27475_, _27474_, _04933_);
  nand (_27476_, _06370_, _04933_);
  and (_27478_, _27476_, _04537_);
  and (_27479_, _27478_, _27475_);
  nand (_27480_, _10079_, _03755_);
  nand (_27481_, _27480_, _10364_);
  or (_27482_, _27481_, _27479_);
  or (_27483_, _27409_, _10364_);
  and (_27484_, _27483_, _03751_);
  and (_27485_, _27484_, _27482_);
  nand (_27486_, _10079_, _03750_);
  nand (_27487_, _27486_, _10375_);
  or (_27489_, _27487_, _27485_);
  or (_27490_, _27409_, _10375_);
  and (_27491_, _27490_, _03692_);
  and (_27492_, _27491_, _27489_);
  and (_27493_, _10079_, _03691_);
  or (_27494_, _27493_, _10379_);
  or (_27495_, _27494_, _27492_);
  nand (_27496_, _06370_, _10379_);
  and (_27497_, _27496_, _04759_);
  and (_27498_, _27497_, _27495_);
  or (_27500_, _27430_, _10423_);
  nand (_27501_, _10423_, _10235_);
  and (_27502_, _27501_, _27500_);
  and (_27503_, _27502_, _10386_);
  and (_27504_, _10079_, _03690_);
  or (_27505_, _27504_, _10387_);
  or (_27506_, _27505_, _27503_);
  or (_27507_, _27506_, _27498_);
  or (_27508_, _27502_, _10388_);
  and (_27509_, _27508_, _03855_);
  and (_27511_, _27509_, _27507_);
  or (_27512_, _27511_, _27434_);
  and (_27513_, _27512_, _10433_);
  nand (_27514_, _27429_, _27160_);
  nand (_27515_, _10446_, _10235_);
  and (_27516_, _27515_, _03847_);
  and (_27517_, _27516_, _27514_);
  and (_27518_, _10462_, _10234_);
  nor (_27519_, _27429_, _10462_);
  or (_27520_, _27519_, _27518_);
  and (_27522_, _27520_, _03773_);
  or (_27523_, _27522_, _27517_);
  and (_27524_, _27409_, _10431_);
  or (_27525_, _27524_, _03684_);
  or (_27526_, _27525_, _27523_);
  or (_27527_, _27526_, _27513_);
  nand (_27528_, _10080_, _03684_);
  and (_27529_, _27528_, _03442_);
  and (_27530_, _27529_, _27527_);
  nor (_27531_, _06370_, _03442_);
  or (_27533_, _27531_, _26076_);
  or (_27534_, _27533_, _27530_);
  and (_27535_, _27534_, _27423_);
  or (_27536_, _27535_, _10481_);
  or (_27537_, _27409_, _10477_);
  and (_27538_, _27537_, _11667_);
  and (_27539_, _27538_, _27536_);
  and (_27540_, _10079_, _03811_);
  or (_27541_, _27540_, _25787_);
  or (_27542_, _27541_, _27539_);
  nand (_27544_, _06370_, _25787_);
  and (_27545_, _27544_, _11666_);
  and (_27546_, _27545_, _27542_);
  nand (_27547_, _10079_, _03810_);
  nand (_27548_, _27547_, _10488_);
  or (_27549_, _27548_, _27546_);
  or (_27550_, _27409_, _10488_);
  and (_27551_, _27550_, _27549_);
  or (_27552_, _27551_, _10493_);
  or (_27553_, _10079_, _10492_);
  and (_27555_, _27553_, _03422_);
  and (_27556_, _27555_, _27552_);
  and (_27557_, _27409_, _03547_);
  or (_27558_, _27557_, _03679_);
  or (_27559_, _27558_, _27556_);
  nand (_27560_, _10080_, _03679_);
  and (_27561_, _27560_, _27559_);
  or (_27562_, _27561_, _03676_);
  nand (_27563_, _06370_, _03676_);
  and (_27564_, _27563_, _09806_);
  and (_27566_, _27564_, _27562_);
  nand (_27567_, _10234_, _03861_);
  nand (_27568_, _27567_, _10510_);
  or (_27569_, _27568_, _27566_);
  or (_27570_, _10510_, _10079_);
  and (_27571_, _27570_, _03415_);
  and (_27572_, _27571_, _27569_);
  or (_27573_, _10235_, _03415_);
  nand (_27574_, _27573_, _10517_);
  or (_27575_, _27574_, _27572_);
  not (_27577_, _03746_);
  or (_27578_, _27409_, _10517_);
  and (_27579_, _27578_, _27577_);
  and (_27580_, _27579_, _27575_);
  nor (_27581_, _10079_, _03487_);
  nor (_27582_, _27581_, _10519_);
  or (_27583_, _27582_, _27580_);
  nand (_27584_, _06370_, _03487_);
  and (_27585_, _27584_, _10526_);
  and (_27586_, _27585_, _27583_);
  and (_27588_, _27445_, _10525_);
  or (_27589_, _27588_, _06306_);
  or (_27590_, _27589_, _27586_);
  and (_27591_, _27590_, _27420_);
  or (_27592_, _27591_, _03839_);
  nand (_27593_, _10235_, _03839_);
  and (_27594_, _27593_, _08457_);
  and (_27595_, _27594_, _27592_);
  and (_27596_, _10079_, _08456_);
  or (_27597_, _27596_, _27595_);
  and (_27599_, _27597_, _10541_);
  or (_27600_, _10553_, _10552_);
  or (_27601_, _27600_, _10560_);
  nand (_27602_, _27600_, _10560_);
  and (_27603_, _27602_, _10540_);
  and (_27604_, _27603_, _27601_);
  or (_27605_, _27604_, _03745_);
  or (_27606_, _27605_, _27599_);
  and (_27607_, _27606_, _27419_);
  or (_27608_, _27607_, _03483_);
  nand (_27610_, _06370_, _03483_);
  and (_27611_, _27610_, _10580_);
  and (_27612_, _27611_, _27608_);
  or (_27613_, _27445_, _08783_);
  or (_27614_, _10079_, _10146_);
  and (_27615_, _27614_, _10145_);
  and (_27616_, _27615_, _27613_);
  or (_27617_, _27616_, _10587_);
  or (_27618_, _27617_, _27612_);
  and (_27619_, _27618_, _27418_);
  or (_27621_, _27619_, _10590_);
  or (_27622_, _10589_, _10079_);
  and (_27623_, _27622_, _04703_);
  and (_27624_, _27623_, _27621_);
  and (_27625_, _10234_, _03838_);
  or (_27626_, _27625_, _03959_);
  or (_27627_, _27626_, _27624_);
  nand (_27628_, _10080_, _03959_);
  and (_27629_, _27628_, _27627_);
  or (_27630_, _27629_, _03486_);
  nand (_27632_, _06370_, _03486_);
  and (_27633_, _27632_, _10602_);
  and (_27634_, _27633_, _27630_);
  or (_27635_, _27445_, _10146_);
  or (_27636_, _10079_, _08783_);
  and (_27637_, _27636_, _10601_);
  and (_27638_, _27637_, _27635_);
  or (_27639_, _27638_, _10616_);
  or (_27640_, _27639_, _27634_);
  and (_27641_, _27640_, _27417_);
  or (_27643_, _27641_, _10615_);
  or (_27644_, _10079_, _10614_);
  and (_27645_, _27644_, _04708_);
  and (_27646_, _27645_, _27643_);
  and (_27647_, _10234_, _03866_);
  or (_27648_, _27647_, _03967_);
  or (_27649_, _27648_, _27646_);
  nand (_27650_, _10080_, _03967_);
  and (_27651_, _27650_, _27649_);
  or (_27652_, _27651_, _03477_);
  nand (_27654_, _06370_, _03477_);
  and (_27655_, _27654_, _10030_);
  and (_27656_, _27655_, _27652_);
  or (_27657_, _27445_, \oc8051_golden_model_1.PSW [7]);
  or (_27658_, _10079_, _08059_);
  and (_27659_, _27658_, _10029_);
  and (_27660_, _27659_, _27657_);
  or (_27661_, _27660_, _10628_);
  or (_27662_, _27661_, _27656_);
  and (_27663_, _27662_, _27416_);
  or (_27665_, _27663_, _08528_);
  or (_27666_, _10079_, _08527_);
  and (_27667_, _27666_, _06532_);
  and (_27668_, _27667_, _27665_);
  and (_27669_, _10234_, _03835_);
  or (_27670_, _27669_, _03954_);
  or (_27671_, _27670_, _27668_);
  nand (_27672_, _10080_, _03954_);
  and (_27673_, _27672_, _27671_);
  or (_27674_, _27673_, _03481_);
  nand (_27676_, _06370_, _03481_);
  and (_27677_, _27676_, _10015_);
  and (_27678_, _27677_, _27674_);
  or (_27679_, _27445_, _08059_);
  or (_27680_, _10079_, \oc8051_golden_model_1.PSW [7]);
  and (_27681_, _27680_, _10014_);
  and (_27682_, _27681_, _27679_);
  or (_27683_, _27682_, _10646_);
  or (_27684_, _27683_, _27678_);
  and (_27685_, _27684_, _27415_);
  or (_27687_, _27685_, _10011_);
  or (_27688_, _10079_, _10010_);
  and (_27689_, _27688_, _08007_);
  and (_27690_, _27689_, _27687_);
  and (_27691_, _27409_, _08006_);
  or (_27692_, _27691_, _03974_);
  or (_27693_, _27692_, _27690_);
  and (_27694_, _27693_, _27414_);
  or (_27695_, _27694_, _03474_);
  nand (_27696_, _06370_, _03474_);
  and (_27697_, _27696_, _04386_);
  and (_27698_, _27697_, _27695_);
  or (_27699_, _10234_, _10860_);
  nand (_27700_, _27429_, _10860_);
  and (_27701_, _27700_, _03831_);
  and (_27702_, _27701_, _27699_);
  or (_27703_, _27702_, _10669_);
  or (_27704_, _27703_, _27698_);
  and (_27705_, _27704_, _27413_);
  or (_27706_, _27705_, _09990_);
  or (_27709_, _10079_, _09989_);
  and (_27710_, _27709_, _10870_);
  and (_27711_, _27710_, _27706_);
  and (_27712_, _27409_, _07964_);
  or (_27713_, _27712_, _03707_);
  or (_27714_, _27713_, _27711_);
  or (_27715_, _06941_, _03708_);
  and (_27716_, _27715_, _27714_);
  or (_27717_, _27716_, _03394_);
  nand (_27718_, _06370_, _03394_);
  and (_27720_, _27718_, _03706_);
  and (_27721_, _27720_, _27717_);
  and (_27722_, _10235_, _10860_);
  nor (_27723_, _27430_, _10860_);
  nor (_27724_, _27723_, _27722_);
  and (_27725_, _27724_, _03705_);
  or (_27726_, _27725_, _10888_);
  or (_27727_, _27726_, _27721_);
  or (_27728_, _27409_, _10887_);
  and (_27729_, _27728_, _03704_);
  and (_27731_, _27729_, _27727_);
  and (_27732_, _10079_, _03703_);
  nor (_27733_, _27732_, _27375_);
  not (_27734_, _27733_);
  nor (_27735_, _27734_, _27731_);
  nor (_27736_, _27735_, _27412_);
  nor (_27737_, _27736_, _05156_);
  and (_27738_, _06370_, _05156_);
  nor (_27739_, _27738_, _03384_);
  not (_27740_, _27739_);
  nor (_27742_, _27740_, _27737_);
  and (_27743_, _27724_, _03384_);
  nor (_27744_, _27743_, _10911_);
  not (_27745_, _27744_);
  nor (_27746_, _27745_, _27742_);
  nor (_27747_, _27409_, _10910_);
  nor (_27748_, _27747_, _03701_);
  not (_27749_, _27748_);
  nor (_27750_, _27749_, _27746_);
  nor (_27751_, _27750_, _27411_);
  nor (_27753_, _27751_, _26323_);
  and (_27754_, _27409_, _26323_);
  nor (_27755_, _27754_, _25672_);
  not (_27756_, _27755_);
  or (_27757_, _27756_, _27753_);
  and (_27758_, _25672_, _06370_);
  nor (_27759_, _27758_, _10928_);
  and (_27760_, _27759_, _27757_);
  or (_27761_, _27760_, _27410_);
  or (_27762_, _27761_, _42912_);
  or (_27764_, _42908_, \oc8051_golden_model_1.PC [5]);
  and (_27765_, _27764_, _41654_);
  and (_43274_, _27765_, _27762_);
  and (_27766_, _06023_, _09991_);
  nor (_27767_, _27766_, \oc8051_golden_model_1.PC [6]);
  nor (_27768_, _27767_, _09992_);
  and (_27769_, _27768_, _10928_);
  and (_27770_, _06406_, _05156_);
  not (_27771_, _27768_);
  and (_27772_, _27771_, _07964_);
  and (_27774_, _10227_, _03835_);
  and (_27775_, _10227_, _03866_);
  and (_27776_, _10227_, _03838_);
  nor (_27777_, _10071_, _06305_);
  and (_27778_, _10072_, _03746_);
  and (_27779_, _27771_, _10431_);
  and (_27780_, _10423_, _10226_);
  and (_27781_, _10271_, _10231_);
  nor (_27782_, _27781_, _10272_);
  not (_27783_, _27782_);
  nor (_27785_, _27783_, _10423_);
  or (_27786_, _27785_, _27780_);
  nor (_27787_, _27786_, _10388_);
  and (_27788_, _10072_, _03691_);
  nor (_27789_, _27768_, _10360_);
  or (_27790_, _10316_, _10227_);
  or (_27791_, _27783_, _10314_);
  nand (_27792_, _27791_, _27790_);
  nand (_27793_, _27792_, _03757_);
  and (_27794_, _06406_, _04111_);
  nor (_27796_, _27768_, _25708_);
  and (_27797_, _10072_, _04109_);
  nor (_27798_, _04615_, \oc8051_golden_model_1.PC [6]);
  and (_27799_, _27798_, _04944_);
  nor (_27800_, _27799_, _27797_);
  nor (_27801_, _27800_, _04234_);
  nor (_27802_, _27801_, _27796_);
  nor (_27803_, _27802_, _04111_);
  nor (_27804_, _27803_, _25715_);
  not (_27805_, _27804_);
  nor (_27807_, _27805_, _27794_);
  nor (_27808_, _27771_, _10344_);
  nor (_27809_, _27808_, _10320_);
  not (_27810_, _27809_);
  nor (_27811_, _27810_, _27807_);
  and (_27812_, _10110_, _10076_);
  nor (_27813_, _27812_, _10111_);
  and (_27814_, _27813_, _10324_);
  and (_27815_, _10326_, _10071_);
  nor (_27816_, _27815_, _27814_);
  and (_27818_, _27816_, _10320_);
  or (_27819_, _27818_, _27811_);
  nand (_27820_, _27819_, _04625_);
  nand (_27821_, _27820_, _04630_);
  and (_27822_, _27821_, _10354_);
  and (_27823_, _27822_, _27793_);
  or (_27824_, _27823_, _27789_);
  nand (_27825_, _27824_, _03697_);
  and (_27826_, _10072_, _03696_);
  nor (_27827_, _27826_, _04933_);
  nand (_27829_, _27827_, _27825_);
  nor (_27830_, _06406_, _03445_);
  nor (_27831_, _27830_, _03755_);
  and (_27832_, _27831_, _27829_);
  and (_27833_, _10072_, _03755_);
  or (_27834_, _27833_, _27832_);
  and (_27835_, _27834_, _10364_);
  nor (_27836_, _27768_, _10364_);
  or (_27837_, _27836_, _27835_);
  nand (_27838_, _27837_, _03751_);
  and (_27840_, _10072_, _03750_);
  nor (_27841_, _27840_, _10377_);
  nand (_27842_, _27841_, _27838_);
  nor (_27843_, _27771_, _10375_);
  nor (_27844_, _27843_, _03691_);
  and (_27845_, _27844_, _27842_);
  or (_27846_, _27845_, _27788_);
  nand (_27847_, _27846_, _03448_);
  and (_27848_, _06406_, _10379_);
  nor (_27849_, _27848_, _03690_);
  nand (_27851_, _27849_, _27847_);
  and (_27852_, _10071_, _03690_);
  nor (_27853_, _27852_, _10425_);
  and (_27854_, _27853_, _27851_);
  or (_27855_, _27854_, _27787_);
  nand (_27856_, _27855_, _03855_);
  and (_27857_, _10226_, _10181_);
  nor (_27858_, _27783_, _10181_);
  or (_27859_, _27858_, _27857_);
  nor (_27860_, _27859_, _03855_);
  nor (_27862_, _27860_, _03773_);
  nand (_27863_, _27862_, _27856_);
  nor (_27864_, _27782_, _10462_);
  and (_27865_, _10462_, _10227_);
  or (_27866_, _27865_, _04216_);
  or (_27867_, _27866_, _27864_);
  nand (_27868_, _27867_, _27863_);
  nand (_27869_, _27868_, _11721_);
  and (_27870_, _10446_, _10226_);
  and (_27871_, _27782_, _27160_);
  or (_27873_, _27871_, _27870_);
  and (_27874_, _27873_, _03847_);
  nor (_27875_, _27874_, _10431_);
  and (_27876_, _27875_, _27869_);
  or (_27877_, _27876_, _27779_);
  nand (_27878_, _27877_, _03685_);
  and (_27879_, _10072_, _03684_);
  nor (_27880_, _27879_, _05105_);
  nand (_27881_, _27880_, _27878_);
  nor (_27882_, _06406_, _03442_);
  nor (_27884_, _27882_, _26076_);
  and (_27885_, _27884_, _27881_);
  nor (_27886_, _26075_, _10071_);
  or (_27887_, _27886_, _27885_);
  nand (_27888_, _27887_, _10477_);
  nor (_27889_, _27768_, _10477_);
  nor (_27890_, _27889_, _03811_);
  nand (_27891_, _27890_, _27888_);
  and (_27892_, _10071_, _03811_);
  nor (_27893_, _27892_, _25787_);
  and (_27895_, _27893_, _27891_);
  and (_27896_, _06406_, _25787_);
  nor (_27897_, _27896_, _27895_);
  and (_27898_, _27897_, _11666_);
  and (_27899_, _10071_, _03810_);
  or (_27900_, _27899_, _10494_);
  or (_27901_, _27900_, _27898_);
  nor (_27902_, _27768_, _10488_);
  nor (_27903_, _27902_, _10493_);
  and (_27904_, _27903_, _27901_);
  nor (_27906_, _10072_, _10492_);
  or (_27907_, _27906_, _03547_);
  nor (_27908_, _27907_, _27904_);
  nor (_27909_, _27768_, _03422_);
  or (_27910_, _27909_, _27908_);
  nand (_27911_, _27910_, _03680_);
  and (_27912_, _10072_, _03679_);
  nor (_27913_, _27912_, _03676_);
  nand (_27914_, _27913_, _27911_);
  nor (_27915_, _06406_, _03418_);
  nor (_27917_, _27915_, _03861_);
  nand (_27918_, _27917_, _27914_);
  and (_27919_, _10227_, _03861_);
  nor (_27920_, _27919_, _11528_);
  nand (_27921_, _27920_, _27918_);
  nor (_27922_, _10510_, _10072_);
  nor (_27923_, _27922_, _07559_);
  nand (_27924_, _27923_, _27921_);
  nor (_27925_, _10226_, _03415_);
  nor (_27926_, _27925_, _10521_);
  nand (_27928_, _27926_, _27924_);
  nor (_27929_, _27771_, _10517_);
  nor (_27930_, _27929_, _03746_);
  and (_27931_, _27930_, _27928_);
  nor (_27932_, _27931_, _27778_);
  or (_27933_, _27932_, _03487_);
  and (_27934_, _06406_, _03487_);
  nor (_27935_, _27934_, _10525_);
  nand (_27936_, _27935_, _27933_);
  and (_27937_, _27813_, _10525_);
  nor (_27939_, _27937_, _06306_);
  and (_27940_, _27939_, _27936_);
  or (_27941_, _27940_, _27777_);
  nand (_27942_, _27941_, _04694_);
  and (_27943_, _10227_, _03839_);
  nor (_27944_, _27943_, _08456_);
  nand (_27945_, _27944_, _27942_);
  and (_27946_, _10071_, _08456_);
  nor (_27947_, _27946_, _10540_);
  nand (_27948_, _27947_, _27945_);
  and (_27950_, _10562_, _10551_);
  nor (_27951_, _27950_, _10563_);
  nor (_27952_, _27951_, _10541_);
  nor (_27953_, _27952_, _03745_);
  nand (_27954_, _27953_, _27948_);
  and (_27955_, _10071_, _03745_);
  nor (_27956_, _27955_, _03483_);
  nand (_27957_, _27956_, _27954_);
  and (_27958_, _06406_, _03483_);
  nor (_27959_, _27958_, _10145_);
  nand (_27961_, _27959_, _27957_);
  and (_27962_, _10071_, _08783_);
  and (_27963_, _27813_, _10146_);
  or (_27964_, _27963_, _27962_);
  and (_27965_, _27964_, _10145_);
  nor (_27966_, _27965_, _10587_);
  nand (_27967_, _27966_, _27961_);
  nor (_27968_, _27768_, _10585_);
  nor (_27969_, _27968_, _10590_);
  nand (_27970_, _27969_, _27967_);
  nor (_27972_, _10589_, _10072_);
  nor (_27973_, _27972_, _03838_);
  and (_27974_, _27973_, _27970_);
  or (_27975_, _27974_, _27776_);
  nand (_27976_, _27975_, _04701_);
  and (_27977_, _10072_, _03959_);
  nor (_27978_, _27977_, _03486_);
  and (_27979_, _27978_, _27976_);
  nor (_27980_, _06406_, _25690_);
  or (_27981_, _27980_, _27979_);
  nand (_27983_, _27981_, _10602_);
  nor (_27984_, _27813_, _10146_);
  nor (_27985_, _10071_, _08783_);
  nor (_27986_, _27985_, _10602_);
  not (_27987_, _27986_);
  nor (_27988_, _27987_, _27984_);
  nor (_27989_, _27988_, _10616_);
  nand (_27990_, _27989_, _27983_);
  nor (_27991_, _27768_, _10612_);
  nor (_27992_, _27991_, _10615_);
  nand (_27994_, _27992_, _27990_);
  nor (_27995_, _10072_, _10614_);
  nor (_27996_, _27995_, _03866_);
  and (_27997_, _27996_, _27994_);
  or (_27998_, _27997_, _27775_);
  nand (_27999_, _27998_, _04706_);
  and (_28000_, _10072_, _03967_);
  nor (_28001_, _28000_, _03477_);
  and (_28002_, _28001_, _27999_);
  nor (_28003_, _06406_, _25686_);
  or (_28005_, _28003_, _28002_);
  nand (_28006_, _28005_, _10030_);
  nor (_28007_, _27813_, \oc8051_golden_model_1.PSW [7]);
  nor (_28008_, _10071_, _08059_);
  nor (_28009_, _28008_, _10030_);
  not (_28010_, _28009_);
  nor (_28011_, _28010_, _28007_);
  nor (_28012_, _28011_, _10628_);
  nand (_28013_, _28012_, _28006_);
  nor (_28014_, _27768_, _10027_);
  nor (_28016_, _28014_, _08528_);
  nand (_28017_, _28016_, _28013_);
  nor (_28018_, _10072_, _08527_);
  nor (_28019_, _28018_, _03835_);
  and (_28020_, _28019_, _28017_);
  or (_28021_, _28020_, _27774_);
  nand (_28022_, _28021_, _06537_);
  and (_28023_, _10072_, _03954_);
  nor (_28024_, _28023_, _03481_);
  and (_28025_, _28024_, _28022_);
  nor (_28027_, _06406_, _25683_);
  or (_28028_, _28027_, _28025_);
  nand (_28029_, _28028_, _10015_);
  nor (_28030_, _27813_, _08059_);
  nor (_28031_, _10071_, \oc8051_golden_model_1.PSW [7]);
  nor (_28032_, _28031_, _10015_);
  not (_28033_, _28032_);
  nor (_28034_, _28033_, _28030_);
  nor (_28035_, _28034_, _10646_);
  nand (_28036_, _28035_, _28029_);
  nor (_28038_, _27768_, _10012_);
  nor (_28039_, _28038_, _10011_);
  nand (_28040_, _28039_, _28036_);
  nor (_28041_, _10072_, _10010_);
  nor (_28042_, _28041_, _08006_);
  nand (_28043_, _28042_, _28040_);
  and (_28044_, _27771_, _08006_);
  nor (_28045_, _28044_, _03974_);
  and (_28046_, _28045_, _28043_);
  and (_28047_, _06933_, _03974_);
  or (_28049_, _28047_, _03474_);
  or (_28050_, _28049_, _28046_);
  and (_28051_, _06406_, _03474_);
  nor (_28052_, _28051_, _03831_);
  nand (_28053_, _28052_, _28050_);
  and (_28054_, _27783_, _10860_);
  nor (_28055_, _10226_, _10860_);
  or (_28056_, _28055_, _04386_);
  nor (_28057_, _28056_, _28054_);
  nor (_28058_, _28057_, _10669_);
  nand (_28060_, _28058_, _28053_);
  nor (_28061_, _27768_, _10008_);
  nor (_28062_, _28061_, _09990_);
  nand (_28063_, _28062_, _28060_);
  nor (_28064_, _10072_, _09989_);
  nor (_28065_, _28064_, _07964_);
  and (_28066_, _28065_, _28063_);
  or (_28067_, _28066_, _27772_);
  nand (_28068_, _28067_, _03708_);
  and (_28069_, _06607_, _03707_);
  nor (_28071_, _28069_, _03394_);
  and (_28072_, _28071_, _28068_);
  nor (_28073_, _06406_, _03395_);
  or (_28074_, _28073_, _03705_);
  nor (_28075_, _28074_, _28072_);
  nor (_28076_, _27782_, _10860_);
  and (_28077_, _10227_, _10860_);
  nor (_28078_, _28077_, _28076_);
  nor (_28079_, _28078_, _03706_);
  or (_28080_, _28079_, _28075_);
  and (_28082_, _28080_, _10887_);
  nor (_28083_, _27768_, _10887_);
  or (_28084_, _28083_, _28082_);
  nand (_28085_, _28084_, _03704_);
  and (_28086_, _10072_, _03703_);
  nor (_28087_, _28086_, _27375_);
  nand (_28088_, _28087_, _28085_);
  nor (_28089_, _27771_, _10894_);
  nor (_28090_, _28089_, _05156_);
  and (_28091_, _28090_, _28088_);
  or (_28093_, _28091_, _27770_);
  nand (_28094_, _28093_, _03385_);
  nor (_28095_, _28078_, _03385_);
  nor (_28096_, _28095_, _10911_);
  nand (_28097_, _28096_, _28094_);
  nor (_28098_, _27771_, _10910_);
  nor (_28099_, _28098_, _03701_);
  nand (_28100_, _28099_, _28097_);
  and (_28101_, _10072_, _03701_);
  nor (_28102_, _28101_, _26323_);
  nand (_28104_, _28102_, _28100_);
  nor (_28105_, _27771_, _10917_);
  nor (_28106_, _28105_, _25672_);
  nand (_28107_, _28106_, _28104_);
  and (_28108_, _25672_, _06406_);
  nor (_28109_, _28108_, _10928_);
  and (_28110_, _28109_, _28107_);
  nor (_28111_, _28110_, _27769_);
  nand (_28112_, _28111_, _42908_);
  or (_28113_, _42908_, \oc8051_golden_model_1.PC [6]);
  and (_28115_, _28113_, _41654_);
  and (_43275_, _28115_, _28112_);
  and (_28116_, _06028_, _03701_);
  and (_28117_, _06028_, _03703_);
  nor (_28118_, _09992_, \oc8051_golden_model_1.PC [7]);
  nor (_28119_, _28118_, _09993_);
  nor (_28120_, _28119_, _10008_);
  nor (_28121_, _28119_, _10012_);
  nor (_28122_, _28119_, _10027_);
  nor (_28123_, _28119_, _10612_);
  nor (_28125_, _28119_, _10585_);
  and (_28126_, _06273_, _03745_);
  nor (_28127_, _06305_, _06028_);
  and (_28128_, _06273_, _03679_);
  nor (_28129_, _28119_, _10488_);
  nor (_28130_, _26075_, _06028_);
  not (_28131_, _28119_);
  and (_28132_, _28131_, _10431_);
  nor (_28133_, _06070_, _03445_);
  and (_28134_, _28131_, _04624_);
  or (_28135_, _10067_, _10068_);
  and (_28136_, _28135_, _10112_);
  nor (_28137_, _28135_, _10112_);
  nor (_28138_, _28137_, _28136_);
  nand (_28139_, _28138_, _10324_);
  or (_28140_, _10324_, _06273_);
  nand (_28141_, _28140_, _28139_);
  nand (_28142_, _28141_, _10320_);
  nand (_28143_, _06070_, _04111_);
  and (_28144_, _25708_, _10344_);
  or (_28147_, _28144_, _28119_);
  nand (_28148_, _06273_, _04109_);
  nor (_28149_, _04615_, \oc8051_golden_model_1.PC [7]);
  nand (_28150_, _28149_, _04944_);
  and (_28151_, _28150_, _28148_);
  nand (_28152_, _27451_, _04235_);
  or (_28153_, _28152_, _28151_);
  and (_28154_, _28153_, _06140_);
  and (_28155_, _28154_, _28147_);
  and (_28156_, _28155_, _28143_);
  nor (_28158_, _28156_, _04624_);
  and (_28159_, _28158_, _28142_);
  nor (_28160_, _28159_, _28134_);
  or (_28161_, _28160_, _03757_);
  and (_28162_, _10314_, _06899_);
  or (_28163_, _10222_, _10223_);
  and (_28164_, _28163_, _10273_);
  nor (_28165_, _28163_, _10273_);
  nor (_28166_, _28165_, _28164_);
  and (_28167_, _28166_, _10316_);
  or (_28169_, _28167_, _28162_);
  or (_28170_, _28169_, _04630_);
  and (_28171_, _28170_, _10354_);
  and (_28172_, _28171_, _28161_);
  nor (_28173_, _28131_, _10354_);
  or (_28174_, _28173_, _03696_);
  or (_28175_, _28174_, _28172_);
  and (_28176_, _06273_, _03696_);
  nor (_28177_, _28176_, _04933_);
  and (_28178_, _28177_, _28175_);
  or (_28180_, _28178_, _28133_);
  nand (_28181_, _28180_, _04537_);
  and (_28182_, _06028_, _03755_);
  nor (_28183_, _28182_, _10365_);
  nand (_28184_, _28183_, _28181_);
  nor (_28185_, _28119_, _10364_);
  nor (_28186_, _28185_, _03750_);
  nand (_28187_, _28186_, _28184_);
  and (_28188_, _06028_, _03750_);
  nor (_28189_, _28188_, _10377_);
  nand (_28191_, _28189_, _28187_);
  nor (_28192_, _28119_, _10375_);
  nor (_28193_, _28192_, _03691_);
  nand (_28194_, _28193_, _28191_);
  and (_28195_, _06028_, _03691_);
  nor (_28196_, _28195_, _10379_);
  nand (_28197_, _28196_, _28194_);
  and (_28198_, _06070_, _10379_);
  nor (_28199_, _28198_, _03690_);
  nand (_28200_, _28199_, _28197_);
  and (_28202_, _06028_, _03690_);
  nor (_28203_, _28202_, _10425_);
  and (_28204_, _28203_, _28200_);
  and (_28205_, _10423_, _06899_);
  not (_28206_, _28166_);
  nor (_28207_, _28206_, _10423_);
  or (_28208_, _28207_, _28205_);
  nor (_28209_, _28208_, _10388_);
  or (_28210_, _28209_, _28204_);
  nand (_28211_, _28210_, _03855_);
  and (_28213_, _10181_, _06899_);
  nor (_28214_, _28206_, _10181_);
  or (_28215_, _28214_, _03855_);
  nor (_28216_, _28215_, _28213_);
  nor (_28217_, _28216_, _03773_);
  nand (_28218_, _28217_, _28211_);
  nor (_28219_, _28166_, _10462_);
  and (_28220_, _10462_, _06900_);
  or (_28221_, _28220_, _04216_);
  or (_28222_, _28221_, _28219_);
  nand (_28224_, _28222_, _28218_);
  nand (_28225_, _28224_, _11721_);
  and (_28226_, _10446_, _06899_);
  and (_28227_, _28166_, _27160_);
  or (_28228_, _28227_, _28226_);
  and (_28229_, _28228_, _03847_);
  nor (_28230_, _28229_, _10431_);
  and (_28231_, _28230_, _28225_);
  or (_28232_, _28231_, _28132_);
  nand (_28233_, _28232_, _03685_);
  and (_28235_, _06273_, _03684_);
  nor (_28236_, _28235_, _05105_);
  nand (_28237_, _28236_, _28233_);
  nor (_28238_, _06070_, _03442_);
  nor (_28239_, _28238_, _26076_);
  and (_28240_, _28239_, _28237_);
  or (_28241_, _28240_, _28130_);
  nand (_28242_, _28241_, _10477_);
  nor (_28243_, _28119_, _10477_);
  nor (_28244_, _28243_, _03811_);
  nand (_28246_, _28244_, _28242_);
  and (_28247_, _06028_, _03811_);
  nor (_28248_, _28247_, _25787_);
  nand (_28249_, _28248_, _28246_);
  and (_28250_, _06070_, _25787_);
  nor (_28251_, _28250_, _03810_);
  nand (_28252_, _28251_, _28249_);
  and (_28253_, _06028_, _03810_);
  nor (_28254_, _28253_, _10494_);
  and (_28255_, _28254_, _28252_);
  or (_28257_, _28255_, _28129_);
  nand (_28258_, _28257_, _10492_);
  nor (_28259_, _10492_, _06028_);
  nor (_28260_, _28259_, _03547_);
  nand (_28261_, _28260_, _28258_);
  nor (_28262_, _28131_, _03422_);
  nor (_28263_, _28262_, _03679_);
  and (_28264_, _28263_, _28261_);
  or (_28265_, _28264_, _28128_);
  nand (_28266_, _28265_, _03418_);
  and (_28268_, _06070_, _03676_);
  nor (_28269_, _28268_, _03861_);
  nand (_28270_, _28269_, _28266_);
  and (_28271_, _06899_, _03861_);
  nor (_28272_, _28271_, _11528_);
  nand (_28273_, _28272_, _28270_);
  nor (_28274_, _10510_, _06028_);
  nor (_28275_, _28274_, _07559_);
  nand (_28276_, _28275_, _28273_);
  nor (_28277_, _06900_, _03415_);
  nor (_28279_, _28277_, _10521_);
  nand (_28280_, _28279_, _28276_);
  nor (_28281_, _28119_, _10517_);
  nor (_28282_, _28281_, _03746_);
  and (_28283_, _28282_, _28280_);
  and (_28284_, _06028_, _03746_);
  or (_28285_, _28284_, _03487_);
  or (_28286_, _28285_, _28283_);
  and (_28287_, _06070_, _03487_);
  nor (_28288_, _28287_, _10525_);
  nand (_28290_, _28288_, _28286_);
  and (_28291_, _28138_, _10525_);
  nor (_28292_, _28291_, _06306_);
  and (_28293_, _28292_, _28290_);
  or (_28294_, _28293_, _28127_);
  nand (_28295_, _28294_, _04694_);
  and (_28296_, _06900_, _03839_);
  nor (_28297_, _28296_, _08456_);
  and (_28298_, _28297_, _28295_);
  and (_28299_, _08456_, _06028_);
  or (_28301_, _28299_, _28298_);
  nand (_28302_, _28301_, _10541_);
  or (_28303_, _10547_, _10546_);
  nor (_28304_, _28303_, _10564_);
  and (_28305_, _28303_, _10564_);
  or (_28306_, _28305_, _10541_);
  or (_28307_, _28306_, _28304_);
  and (_28308_, _28307_, _04336_);
  and (_28309_, _28308_, _28302_);
  or (_28310_, _28309_, _28126_);
  nand (_28312_, _28310_, _11594_);
  and (_28313_, _06070_, _03483_);
  nor (_28314_, _28313_, _10145_);
  nand (_28315_, _28314_, _28312_);
  and (_28316_, _08783_, _06028_);
  and (_28317_, _28138_, _10146_);
  or (_28318_, _28317_, _28316_);
  and (_28319_, _28318_, _10145_);
  nor (_28320_, _28319_, _10587_);
  and (_28321_, _28320_, _28315_);
  or (_28322_, _28321_, _28125_);
  nand (_28323_, _28322_, _10589_);
  nor (_28324_, _10589_, _06028_);
  nor (_28325_, _28324_, _03838_);
  and (_28326_, _28325_, _28323_);
  and (_28327_, _06899_, _03838_);
  or (_28328_, _28327_, _03959_);
  nor (_28329_, _28328_, _28326_);
  and (_28330_, _06273_, _03959_);
  or (_28331_, _28330_, _28329_);
  nand (_28334_, _28331_, _25690_);
  and (_28335_, _06070_, _03486_);
  nor (_28336_, _28335_, _10601_);
  nand (_28337_, _28336_, _28334_);
  nor (_28338_, _28138_, _10146_);
  nor (_28339_, _08783_, _06028_);
  nor (_28340_, _28339_, _10602_);
  not (_28341_, _28340_);
  nor (_28342_, _28341_, _28338_);
  nor (_28343_, _28342_, _10616_);
  and (_28345_, _28343_, _28337_);
  or (_28346_, _28345_, _28123_);
  nand (_28347_, _28346_, _10614_);
  nor (_28348_, _10614_, _06028_);
  nor (_28349_, _28348_, _03866_);
  and (_28350_, _28349_, _28347_);
  and (_28351_, _06899_, _03866_);
  or (_28352_, _28351_, _03967_);
  nor (_28353_, _28352_, _28350_);
  and (_28354_, _06273_, _03967_);
  or (_28356_, _28354_, _28353_);
  nand (_28357_, _28356_, _25686_);
  and (_28358_, _06070_, _03477_);
  nor (_28359_, _28358_, _10029_);
  nand (_28360_, _28359_, _28357_);
  nor (_28361_, _28138_, \oc8051_golden_model_1.PSW [7]);
  nor (_28362_, _06028_, _08059_);
  nor (_28363_, _28362_, _10030_);
  not (_28364_, _28363_);
  nor (_28365_, _28364_, _28361_);
  nor (_28367_, _28365_, _10628_);
  and (_28368_, _28367_, _28360_);
  or (_28369_, _28368_, _28122_);
  nand (_28370_, _28369_, _08527_);
  nor (_28371_, _08527_, _06028_);
  nor (_28372_, _28371_, _03835_);
  and (_28373_, _28372_, _28370_);
  and (_28374_, _06899_, _03835_);
  or (_28375_, _28374_, _03954_);
  nor (_28376_, _28375_, _28373_);
  and (_28378_, _06273_, _03954_);
  or (_28379_, _28378_, _28376_);
  nand (_28380_, _28379_, _25683_);
  and (_28381_, _06070_, _03481_);
  nor (_28382_, _28381_, _10014_);
  nand (_28383_, _28382_, _28380_);
  nor (_28384_, _28138_, _08059_);
  nor (_28385_, _06028_, \oc8051_golden_model_1.PSW [7]);
  nor (_28386_, _28385_, _10015_);
  not (_28387_, _28386_);
  nor (_28389_, _28387_, _28384_);
  nor (_28390_, _28389_, _10646_);
  and (_28391_, _28390_, _28383_);
  or (_28392_, _28391_, _28121_);
  nand (_28393_, _28392_, _10010_);
  nor (_28394_, _10010_, _06028_);
  nor (_28395_, _28394_, _08006_);
  nand (_28396_, _28395_, _28393_);
  and (_28397_, _28119_, _08006_);
  nor (_28398_, _28397_, _03974_);
  and (_28400_, _28398_, _28396_);
  and (_28401_, _06280_, _03974_);
  or (_28402_, _28401_, _28400_);
  nand (_28403_, _28402_, _06543_);
  and (_28404_, _06070_, _03474_);
  nor (_28405_, _28404_, _03831_);
  nand (_28406_, _28405_, _28403_);
  and (_28407_, _28206_, _10860_);
  nor (_28408_, _06899_, _10860_);
  or (_28409_, _28408_, _04386_);
  or (_28411_, _28409_, _28407_);
  and (_28412_, _28411_, _10008_);
  and (_28413_, _28412_, _28406_);
  or (_28414_, _28413_, _28120_);
  nand (_28415_, _28414_, _09989_);
  nor (_28416_, _09989_, _06028_);
  nor (_28417_, _28416_, _07964_);
  and (_28418_, _28417_, _28415_);
  and (_28419_, _28119_, _07964_);
  or (_28420_, _28419_, _03707_);
  nor (_28422_, _28420_, _28418_);
  and (_28423_, _06280_, _03707_);
  or (_28424_, _28423_, _28422_);
  nand (_28425_, _28424_, _03395_);
  and (_28426_, _06070_, _03394_);
  nor (_28427_, _28426_, _03705_);
  nand (_28428_, _28427_, _28425_);
  and (_28429_, _06900_, _10860_);
  nor (_28430_, _28166_, _10860_);
  nor (_28431_, _28430_, _28429_);
  and (_28433_, _28431_, _03705_);
  nor (_28434_, _28433_, _10888_);
  nand (_28435_, _28434_, _28428_);
  nor (_28436_, _28119_, _10887_);
  nor (_28437_, _28436_, _03703_);
  and (_28438_, _28437_, _28435_);
  or (_28439_, _28438_, _28117_);
  nand (_28440_, _28439_, _10894_);
  nor (_28441_, _28131_, _10894_);
  nor (_28442_, _28441_, _05156_);
  nand (_28444_, _28442_, _28440_);
  and (_28445_, _06070_, _05156_);
  nor (_28446_, _28445_, _03384_);
  nand (_28447_, _28446_, _28444_);
  and (_28448_, _28431_, _03384_);
  nor (_28449_, _28448_, _10911_);
  nand (_28450_, _28449_, _28447_);
  nor (_28451_, _28119_, _10910_);
  nor (_28452_, _28451_, _03701_);
  and (_28453_, _28452_, _28450_);
  or (_28455_, _28453_, _28116_);
  nand (_28456_, _28455_, _10917_);
  nor (_28457_, _28131_, _10917_);
  nor (_28458_, _28457_, _25672_);
  nand (_28459_, _28458_, _28456_);
  and (_28460_, _25672_, _06070_);
  nor (_28461_, _28460_, _10928_);
  and (_28462_, _28461_, _28459_);
  and (_28463_, _28119_, _10928_);
  or (_28464_, _28463_, _28462_);
  or (_28466_, _28464_, _42912_);
  or (_28467_, _42908_, \oc8051_golden_model_1.PC [7]);
  and (_28468_, _28467_, _41654_);
  and (_43276_, _28468_, _28466_);
  nor (_28469_, _04211_, _10921_);
  nor (_28470_, _04211_, _06956_);
  nor (_28471_, _10014_, _03481_);
  and (_28472_, _10278_, _03866_);
  nor (_28473_, _10116_, _06305_);
  and (_28474_, _10116_, _03746_);
  or (_28476_, _26075_, _10116_);
  nor (_28477_, _09993_, \oc8051_golden_model_1.PC [8]);
  nor (_28478_, _28477_, _09994_);
  and (_28479_, _28478_, _10431_);
  nor (_28480_, _10281_, _10275_);
  nor (_28481_, _28480_, _10282_);
  or (_28482_, _28481_, _10446_);
  nand (_28483_, _10446_, _10278_);
  and (_28484_, _28483_, _03847_);
  and (_28485_, _28484_, _28482_);
  or (_28487_, _28481_, _10462_);
  nand (_28488_, _10462_, _10278_);
  and (_28489_, _28488_, _03773_);
  and (_28490_, _28489_, _28487_);
  or (_28491_, _28490_, _28485_);
  or (_28492_, _28491_, _28479_);
  not (_28493_, _28481_);
  nor (_28494_, _28493_, _10181_);
  and (_28495_, _10277_, _10181_);
  or (_28496_, _28495_, _28494_);
  and (_28498_, _28496_, _03854_);
  and (_28499_, _10116_, _03691_);
  nor (_28500_, _25971_, _10278_);
  and (_28501_, _28481_, _10316_);
  or (_28502_, _28501_, _04630_);
  or (_28503_, _28502_, _28500_);
  not (_28504_, _28478_);
  nand (_28505_, _28504_, _04624_);
  nor (_28506_, _10119_, _10114_);
  nor (_28507_, _28506_, _10120_);
  and (_28509_, _28507_, _10324_);
  and (_28510_, _10326_, _10116_);
  or (_28511_, _28510_, _28509_);
  and (_28512_, _28511_, _10320_);
  not (_28513_, _10116_);
  nand (_28514_, _28513_, _04109_);
  nor (_28515_, _04615_, \oc8051_golden_model_1.PC [8]);
  nand (_28516_, _28515_, _04944_);
  and (_28517_, _28516_, _28514_);
  or (_28518_, _28517_, _04234_);
  or (_28520_, _28478_, _25708_);
  and (_28521_, _28520_, _28518_);
  or (_28522_, _28521_, _27452_);
  or (_28523_, _28478_, _10344_);
  and (_28524_, _28523_, _06140_);
  and (_28525_, _28524_, _28522_);
  or (_28526_, _28525_, _04624_);
  or (_28527_, _28526_, _28512_);
  and (_28528_, _28527_, _28505_);
  or (_28529_, _28528_, _03757_);
  and (_28531_, _28529_, _10354_);
  and (_28532_, _28531_, _28503_);
  nor (_28533_, _28504_, _10354_);
  or (_28534_, _28533_, _03696_);
  or (_28535_, _28534_, _28532_);
  and (_28536_, _28513_, _03696_);
  nor (_28537_, _28536_, _10358_);
  and (_28538_, _28537_, _28535_);
  nand (_28539_, _10116_, _03755_);
  nand (_28540_, _28539_, _10364_);
  or (_28542_, _28540_, _28538_);
  or (_28543_, _28478_, _10364_);
  and (_28544_, _28543_, _03751_);
  and (_28545_, _28544_, _28542_);
  nand (_28546_, _10116_, _03750_);
  nand (_28547_, _28546_, _10375_);
  or (_28548_, _28547_, _28545_);
  or (_28549_, _28478_, _10375_);
  and (_28550_, _28549_, _03692_);
  and (_28551_, _28550_, _28548_);
  or (_28553_, _28551_, _28499_);
  and (_28554_, _28553_, _10380_);
  or (_28555_, _28481_, _10423_);
  nand (_28556_, _10423_, _10278_);
  and (_28557_, _28556_, _28555_);
  and (_28558_, _28557_, _10386_);
  and (_28559_, _10116_, _03690_);
  or (_28560_, _28559_, _10387_);
  or (_28561_, _28560_, _28558_);
  or (_28562_, _28561_, _28554_);
  or (_28564_, _28557_, _10388_);
  and (_28565_, _28564_, _03855_);
  and (_28566_, _28565_, _28562_);
  or (_28567_, _28566_, _28498_);
  and (_28568_, _28567_, _10433_);
  or (_28569_, _28568_, _28492_);
  and (_28570_, _28569_, _03685_);
  and (_28571_, _10116_, _03684_);
  nor (_28572_, _28571_, _05105_);
  nand (_28573_, _28572_, _26075_);
  or (_28575_, _28573_, _28570_);
  and (_28576_, _28575_, _28476_);
  or (_28577_, _28576_, _10481_);
  or (_28578_, _28478_, _10477_);
  and (_28579_, _28578_, _11667_);
  and (_28580_, _28579_, _28577_);
  and (_28581_, _10116_, _03811_);
  or (_28582_, _28581_, _25787_);
  or (_28583_, _28582_, _28580_);
  and (_28584_, _28583_, _11666_);
  nand (_28586_, _10116_, _03810_);
  nand (_28587_, _28586_, _10488_);
  or (_28588_, _28587_, _28584_);
  or (_28589_, _28478_, _10488_);
  and (_28590_, _28589_, _10492_);
  and (_28591_, _28590_, _28588_);
  nor (_28592_, _28513_, _10492_);
  or (_28593_, _28592_, _03547_);
  or (_28594_, _28593_, _28591_);
  or (_28595_, _28478_, _03422_);
  and (_28597_, _28595_, _28594_);
  or (_28598_, _28597_, _03679_);
  nand (_28599_, _28513_, _03679_);
  nor (_28600_, _03861_, _03676_);
  and (_28601_, _28600_, _28599_);
  and (_28602_, _28601_, _28598_);
  and (_28603_, _10277_, _03861_);
  or (_28604_, _28603_, _11528_);
  or (_28605_, _28604_, _28602_);
  nor (_28606_, _10510_, _10116_);
  nor (_28608_, _28606_, _07559_);
  nand (_28609_, _28608_, _28605_);
  nor (_28610_, _10278_, _03415_);
  nor (_28611_, _28610_, _10521_);
  nand (_28612_, _28611_, _28609_);
  nor (_28613_, _28478_, _10517_);
  nor (_28614_, _28613_, _03746_);
  and (_28615_, _28614_, _28612_);
  or (_28616_, _28615_, _28474_);
  nand (_28617_, _28616_, _25812_);
  and (_28619_, _28507_, _10525_);
  nor (_28620_, _28619_, _06306_);
  and (_28621_, _28620_, _28617_);
  or (_28622_, _28621_, _28473_);
  nand (_28623_, _28622_, _04694_);
  and (_28624_, _10278_, _03839_);
  nor (_28625_, _28624_, _08456_);
  nand (_28626_, _28625_, _28623_);
  and (_28627_, _10116_, _08456_);
  nor (_28628_, _28627_, _10540_);
  nand (_28630_, _28628_, _28626_);
  and (_28631_, _10566_, _10545_);
  nor (_28632_, _28631_, _10567_);
  nor (_28633_, _28632_, _10541_);
  nor (_28634_, _28633_, _03745_);
  nand (_28635_, _28634_, _28630_);
  and (_28636_, _10116_, _03745_);
  nor (_28637_, _28636_, _03483_);
  nand (_28638_, _28637_, _28635_);
  nand (_28639_, _28638_, _10580_);
  and (_28641_, _10116_, _08783_);
  and (_28642_, _28507_, _10146_);
  or (_28643_, _28642_, _28641_);
  and (_28644_, _28643_, _10145_);
  nor (_28645_, _28644_, _10587_);
  nand (_28646_, _28645_, _28639_);
  nor (_28647_, _28478_, _10585_);
  nor (_28648_, _28647_, _10590_);
  and (_28649_, _28648_, _28646_);
  nor (_28650_, _10589_, _28513_);
  or (_28652_, _28650_, _03838_);
  or (_28653_, _28652_, _28649_);
  and (_28654_, _10278_, _03838_);
  nor (_28655_, _28654_, _03959_);
  nand (_28656_, _28655_, _28653_);
  nor (_28657_, _10116_, _03486_);
  or (_28658_, _28657_, _10597_);
  nand (_28659_, _28658_, _28656_);
  nand (_28660_, _28659_, _10602_);
  nor (_28661_, _28507_, _10146_);
  nor (_28663_, _10116_, _08783_);
  nor (_28664_, _28663_, _10602_);
  not (_28665_, _28664_);
  nor (_28666_, _28665_, _28661_);
  nor (_28667_, _28666_, _10616_);
  nand (_28668_, _28667_, _28660_);
  nor (_28669_, _28478_, _10612_);
  nor (_28670_, _28669_, _10615_);
  nand (_28671_, _28670_, _28668_);
  nor (_28672_, _28513_, _10614_);
  nor (_28674_, _28672_, _03866_);
  and (_28675_, _28674_, _28671_);
  or (_28676_, _28675_, _28472_);
  nand (_28677_, _28676_, _04706_);
  nor (_28678_, _10029_, _03477_);
  not (_28679_, _28678_);
  and (_28680_, _28513_, _03967_);
  nor (_28681_, _28680_, _28679_);
  nand (_28682_, _28681_, _28677_);
  nor (_28683_, _28507_, \oc8051_golden_model_1.PSW [7]);
  nor (_28685_, _10116_, _08059_);
  nor (_28686_, _28685_, _10030_);
  not (_28687_, _28686_);
  nor (_28688_, _28687_, _28683_);
  nor (_28689_, _28688_, _10628_);
  nand (_28690_, _28689_, _28682_);
  nor (_28691_, _28478_, _10027_);
  nor (_28692_, _28691_, _08528_);
  and (_28693_, _28692_, _28690_);
  nor (_28694_, _28513_, _08527_);
  or (_28696_, _28694_, _03835_);
  or (_28697_, _28696_, _28693_);
  and (_28698_, _10278_, _03835_);
  nor (_28699_, _28698_, _03954_);
  and (_28700_, _28699_, _28697_);
  and (_28701_, _10116_, _03954_);
  or (_28702_, _28701_, _28700_);
  nand (_28703_, _28702_, _28471_);
  nor (_28704_, _28507_, _08059_);
  nor (_28705_, _10116_, \oc8051_golden_model_1.PSW [7]);
  nor (_28707_, _28705_, _10015_);
  not (_28708_, _28707_);
  nor (_28709_, _28708_, _28704_);
  nor (_28710_, _28709_, _10646_);
  nand (_28711_, _28710_, _28703_);
  nor (_28712_, _28478_, _10012_);
  nor (_28713_, _28712_, _10011_);
  and (_28714_, _28713_, _28711_);
  nor (_28715_, _28513_, _10010_);
  or (_28716_, _28715_, _08006_);
  or (_28718_, _28716_, _28714_);
  and (_28719_, _28504_, _08006_);
  nor (_28720_, _28719_, _03974_);
  nand (_28721_, _28720_, _28718_);
  and (_28722_, _04608_, _03974_);
  nor (_28723_, _28722_, _03474_);
  nand (_28724_, _28723_, _28721_);
  nand (_28725_, _28724_, _04386_);
  and (_28726_, _28493_, _10860_);
  nor (_28727_, _10277_, _10860_);
  or (_28729_, _28727_, _04386_);
  or (_28730_, _28729_, _28726_);
  and (_28731_, _28730_, _10008_);
  nand (_28732_, _28731_, _28725_);
  nor (_28733_, _28478_, _10008_);
  nor (_28734_, _28733_, _09990_);
  and (_28735_, _28734_, _28732_);
  nor (_28736_, _28513_, _09989_);
  or (_28737_, _28736_, _07964_);
  or (_28738_, _28737_, _28735_);
  and (_28740_, _28504_, _07964_);
  nor (_28741_, _28740_, _03707_);
  nand (_28742_, _28741_, _28738_);
  and (_28743_, _04608_, _03707_);
  nor (_28744_, _28743_, _03394_);
  nand (_28745_, _28744_, _28742_);
  nand (_28746_, _28745_, _03706_);
  and (_28747_, _10278_, _10860_);
  nor (_28748_, _28481_, _10860_);
  nor (_28749_, _28748_, _28747_);
  and (_28751_, _28749_, _03705_);
  nor (_28752_, _28751_, _10888_);
  nand (_28753_, _28752_, _28746_);
  nor (_28754_, _28478_, _10887_);
  nor (_28755_, _28754_, _03703_);
  nand (_28756_, _28755_, _28753_);
  and (_28757_, _10116_, _03703_);
  nor (_28758_, _28757_, _27375_);
  nand (_28759_, _28758_, _28756_);
  nor (_28760_, _28478_, _10894_);
  nor (_28762_, _28760_, _03833_);
  and (_28763_, _28762_, _28759_);
  or (_28764_, _28763_, _28470_);
  nor (_28765_, _03400_, _03384_);
  nand (_28766_, _28765_, _28764_);
  and (_28767_, _28749_, _03384_);
  nor (_28768_, _28767_, _10911_);
  nand (_28769_, _28768_, _28766_);
  nor (_28770_, _28478_, _10910_);
  nor (_28771_, _28770_, _03701_);
  nand (_28773_, _28771_, _28769_);
  and (_28774_, _10116_, _03701_);
  nor (_28775_, _28774_, _26323_);
  nand (_28776_, _28775_, _28773_);
  nor (_28777_, _28478_, _10917_);
  nor (_28778_, _28777_, _03841_);
  and (_28779_, _28778_, _28776_);
  or (_28780_, _28779_, _28469_);
  nor (_28781_, _10928_, _03399_);
  and (_28782_, _28781_, _28780_);
  and (_28784_, _28478_, _10928_);
  or (_28785_, _28784_, _28782_);
  or (_28786_, _28785_, _42912_);
  or (_28787_, _42908_, \oc8051_golden_model_1.PC [8]);
  and (_28788_, _28787_, _41654_);
  and (_43277_, _28788_, _28786_);
  nor (_28789_, _09994_, \oc8051_golden_model_1.PC [9]);
  nor (_28790_, _28789_, _09995_);
  and (_28791_, _28790_, _10928_);
  nor (_28792_, _28790_, _10917_);
  nor (_28794_, _04482_, _06956_);
  nor (_28795_, _28790_, _10008_);
  nor (_28796_, _28790_, _10012_);
  and (_28797_, _10217_, _03835_);
  nor (_28798_, _28790_, _10027_);
  and (_28799_, _10217_, _03866_);
  nor (_28800_, _28790_, _10612_);
  and (_28801_, _10217_, _03838_);
  nor (_28802_, _28790_, _10585_);
  nor (_28803_, _10063_, _06305_);
  and (_28805_, _10063_, _03746_);
  nor (_28806_, _28790_, _10477_);
  and (_28807_, _10217_, _10181_);
  nor (_28808_, _10282_, _10279_);
  and (_28809_, _28808_, _10221_);
  nor (_28810_, _28808_, _10221_);
  nor (_28811_, _28810_, _28809_);
  nor (_28812_, _28811_, _10181_);
  nor (_28813_, _28812_, _28807_);
  nor (_28814_, _28813_, _03855_);
  and (_28816_, _10063_, _03690_);
  and (_28817_, _10063_, _03755_);
  not (_28818_, _28811_);
  and (_28819_, _28818_, _10316_);
  nor (_28820_, _25971_, _10218_);
  or (_28821_, _28820_, _04630_);
  or (_28822_, _28821_, _28819_);
  nor (_28823_, _10120_, _10117_);
  and (_28824_, _28823_, _10066_);
  nor (_28825_, _28823_, _10066_);
  nor (_28827_, _28825_, _28824_);
  nor (_28828_, _28827_, _10326_);
  and (_28829_, _10326_, _10063_);
  or (_28830_, _28829_, _28828_);
  nor (_28831_, _28830_, _06140_);
  and (_28832_, _10344_, _04944_);
  or (_28833_, _28832_, _28790_);
  not (_28834_, _10063_);
  and (_28835_, _28834_, _04615_);
  nor (_28836_, _28835_, _04234_);
  nor (_28838_, _04615_, \oc8051_golden_model_1.PC [9]);
  nand (_28839_, _28838_, _04944_);
  nand (_28840_, _28839_, _28836_);
  nand (_28841_, _28840_, _27451_);
  and (_28842_, _28841_, _28833_);
  and (_28843_, _28790_, _04234_);
  nor (_28844_, _28843_, _10320_);
  not (_28845_, _28844_);
  nor (_28846_, _28845_, _28842_);
  or (_28847_, _28846_, _04624_);
  nor (_28849_, _28847_, _28831_);
  and (_28850_, _28790_, _04624_);
  or (_28851_, _28850_, _03757_);
  or (_28852_, _28851_, _28849_);
  and (_28853_, _28852_, _28822_);
  nor (_28854_, _28853_, _10355_);
  nor (_28855_, _28790_, _10354_);
  nor (_28856_, _28855_, _03696_);
  not (_28857_, _28856_);
  nor (_28858_, _28857_, _28854_);
  and (_28859_, _10063_, _03696_);
  or (_28860_, _28859_, _04933_);
  nor (_28861_, _28860_, _28858_);
  nor (_28862_, _28861_, _03755_);
  or (_28863_, _28862_, _10365_);
  nor (_28864_, _28863_, _28817_);
  nor (_28865_, _28790_, _10364_);
  nor (_28866_, _28865_, _03750_);
  not (_28867_, _28866_);
  nor (_28868_, _28867_, _28864_);
  and (_28871_, _10063_, _03750_);
  nor (_28872_, _28871_, _10377_);
  not (_28873_, _28872_);
  nor (_28874_, _28873_, _28868_);
  nor (_28875_, _28790_, _10375_);
  nor (_28876_, _28875_, _03691_);
  not (_28877_, _28876_);
  nor (_28878_, _28877_, _28874_);
  and (_28879_, _10063_, _03691_);
  or (_28880_, _28879_, _10379_);
  or (_28882_, _28880_, _28878_);
  and (_28883_, _28882_, _04759_);
  or (_28884_, _28883_, _10425_);
  or (_28885_, _28884_, _28816_);
  and (_28886_, _10423_, _10217_);
  nor (_28887_, _28811_, _10423_);
  or (_28888_, _28887_, _28886_);
  nor (_28889_, _28888_, _10388_);
  nor (_28890_, _28889_, _03854_);
  and (_28891_, _28890_, _28885_);
  or (_28893_, _28891_, _28814_);
  nand (_28894_, _28893_, _10433_);
  and (_28895_, _10446_, _10217_);
  nor (_28896_, _28811_, _10446_);
  or (_28897_, _28896_, _28895_);
  and (_28898_, _28897_, _03847_);
  nor (_28899_, _28811_, _10462_);
  and (_28900_, _10462_, _10217_);
  nor (_28901_, _28900_, _28899_);
  nor (_28902_, _28901_, _04216_);
  nor (_28904_, _28902_, _28898_);
  and (_28905_, _28790_, _10431_);
  nor (_28906_, _28905_, _03684_);
  and (_28907_, _28906_, _28904_);
  nand (_28908_, _28907_, _28894_);
  and (_28909_, _28834_, _03684_);
  nor (_28910_, _28909_, _05105_);
  and (_28911_, _28910_, _26075_);
  nand (_28912_, _28911_, _28908_);
  nor (_28913_, _26075_, _28834_);
  nor (_28915_, _28913_, _10481_);
  and (_28916_, _28915_, _28912_);
  nor (_28917_, _28916_, _28806_);
  or (_28918_, _28917_, _03811_);
  and (_28919_, _28834_, _03811_);
  nor (_28920_, _28919_, _10483_);
  nand (_28921_, _28920_, _28918_);
  and (_28922_, _10063_, _03810_);
  nor (_28923_, _28922_, _10494_);
  and (_28924_, _28923_, _28921_);
  nor (_28926_, _28790_, _10488_);
  or (_28927_, _28926_, _28924_);
  nand (_28928_, _28927_, _10492_);
  nor (_28929_, _10063_, _10492_);
  nor (_28930_, _28929_, _03547_);
  nand (_28931_, _28930_, _28928_);
  and (_28932_, _28790_, _03547_);
  nor (_28933_, _28932_, _03679_);
  nand (_28934_, _28933_, _28931_);
  not (_28935_, _28600_);
  and (_28937_, _28834_, _03679_);
  nor (_28938_, _28937_, _28935_);
  nand (_28939_, _28938_, _28934_);
  and (_28940_, _10217_, _03861_);
  nor (_28941_, _28940_, _11528_);
  nand (_28942_, _28941_, _28939_);
  nor (_28943_, _10510_, _10063_);
  nor (_28944_, _28943_, _07559_);
  nand (_28945_, _28944_, _28942_);
  nor (_28946_, _10218_, _03415_);
  nor (_28948_, _28946_, _10521_);
  nand (_28949_, _28948_, _28945_);
  nor (_28950_, _28790_, _10517_);
  nor (_28951_, _28950_, _03746_);
  and (_28952_, _28951_, _28949_);
  or (_28953_, _28952_, _28805_);
  nand (_28954_, _28953_, _25812_);
  nor (_28955_, _28827_, _10526_);
  nor (_28956_, _28955_, _06306_);
  and (_28957_, _28956_, _28954_);
  or (_28959_, _28957_, _28803_);
  nand (_28960_, _28959_, _04694_);
  and (_28961_, _10218_, _03839_);
  nor (_28962_, _28961_, _08456_);
  nand (_28963_, _28962_, _28960_);
  and (_28964_, _10063_, _08456_);
  nor (_28965_, _28964_, _10540_);
  nand (_28966_, _28965_, _28963_);
  nor (_28967_, _10567_, \oc8051_golden_model_1.DPH [1]);
  nor (_28968_, _28967_, _10568_);
  nor (_28970_, _28968_, _10541_);
  nor (_28971_, _28970_, _03745_);
  nand (_28972_, _28971_, _28966_);
  and (_28973_, _10063_, _03745_);
  nor (_28974_, _28973_, _03483_);
  nand (_28975_, _28974_, _28972_);
  nand (_28976_, _28975_, _10580_);
  and (_28977_, _10063_, _08783_);
  nor (_28978_, _28827_, _08783_);
  or (_28979_, _28978_, _28977_);
  and (_28981_, _28979_, _10145_);
  nor (_28982_, _28981_, _10587_);
  and (_28983_, _28982_, _28976_);
  or (_28984_, _28983_, _28802_);
  nand (_28985_, _28984_, _10589_);
  nor (_28986_, _10589_, _10063_);
  nor (_28987_, _28986_, _03838_);
  and (_28988_, _28987_, _28985_);
  or (_28989_, _28988_, _28801_);
  nand (_28990_, _28989_, _04701_);
  and (_28992_, _10063_, _03959_);
  nor (_28993_, _28992_, _03486_);
  nand (_28994_, _28993_, _28990_);
  nand (_28995_, _28994_, _10602_);
  and (_28996_, _28827_, _08783_);
  nor (_28997_, _10063_, _08783_);
  nor (_28998_, _28997_, _10602_);
  not (_28999_, _28998_);
  nor (_29000_, _28999_, _28996_);
  nor (_29001_, _29000_, _10616_);
  and (_29003_, _29001_, _28995_);
  or (_29004_, _29003_, _28800_);
  nand (_29005_, _29004_, _10614_);
  nor (_29006_, _10063_, _10614_);
  nor (_29007_, _29006_, _03866_);
  and (_29008_, _29007_, _29005_);
  or (_29009_, _29008_, _28799_);
  nand (_29010_, _29009_, _04706_);
  and (_29011_, _10063_, _03967_);
  nor (_29012_, _29011_, _03477_);
  nand (_29014_, _29012_, _29010_);
  nand (_29015_, _29014_, _10030_);
  and (_29016_, _28827_, _08059_);
  nor (_29017_, _10063_, _08059_);
  nor (_29018_, _29017_, _10030_);
  not (_29019_, _29018_);
  nor (_29020_, _29019_, _29016_);
  nor (_29021_, _29020_, _10628_);
  and (_29022_, _29021_, _29015_);
  or (_29023_, _29022_, _28798_);
  nand (_29025_, _29023_, _08527_);
  nor (_29026_, _10063_, _08527_);
  nor (_29027_, _29026_, _03835_);
  and (_29028_, _29027_, _29025_);
  or (_29029_, _29028_, _28797_);
  nand (_29030_, _29029_, _06537_);
  and (_29031_, _10063_, _03954_);
  nor (_29032_, _29031_, _03481_);
  nand (_29033_, _29032_, _29030_);
  nand (_29034_, _29033_, _10015_);
  and (_29036_, _28827_, \oc8051_golden_model_1.PSW [7]);
  nor (_29037_, _10063_, \oc8051_golden_model_1.PSW [7]);
  nor (_29038_, _29037_, _10015_);
  not (_29039_, _29038_);
  nor (_29040_, _29039_, _29036_);
  nor (_29041_, _29040_, _10646_);
  and (_29042_, _29041_, _29034_);
  or (_29043_, _29042_, _28796_);
  nand (_29044_, _29043_, _10010_);
  nor (_29045_, _10063_, _10010_);
  nor (_29047_, _29045_, _08006_);
  nand (_29048_, _29047_, _29044_);
  and (_29049_, _28790_, _08006_);
  nor (_29050_, _29049_, _03974_);
  nand (_29051_, _29050_, _29048_);
  nor (_29052_, _03831_, _03474_);
  not (_29053_, _29052_);
  and (_29054_, _04842_, _03974_);
  nor (_29055_, _29054_, _29053_);
  nand (_29056_, _29055_, _29051_);
  nor (_29058_, _10217_, _10860_);
  and (_29059_, _28811_, _10860_);
  or (_29060_, _29059_, _04386_);
  or (_29061_, _29060_, _29058_);
  and (_29062_, _29061_, _10008_);
  and (_29063_, _29062_, _29056_);
  or (_29064_, _29063_, _28795_);
  nand (_29065_, _29064_, _09989_);
  nor (_29066_, _10063_, _09989_);
  nor (_29067_, _29066_, _07964_);
  nand (_29069_, _29067_, _29065_);
  and (_29070_, _28790_, _07964_);
  nor (_29071_, _29070_, _03707_);
  nand (_29072_, _29071_, _29069_);
  and (_29073_, _04842_, _03707_);
  nor (_29074_, _03705_, _03394_);
  not (_29075_, _29074_);
  nor (_29076_, _29075_, _29073_);
  nand (_29077_, _29076_, _29072_);
  nor (_29078_, _28818_, _10860_);
  and (_29080_, _10218_, _10860_);
  nor (_29081_, _29080_, _29078_);
  and (_29082_, _29081_, _03705_);
  nor (_29083_, _29082_, _10888_);
  nand (_29084_, _29083_, _29077_);
  nor (_29085_, _28790_, _10887_);
  nor (_29086_, _29085_, _03703_);
  nand (_29087_, _29086_, _29084_);
  and (_29088_, _10063_, _03703_);
  nor (_29089_, _29088_, _27375_);
  nand (_29091_, _29089_, _29087_);
  nor (_29092_, _28790_, _10894_);
  nor (_29093_, _29092_, _03833_);
  and (_29094_, _29093_, _29091_);
  or (_29095_, _29094_, _28794_);
  nand (_29096_, _29095_, _28765_);
  and (_29097_, _29081_, _03384_);
  nor (_29098_, _29097_, _10911_);
  nand (_29099_, _29098_, _29096_);
  nor (_29100_, _28790_, _10910_);
  nor (_29102_, _29100_, _03701_);
  nand (_29103_, _29102_, _29099_);
  and (_29104_, _10063_, _03701_);
  nor (_29105_, _29104_, _26323_);
  and (_29106_, _29105_, _29103_);
  or (_29107_, _29106_, _28792_);
  nand (_29108_, _29107_, _10921_);
  not (_29109_, _28781_);
  and (_29110_, _04482_, _03841_);
  nor (_29111_, _29110_, _29109_);
  and (_29113_, _29111_, _29108_);
  or (_29114_, _29113_, _28791_);
  or (_29115_, _29114_, _42912_);
  or (_29116_, _42908_, \oc8051_golden_model_1.PC [9]);
  and (_29117_, _29116_, _41654_);
  and (_43278_, _29117_, _29115_);
  and (_29118_, _04165_, _03833_);
  nor (_29119_, _09995_, \oc8051_golden_model_1.PC [10]);
  nor (_29120_, _29119_, _09996_);
  nor (_29121_, _29120_, _10887_);
  not (_29123_, _29120_);
  and (_29124_, _29123_, _07964_);
  and (_29125_, _29123_, _08006_);
  and (_29126_, _10211_, _03835_);
  and (_29127_, _10211_, _03866_);
  and (_29128_, _10211_, _03838_);
  or (_29129_, _10145_, _03483_);
  nor (_29130_, _29120_, _10488_);
  not (_29131_, _10051_);
  and (_29132_, _29131_, _03810_);
  and (_29134_, _29120_, _10431_);
  and (_29135_, _10446_, _10210_);
  not (_29136_, _10214_);
  nor (_29137_, _10286_, _10283_);
  nor (_29138_, _29137_, _29136_);
  and (_29139_, _29137_, _29136_);
  nor (_29140_, _29139_, _29138_);
  and (_29141_, _29140_, _27160_);
  or (_29142_, _29141_, _29135_);
  and (_29143_, _29142_, _03847_);
  nand (_29145_, _10462_, _10211_);
  or (_29146_, _29140_, _10462_);
  and (_29147_, _29146_, _03773_);
  and (_29148_, _29147_, _29145_);
  or (_29149_, _29148_, _29143_);
  or (_29150_, _29149_, _29134_);
  nand (_29151_, _10211_, _10181_);
  or (_29152_, _29140_, _10181_);
  and (_29153_, _29152_, _03854_);
  and (_29154_, _29153_, _29151_);
  or (_29156_, _29120_, _10364_);
  nand (_29157_, _29131_, _04109_);
  nor (_29158_, _04615_, \oc8051_golden_model_1.PC [10]);
  nand (_29159_, _29158_, _04944_);
  and (_29160_, _29159_, _29157_);
  or (_29161_, _29160_, _04234_);
  or (_29162_, _29120_, _28144_);
  and (_29163_, _29162_, _29161_);
  nor (_29164_, _29123_, _10344_);
  nand (_29165_, _06140_, _04948_);
  or (_29167_, _29165_, _29164_);
  or (_29168_, _29167_, _29163_);
  not (_29169_, _10060_);
  nor (_29170_, _10124_, _10121_);
  nor (_29171_, _29170_, _29169_);
  and (_29172_, _29170_, _29169_);
  nor (_29173_, _29172_, _29171_);
  and (_29174_, _29173_, _10324_);
  and (_29175_, _10326_, _10051_);
  or (_29176_, _29175_, _29174_);
  or (_29178_, _29176_, _06140_);
  and (_29179_, _29178_, _29168_);
  or (_29180_, _29179_, _04624_);
  nand (_29181_, _29123_, _04624_);
  and (_29182_, _29181_, _04630_);
  and (_29183_, _29182_, _29180_);
  and (_29184_, _10314_, _10210_);
  and (_29185_, _29140_, _10316_);
  or (_29186_, _29185_, _29184_);
  and (_29187_, _29186_, _03757_);
  or (_29189_, _29187_, _29183_);
  or (_29190_, _29189_, _10355_);
  or (_29191_, _29120_, _10354_);
  and (_29192_, _29191_, _03697_);
  and (_29193_, _29192_, _29190_);
  or (_29194_, _29193_, _04933_);
  and (_29195_, _29194_, _04537_);
  nor (_29196_, _29131_, _03761_);
  or (_29197_, _29196_, _10365_);
  or (_29198_, _29197_, _29195_);
  and (_29200_, _29198_, _29156_);
  or (_29201_, _29200_, _03750_);
  nand (_29202_, _29131_, _03750_);
  and (_29203_, _29202_, _10375_);
  and (_29204_, _29203_, _29201_);
  nor (_29205_, _29123_, _10375_);
  or (_29206_, _29205_, _29204_);
  and (_29207_, _29206_, _03692_);
  and (_29208_, _10051_, _03691_);
  or (_29209_, _29208_, _10379_);
  or (_29211_, _29209_, _29207_);
  and (_29212_, _29211_, _04759_);
  or (_29213_, _29140_, _10423_);
  nand (_29214_, _10423_, _10211_);
  and (_29215_, _29214_, _29213_);
  and (_29216_, _29215_, _10386_);
  and (_29217_, _10051_, _03690_);
  or (_29218_, _29217_, _10387_);
  or (_29219_, _29218_, _29216_);
  or (_29220_, _29219_, _29212_);
  or (_29221_, _29215_, _10388_);
  and (_29222_, _29221_, _03855_);
  and (_29223_, _29222_, _29220_);
  or (_29224_, _29223_, _29154_);
  and (_29225_, _29224_, _10433_);
  nor (_29226_, _29225_, _29150_);
  and (_29227_, _26075_, _03685_);
  not (_29228_, _29227_);
  or (_29229_, _29228_, _29226_);
  nor (_29230_, _29227_, _29131_);
  nand (_29232_, _10477_, _03442_);
  nor (_29233_, _29232_, _29230_);
  and (_29234_, _29233_, _29229_);
  nor (_29235_, _29120_, _10477_);
  nor (_29236_, _29235_, _03811_);
  not (_29237_, _29236_);
  nor (_29238_, _29237_, _29234_);
  and (_29239_, _10051_, _03811_);
  or (_29240_, _29239_, _10483_);
  nor (_29241_, _29240_, _29238_);
  nor (_29243_, _29241_, _29132_);
  nor (_29244_, _29243_, _10494_);
  or (_29245_, _29244_, _10493_);
  or (_29246_, _29245_, _29130_);
  nor (_29247_, _29131_, _10492_);
  nor (_29248_, _29247_, _03547_);
  nand (_29249_, _29248_, _29246_);
  nor (_29250_, _29120_, _03422_);
  nor (_29251_, _29250_, _03679_);
  and (_29252_, _29251_, _29249_);
  and (_29254_, _10051_, _03679_);
  nor (_29255_, _29254_, _29252_);
  and (_29256_, _29255_, _28600_);
  and (_29257_, _10211_, _03861_);
  or (_29258_, _29257_, _29256_);
  and (_29259_, _29258_, _10510_);
  nor (_29260_, _10510_, _10051_);
  or (_29261_, _29260_, _29259_);
  nand (_29262_, _29261_, _03415_);
  nor (_29263_, _10210_, _03415_);
  nor (_29265_, _29263_, _10521_);
  and (_29266_, _29265_, _29262_);
  nor (_29267_, _29123_, _10517_);
  or (_29268_, _29267_, _29266_);
  nand (_29269_, _29268_, _27577_);
  and (_29270_, _10051_, _03746_);
  nor (_29271_, _29270_, _25813_);
  nand (_29272_, _29271_, _29269_);
  nor (_29273_, _29173_, _10526_);
  nor (_29274_, _29273_, _06306_);
  and (_29276_, _29274_, _29272_);
  nor (_29277_, _29131_, _06305_);
  or (_29278_, _29277_, _03839_);
  or (_29279_, _29278_, _29276_);
  and (_29280_, _10211_, _03839_);
  nor (_29281_, _29280_, _08456_);
  nand (_29282_, _29281_, _29279_);
  and (_29283_, _10051_, _08456_);
  nor (_29284_, _29283_, _10540_);
  nand (_29285_, _29284_, _29282_);
  nor (_29287_, _10568_, \oc8051_golden_model_1.DPH [2]);
  nor (_29288_, _29287_, _10569_);
  nor (_29289_, _29288_, _10541_);
  nor (_29290_, _29289_, _03745_);
  and (_29291_, _29290_, _29285_);
  and (_29292_, _10051_, _03745_);
  nor (_29293_, _29292_, _29291_);
  or (_29294_, _29293_, _29129_);
  and (_29295_, _10051_, _08783_);
  and (_29296_, _29173_, _10146_);
  or (_29298_, _29296_, _29295_);
  and (_29299_, _29298_, _10145_);
  nor (_29300_, _29299_, _10587_);
  nand (_29301_, _29300_, _29294_);
  nor (_29302_, _29120_, _10585_);
  nor (_29303_, _29302_, _10590_);
  nand (_29304_, _29303_, _29301_);
  nor (_29305_, _10589_, _29131_);
  nor (_29306_, _29305_, _03838_);
  and (_29307_, _29306_, _29304_);
  or (_29309_, _29307_, _29128_);
  nand (_29310_, _29309_, _04701_);
  and (_29311_, _29131_, _03959_);
  nor (_29312_, _10601_, _03486_);
  not (_29313_, _29312_);
  nor (_29314_, _29313_, _29311_);
  nand (_29315_, _29314_, _29310_);
  nor (_29316_, _29173_, _10146_);
  nor (_29317_, _10051_, _08783_);
  nor (_29318_, _29317_, _10602_);
  not (_29320_, _29318_);
  nor (_29321_, _29320_, _29316_);
  nor (_29322_, _29321_, _10616_);
  nand (_29323_, _29322_, _29315_);
  nor (_29324_, _29120_, _10612_);
  nor (_29325_, _29324_, _10615_);
  nand (_29326_, _29325_, _29323_);
  nor (_29327_, _29131_, _10614_);
  nor (_29328_, _29327_, _03866_);
  and (_29329_, _29328_, _29326_);
  or (_29331_, _29329_, _29127_);
  nand (_29332_, _29331_, _04706_);
  and (_29333_, _29131_, _03967_);
  nor (_29334_, _29333_, _28679_);
  nand (_29335_, _29334_, _29332_);
  nor (_29336_, _29173_, \oc8051_golden_model_1.PSW [7]);
  nor (_29337_, _10051_, _08059_);
  nor (_29338_, _29337_, _10030_);
  not (_29339_, _29338_);
  nor (_29340_, _29339_, _29336_);
  nor (_29342_, _29340_, _10628_);
  nand (_29343_, _29342_, _29335_);
  nor (_29344_, _29120_, _10027_);
  nor (_29345_, _29344_, _08528_);
  nand (_29346_, _29345_, _29343_);
  nor (_29347_, _29131_, _08527_);
  nor (_29348_, _29347_, _03835_);
  and (_29349_, _29348_, _29346_);
  or (_29350_, _29349_, _29126_);
  nand (_29351_, _29350_, _06537_);
  and (_29353_, _29131_, _03954_);
  not (_29354_, _29353_);
  and (_29355_, _29354_, _28471_);
  nand (_29356_, _29355_, _29351_);
  nand (_29357_, _10051_, _08059_);
  nand (_29358_, _29173_, \oc8051_golden_model_1.PSW [7]);
  and (_29359_, _29358_, _29357_);
  or (_29360_, _29359_, _10015_);
  and (_29361_, _29360_, _29356_);
  nand (_29362_, _29361_, _10012_);
  nor (_29364_, _29120_, _10012_);
  nor (_29365_, _29364_, _10011_);
  nand (_29366_, _29365_, _29362_);
  nor (_29367_, _29131_, _10010_);
  nor (_29368_, _29367_, _08006_);
  and (_29369_, _29368_, _29366_);
  or (_29370_, _29369_, _29125_);
  nand (_29371_, _29370_, _11621_);
  and (_29372_, _05236_, _03974_);
  nor (_29373_, _29372_, _29053_);
  nand (_29375_, _29373_, _29371_);
  nor (_29376_, _10211_, _10860_);
  and (_29377_, _29140_, _10860_);
  or (_29378_, _29377_, _29376_);
  and (_29379_, _29378_, _03831_);
  nor (_29380_, _29379_, _10669_);
  nand (_29381_, _29380_, _29375_);
  nor (_29382_, _29120_, _10008_);
  nor (_29383_, _29382_, _09990_);
  nand (_29384_, _29383_, _29381_);
  nor (_29386_, _29131_, _09989_);
  nor (_29387_, _29386_, _07964_);
  and (_29388_, _29387_, _29384_);
  or (_29389_, _29388_, _29124_);
  nand (_29390_, _29389_, _03708_);
  and (_29391_, _05236_, _03707_);
  nor (_29392_, _29391_, _29075_);
  nand (_29393_, _29392_, _29390_);
  nor (_29394_, _29140_, _10860_);
  and (_29395_, _10211_, _10860_);
  nor (_29397_, _29395_, _29394_);
  and (_29398_, _29397_, _03705_);
  nor (_29399_, _29398_, _10888_);
  and (_29400_, _29399_, _29393_);
  or (_29401_, _29400_, _29121_);
  nand (_29402_, _29401_, _03704_);
  and (_29403_, _29131_, _03703_);
  nor (_29404_, _29403_, _27375_);
  nand (_29405_, _29404_, _29402_);
  nor (_29406_, _29123_, _10894_);
  nor (_29407_, _29406_, _03833_);
  nand (_29408_, _29407_, _29405_);
  nand (_29409_, _29408_, _28765_);
  or (_29410_, _29409_, _29118_);
  and (_29411_, _29397_, _03384_);
  nor (_29412_, _29411_, _10911_);
  and (_29413_, _29412_, _29410_);
  nor (_29414_, _29120_, _10910_);
  or (_29415_, _29414_, _29413_);
  nand (_29416_, _29415_, _03702_);
  and (_29419_, _29131_, _03701_);
  nor (_29420_, _29419_, _26323_);
  nand (_29421_, _29420_, _29416_);
  nor (_29422_, _29123_, _10917_);
  nor (_29423_, _29422_, _03841_);
  nand (_29424_, _29423_, _29421_);
  and (_29425_, _04165_, _03841_);
  nor (_29426_, _29425_, _29109_);
  and (_29427_, _29426_, _29424_);
  and (_29428_, _29120_, _10928_);
  or (_29430_, _29428_, _29427_);
  or (_29431_, _29430_, _42912_);
  or (_29432_, _42908_, \oc8051_golden_model_1.PC [10]);
  and (_29433_, _29432_, _41654_);
  and (_43279_, _29433_, _29431_);
  nor (_29434_, _09996_, \oc8051_golden_model_1.PC [11]);
  nor (_29435_, _29434_, _09997_);
  and (_29436_, _29435_, _10928_);
  or (_29437_, _29435_, _10008_);
  or (_29438_, _29435_, _10012_);
  or (_29440_, _10055_, _10016_);
  and (_29441_, _29440_, _10015_);
  or (_29442_, _29435_, _10027_);
  or (_29443_, _10055_, _10031_);
  and (_29444_, _29443_, _10030_);
  or (_29445_, _29435_, _10585_);
  nor (_29446_, _10205_, _03415_);
  nor (_29447_, _29138_, _10212_);
  and (_29448_, _29447_, _10208_);
  nor (_29449_, _29447_, _10208_);
  or (_29451_, _29449_, _29448_);
  or (_29452_, _29451_, _10446_);
  nand (_29453_, _10446_, _10205_);
  and (_29454_, _29453_, _03847_);
  and (_29455_, _29454_, _29452_);
  nand (_29456_, _10205_, _10181_);
  or (_29457_, _29451_, _10181_);
  and (_29458_, _29457_, _03854_);
  and (_29459_, _29458_, _29456_);
  nand (_29460_, _10423_, _10205_);
  or (_29462_, _29451_, _10423_);
  and (_29463_, _29462_, _10425_);
  and (_29464_, _29463_, _29460_);
  and (_29465_, _10055_, _03750_);
  and (_29466_, _10314_, _10204_);
  and (_29467_, _29451_, _10316_);
  or (_29468_, _29467_, _29466_);
  and (_29469_, _29468_, _03757_);
  nor (_29470_, _29171_, _10052_);
  nor (_29471_, _29470_, _10058_);
  and (_29473_, _29470_, _10058_);
  or (_29474_, _29473_, _29471_);
  and (_29475_, _29474_, _10324_);
  and (_29476_, _10326_, _10055_);
  or (_29477_, _29476_, _29475_);
  and (_29478_, _29477_, _10320_);
  or (_29479_, _29435_, _28144_);
  or (_29480_, _10055_, _10331_);
  nor (_29481_, _04615_, \oc8051_golden_model_1.PC [11]);
  nand (_29482_, _29481_, _04944_);
  and (_29484_, _29482_, _29480_);
  or (_29485_, _29484_, _04234_);
  and (_29486_, _29485_, _04948_);
  and (_29487_, _29486_, _29479_);
  and (_29488_, _10055_, _04111_);
  and (_29489_, _29435_, _25715_);
  or (_29490_, _29489_, _29488_);
  or (_29491_, _29490_, _29487_);
  and (_29492_, _29491_, _06140_);
  or (_29493_, _29492_, _04624_);
  or (_29495_, _29493_, _29478_);
  and (_29496_, _29495_, _04630_);
  or (_29497_, _29496_, _10355_);
  or (_29498_, _29497_, _29469_);
  or (_29499_, _29435_, _10360_);
  and (_29500_, _29499_, _10359_);
  and (_29501_, _29500_, _29498_);
  and (_29502_, _10366_, _10055_);
  or (_29503_, _29502_, _10365_);
  or (_29504_, _29503_, _29501_);
  or (_29506_, _29435_, _10364_);
  and (_29507_, _29506_, _03751_);
  and (_29508_, _29507_, _29504_);
  or (_29509_, _29508_, _29465_);
  and (_29510_, _29509_, _10375_);
  and (_29511_, _29435_, _10377_);
  or (_29512_, _29511_, _10382_);
  or (_29513_, _29512_, _29510_);
  or (_29514_, _10381_, _10055_);
  and (_29515_, _29514_, _10388_);
  and (_29517_, _29515_, _29513_);
  or (_29518_, _29517_, _29464_);
  and (_29519_, _29518_, _03855_);
  or (_29520_, _29519_, _03773_);
  or (_29521_, _29520_, _29459_);
  and (_29522_, _10462_, _10204_);
  not (_29523_, _10462_);
  and (_29524_, _29451_, _29523_);
  or (_29525_, _29524_, _04216_);
  or (_29526_, _29525_, _29522_);
  and (_29528_, _29526_, _11721_);
  and (_29529_, _29528_, _29521_);
  or (_29530_, _29529_, _29455_);
  and (_29531_, _29530_, _10432_);
  nand (_29532_, _29435_, _10431_);
  nand (_29533_, _29532_, _10470_);
  or (_29534_, _29533_, _29531_);
  or (_29535_, _10470_, _10055_);
  and (_29536_, _29535_, _10477_);
  and (_29537_, _29536_, _29534_);
  and (_29539_, _29435_, _10481_);
  or (_29540_, _29539_, _10485_);
  or (_29541_, _29540_, _29537_);
  or (_29542_, _10484_, _10055_);
  and (_29543_, _29542_, _10488_);
  and (_29544_, _29543_, _29541_);
  and (_29545_, _29435_, _10494_);
  or (_29546_, _29545_, _10493_);
  or (_29547_, _29546_, _29544_);
  or (_29548_, _10055_, _10492_);
  and (_29550_, _29548_, _03422_);
  and (_29551_, _29550_, _29547_);
  nand (_29552_, _29435_, _03547_);
  nand (_29553_, _29552_, _10502_);
  or (_29554_, _29553_, _29551_);
  or (_29555_, _10502_, _10055_);
  and (_29556_, _29555_, _09806_);
  and (_29557_, _29556_, _29554_);
  nand (_29558_, _10204_, _03861_);
  nand (_29559_, _29558_, _10510_);
  or (_29561_, _29559_, _29557_);
  or (_29562_, _10510_, _10055_);
  and (_29563_, _29562_, _03415_);
  and (_29564_, _29563_, _29561_);
  or (_29565_, _29564_, _29446_);
  and (_29566_, _29565_, _10517_);
  and (_29567_, _29435_, _10521_);
  or (_29568_, _29567_, _10520_);
  or (_29569_, _29568_, _29566_);
  or (_29570_, _10519_, _10055_);
  and (_29572_, _29570_, _10526_);
  and (_29573_, _29572_, _29569_);
  and (_29574_, _29474_, _10525_);
  or (_29575_, _29574_, _06306_);
  or (_29576_, _29575_, _29573_);
  or (_29577_, _10055_, _06305_);
  and (_29578_, _29577_, _04694_);
  and (_29579_, _29578_, _29576_);
  and (_29580_, _10204_, _03839_);
  or (_29581_, _29580_, _08456_);
  or (_29583_, _29581_, _29579_);
  or (_29584_, _10055_, _08457_);
  and (_29585_, _29584_, _10541_);
  and (_29586_, _29585_, _29583_);
  or (_29587_, _10569_, \oc8051_golden_model_1.DPH [3]);
  nor (_29588_, _10570_, _10541_);
  and (_29589_, _29588_, _29587_);
  or (_29590_, _29589_, _10544_);
  or (_29591_, _29590_, _29586_);
  or (_29592_, _10543_, _10055_);
  and (_29594_, _29592_, _10580_);
  and (_29595_, _29594_, _29591_);
  or (_29596_, _29474_, _08783_);
  or (_29597_, _10055_, _10146_);
  and (_29598_, _29597_, _10145_);
  and (_29599_, _29598_, _29596_);
  or (_29600_, _29599_, _10587_);
  or (_29601_, _29600_, _29595_);
  and (_29602_, _29601_, _29445_);
  or (_29603_, _29602_, _10590_);
  or (_29605_, _10589_, _10055_);
  and (_29606_, _29605_, _04703_);
  and (_29607_, _29606_, _29603_);
  nand (_29608_, _10204_, _03838_);
  nand (_29609_, _29608_, _10597_);
  or (_29610_, _29609_, _29607_);
  or (_29611_, _10597_, _10055_);
  and (_29612_, _29611_, _10602_);
  and (_29613_, _29612_, _29610_);
  or (_29614_, _29474_, _10146_);
  or (_29616_, _10055_, _08783_);
  and (_29617_, _29616_, _10601_);
  and (_29618_, _29617_, _29614_);
  or (_29619_, _29618_, _29613_);
  and (_29620_, _29619_, _10612_);
  and (_29621_, _29435_, _10616_);
  or (_29622_, _29621_, _10615_);
  or (_29623_, _29622_, _29620_);
  or (_29624_, _10055_, _10614_);
  and (_29625_, _29624_, _04708_);
  and (_29627_, _29625_, _29623_);
  nand (_29628_, _10204_, _03866_);
  nand (_29629_, _29628_, _10031_);
  or (_29630_, _29629_, _29627_);
  and (_29631_, _29630_, _29444_);
  or (_29632_, _29474_, \oc8051_golden_model_1.PSW [7]);
  or (_29633_, _10055_, _08059_);
  and (_29634_, _29633_, _10029_);
  and (_29635_, _29634_, _29632_);
  or (_29636_, _29635_, _10628_);
  or (_29638_, _29636_, _29631_);
  and (_29639_, _29638_, _29442_);
  or (_29640_, _29639_, _08528_);
  or (_29641_, _10055_, _08527_);
  and (_29642_, _29641_, _06532_);
  and (_29643_, _29642_, _29640_);
  nand (_29644_, _10204_, _03835_);
  nand (_29645_, _29644_, _10016_);
  or (_29646_, _29645_, _29643_);
  and (_29647_, _29646_, _29441_);
  or (_29649_, _29474_, _08059_);
  or (_29650_, _10055_, \oc8051_golden_model_1.PSW [7]);
  and (_29651_, _29650_, _10014_);
  and (_29652_, _29651_, _29649_);
  or (_29653_, _29652_, _10646_);
  or (_29654_, _29653_, _29647_);
  and (_29655_, _29654_, _29438_);
  or (_29656_, _29655_, _10011_);
  or (_29657_, _10055_, _10010_);
  and (_29658_, _29657_, _08007_);
  and (_29660_, _29658_, _29656_);
  and (_29661_, _29435_, _08006_);
  or (_29662_, _29661_, _03974_);
  or (_29663_, _29662_, _29660_);
  nand (_29664_, _05050_, _03974_);
  and (_29665_, _29664_, _29663_);
  or (_29666_, _29665_, _03474_);
  or (_29667_, _10055_, _06543_);
  and (_29668_, _29667_, _04386_);
  and (_29669_, _29668_, _29666_);
  or (_29670_, _29451_, _10861_);
  or (_29671_, _10204_, _10860_);
  and (_29672_, _29671_, _03831_);
  and (_29673_, _29672_, _29670_);
  or (_29674_, _29673_, _10669_);
  or (_29675_, _29674_, _29669_);
  and (_29676_, _29675_, _29437_);
  or (_29677_, _29676_, _09990_);
  or (_29678_, _10055_, _09989_);
  and (_29679_, _29678_, _10870_);
  and (_29682_, _29679_, _29677_);
  and (_29683_, _29435_, _07964_);
  or (_29684_, _29683_, _03707_);
  or (_29685_, _29684_, _29682_);
  nand (_29686_, _05050_, _03707_);
  and (_29687_, _29686_, _29685_);
  or (_29688_, _29687_, _03394_);
  or (_29689_, _10055_, _03395_);
  and (_29690_, _29689_, _03706_);
  and (_29691_, _29690_, _29688_);
  or (_29693_, _29451_, _10860_);
  nand (_29694_, _10205_, _10860_);
  and (_29695_, _29694_, _29693_);
  and (_29696_, _29695_, _03705_);
  or (_29697_, _29696_, _10888_);
  or (_29698_, _29697_, _29691_);
  or (_29699_, _29435_, _10887_);
  and (_29700_, _29699_, _03704_);
  and (_29701_, _29700_, _29698_);
  nand (_29702_, _10055_, _03703_);
  nand (_29704_, _29702_, _10894_);
  or (_29705_, _29704_, _29701_);
  or (_29706_, _29435_, _10894_);
  and (_29707_, _29706_, _06956_);
  and (_29708_, _29707_, _29705_);
  nor (_29709_, _06956_, _03669_);
  or (_29710_, _29709_, _03400_);
  or (_29711_, _29710_, _29708_);
  or (_29712_, _10055_, _10904_);
  and (_29713_, _29712_, _03385_);
  and (_29715_, _29713_, _29711_);
  and (_29716_, _29695_, _03384_);
  or (_29717_, _29716_, _10911_);
  or (_29718_, _29717_, _29715_);
  or (_29719_, _29435_, _10910_);
  and (_29720_, _29719_, _03702_);
  and (_29721_, _29720_, _29718_);
  nand (_29722_, _10055_, _03701_);
  nand (_29723_, _29722_, _10917_);
  or (_29724_, _29723_, _29721_);
  or (_29726_, _29435_, _10917_);
  and (_29727_, _29726_, _10921_);
  and (_29728_, _29727_, _29724_);
  nor (_29729_, _10921_, _03669_);
  or (_29730_, _29729_, _03399_);
  or (_29731_, _29730_, _29728_);
  or (_29732_, _10055_, _10930_);
  and (_29733_, _29732_, _10929_);
  and (_29734_, _29733_, _29731_);
  or (_29735_, _29734_, _29436_);
  or (_29737_, _29735_, _42912_);
  or (_29738_, _42908_, \oc8051_golden_model_1.PC [11]);
  and (_29739_, _29738_, _41654_);
  and (_43282_, _29739_, _29737_);
  nor (_29740_, _09997_, \oc8051_golden_model_1.PC [12]);
  nor (_29741_, _29740_, _09998_);
  not (_29742_, _29741_);
  and (_29743_, _29742_, _10928_);
  and (_29744_, _04446_, _03841_);
  or (_29745_, _29744_, _03399_);
  and (_29747_, _29742_, _07964_);
  not (_29748_, _10048_);
  nor (_29749_, _29748_, _10016_);
  nor (_29750_, _29748_, _10031_);
  nor (_29751_, _10597_, _29748_);
  nor (_29752_, _10543_, _29748_);
  nor (_29753_, _10048_, _10492_);
  nor (_29754_, _29741_, _10477_);
  nor (_29755_, _29741_, _10364_);
  and (_29756_, _10131_, _10128_);
  nor (_29758_, _29756_, _10132_);
  and (_29759_, _29758_, _10324_);
  and (_29760_, _10326_, _10048_);
  or (_29761_, _29760_, _29759_);
  nor (_29762_, _29761_, _06140_);
  and (_29763_, _29748_, _04111_);
  or (_29764_, _29763_, _25715_);
  or (_29765_, _29741_, _25708_);
  nand (_29766_, _29748_, _04109_);
  nor (_29767_, _04615_, \oc8051_golden_model_1.PC [12]);
  nand (_29768_, _29767_, _04944_);
  and (_29769_, _29768_, _29766_);
  or (_29770_, _29769_, _04234_);
  and (_29771_, _29770_, _29765_);
  nor (_29772_, _29771_, _04111_);
  nor (_29773_, _29772_, _29764_);
  nor (_29774_, _29742_, _10344_);
  nor (_29775_, _29774_, _10320_);
  not (_29776_, _29775_);
  nor (_29777_, _29776_, _29773_);
  nor (_29779_, _29777_, _29762_);
  nor (_29780_, _29779_, _04624_);
  and (_29781_, _29742_, _04624_);
  nor (_29782_, _29781_, _03757_);
  not (_29783_, _29782_);
  nor (_29784_, _29783_, _29780_);
  and (_29785_, _10314_, _10200_);
  and (_29786_, _10293_, _10290_);
  nor (_29787_, _29786_, _10294_);
  and (_29788_, _29787_, _10316_);
  or (_29790_, _29788_, _29785_);
  and (_29791_, _29790_, _03757_);
  nor (_29792_, _29791_, _29784_);
  and (_29793_, _29792_, _10354_);
  nor (_29794_, _29741_, _10354_);
  nor (_29795_, _29794_, _10366_);
  not (_29796_, _29795_);
  or (_29797_, _29796_, _29793_);
  nor (_29798_, _10359_, _29748_);
  nor (_29799_, _29798_, _10365_);
  and (_29801_, _29799_, _29797_);
  or (_29802_, _29801_, _29755_);
  nand (_29803_, _29802_, _03751_);
  and (_29804_, _29748_, _03750_);
  nor (_29805_, _29804_, _10377_);
  and (_29806_, _29805_, _29803_);
  nor (_29807_, _29742_, _10375_);
  or (_29808_, _29807_, _29806_);
  nand (_29809_, _29808_, _10381_);
  nor (_29810_, _10381_, _29748_);
  nor (_29812_, _29810_, _10425_);
  and (_29813_, _29812_, _29809_);
  and (_29814_, _10423_, _10200_);
  not (_29815_, _29787_);
  nor (_29816_, _29815_, _10423_);
  or (_29817_, _29816_, _29814_);
  nor (_29818_, _29817_, _10388_);
  or (_29819_, _29818_, _29813_);
  nand (_29820_, _29819_, _03855_);
  and (_29821_, _10200_, _10181_);
  nor (_29823_, _29815_, _10181_);
  or (_29824_, _29823_, _29821_);
  nor (_29825_, _29824_, _03855_);
  nor (_29826_, _29825_, _03773_);
  nand (_29827_, _29826_, _29820_);
  and (_29828_, _10462_, _10201_);
  nor (_29829_, _29787_, _10462_);
  or (_29830_, _29829_, _04216_);
  or (_29831_, _29830_, _29828_);
  nand (_29832_, _29831_, _29827_);
  nand (_29834_, _29832_, _11721_);
  and (_29835_, _10446_, _10200_);
  and (_29836_, _29787_, _27160_);
  or (_29837_, _29836_, _29835_);
  and (_29838_, _29837_, _03847_);
  nor (_29839_, _29838_, _10431_);
  nand (_29840_, _29839_, _29834_);
  and (_29841_, _29742_, _10431_);
  not (_29842_, _29841_);
  and (_29843_, _29842_, _10470_);
  nand (_29845_, _29843_, _29840_);
  nor (_29846_, _10470_, _29748_);
  nor (_29847_, _29846_, _10481_);
  and (_29848_, _29847_, _29845_);
  or (_29849_, _29848_, _29754_);
  nand (_29850_, _29849_, _10484_);
  nor (_29851_, _10484_, _10048_);
  nor (_29852_, _29851_, _10494_);
  nand (_29853_, _29852_, _29850_);
  nor (_29854_, _29742_, _10488_);
  nor (_29856_, _29854_, _10493_);
  and (_29857_, _29856_, _29853_);
  or (_29858_, _29857_, _29753_);
  nand (_29859_, _29858_, _03422_);
  nor (_29860_, _29741_, _03422_);
  nor (_29861_, _29860_, _10503_);
  nand (_29862_, _29861_, _29859_);
  nor (_29863_, _10502_, _29748_);
  nor (_29864_, _29863_, _03861_);
  nand (_29865_, _29864_, _29862_);
  and (_29867_, _10201_, _03861_);
  nor (_29868_, _29867_, _11528_);
  nand (_29869_, _29868_, _29865_);
  nor (_29870_, _10510_, _29748_);
  nor (_29871_, _29870_, _07559_);
  nand (_29872_, _29871_, _29869_);
  nor (_29873_, _10200_, _03415_);
  nor (_29874_, _29873_, _10521_);
  nand (_29875_, _29874_, _29872_);
  nor (_29876_, _29742_, _10517_);
  nor (_29878_, _29876_, _10520_);
  nand (_29879_, _29878_, _29875_);
  nor (_29880_, _10519_, _10048_);
  nor (_29881_, _29880_, _10525_);
  and (_29882_, _29881_, _29879_);
  and (_29883_, _29758_, _10525_);
  nor (_29884_, _29883_, _29882_);
  or (_29885_, _29884_, _06306_);
  or (_29886_, _29748_, _06305_);
  and (_29887_, _29886_, _04694_);
  nand (_29889_, _29887_, _29885_);
  and (_29890_, _10201_, _03839_);
  nor (_29891_, _29890_, _08456_);
  nand (_29892_, _29891_, _29889_);
  and (_29893_, _10048_, _08456_);
  nor (_29894_, _29893_, _10540_);
  nand (_29895_, _29894_, _29892_);
  nor (_29896_, _10570_, \oc8051_golden_model_1.DPH [4]);
  nor (_29897_, _29896_, _10571_);
  nor (_29898_, _29897_, _10541_);
  nor (_29900_, _29898_, _10544_);
  and (_29901_, _29900_, _29895_);
  or (_29902_, _29901_, _29752_);
  nand (_29903_, _29902_, _10580_);
  and (_29904_, _10048_, _08783_);
  and (_29905_, _29758_, _10146_);
  or (_29906_, _29905_, _29904_);
  and (_29907_, _29906_, _10145_);
  nor (_29908_, _29907_, _10587_);
  nand (_29909_, _29908_, _29903_);
  nor (_29911_, _29741_, _10585_);
  nor (_29912_, _29911_, _10590_);
  nand (_29913_, _29912_, _29909_);
  nor (_29914_, _10589_, _29748_);
  nor (_29915_, _29914_, _03838_);
  nand (_29916_, _29915_, _29913_);
  and (_29917_, _10201_, _03838_);
  nor (_29918_, _29917_, _10598_);
  and (_29919_, _29918_, _29916_);
  or (_29920_, _29919_, _29751_);
  nand (_29922_, _29920_, _10602_);
  nor (_29923_, _29758_, _10146_);
  nor (_29924_, _10048_, _08783_);
  nor (_29925_, _29924_, _10602_);
  not (_29926_, _29925_);
  nor (_29927_, _29926_, _29923_);
  nor (_29928_, _29927_, _10616_);
  nand (_29929_, _29928_, _29922_);
  nor (_29930_, _29741_, _10612_);
  nor (_29931_, _29930_, _10615_);
  nand (_29933_, _29931_, _29929_);
  nor (_29934_, _29748_, _10614_);
  nor (_29935_, _29934_, _03866_);
  nand (_29936_, _29935_, _29933_);
  and (_29937_, _10201_, _03866_);
  nor (_29938_, _29937_, _10623_);
  and (_29939_, _29938_, _29936_);
  or (_29940_, _29939_, _29750_);
  nand (_29941_, _29940_, _10030_);
  nor (_29942_, _29758_, \oc8051_golden_model_1.PSW [7]);
  nor (_29944_, _10048_, _08059_);
  nor (_29945_, _29944_, _10030_);
  not (_29946_, _29945_);
  nor (_29947_, _29946_, _29942_);
  nor (_29948_, _29947_, _10628_);
  nand (_29949_, _29948_, _29941_);
  nor (_29950_, _29741_, _10027_);
  nor (_29951_, _29950_, _08528_);
  nand (_29952_, _29951_, _29949_);
  nor (_29953_, _29748_, _08527_);
  nor (_29955_, _29953_, _03835_);
  nand (_29956_, _29955_, _29952_);
  and (_29957_, _10201_, _03835_);
  nor (_29958_, _29957_, _10640_);
  and (_29959_, _29958_, _29956_);
  or (_29960_, _29959_, _29749_);
  nand (_29961_, _29960_, _10015_);
  nor (_29962_, _29758_, _08059_);
  nor (_29963_, _10048_, \oc8051_golden_model_1.PSW [7]);
  nor (_29964_, _29963_, _10015_);
  not (_29966_, _29964_);
  nor (_29967_, _29966_, _29962_);
  nor (_29968_, _29967_, _10646_);
  nand (_29969_, _29968_, _29961_);
  nor (_29970_, _29741_, _10012_);
  nor (_29971_, _29970_, _10011_);
  nand (_29972_, _29971_, _29969_);
  nor (_29973_, _29748_, _10010_);
  nor (_29974_, _29973_, _08006_);
  nand (_29975_, _29974_, _29972_);
  and (_29976_, _29742_, _08006_);
  nor (_29977_, _29976_, _03974_);
  and (_29978_, _29977_, _29975_);
  nor (_29979_, _05898_, _11621_);
  or (_29980_, _29979_, _03474_);
  or (_29981_, _29980_, _29978_);
  and (_29982_, _29748_, _03474_);
  nor (_29983_, _29982_, _03831_);
  nand (_29984_, _29983_, _29981_);
  nor (_29985_, _10200_, _10860_);
  and (_29988_, _29815_, _10860_);
  or (_29989_, _29988_, _04386_);
  nor (_29990_, _29989_, _29985_);
  nor (_29991_, _29990_, _10669_);
  nand (_29992_, _29991_, _29984_);
  nor (_29993_, _29741_, _10008_);
  nor (_29994_, _29993_, _09990_);
  nand (_29995_, _29994_, _29992_);
  nor (_29996_, _29748_, _09989_);
  nor (_29997_, _29996_, _07964_);
  and (_29999_, _29997_, _29995_);
  or (_30000_, _29999_, _29747_);
  nand (_30001_, _30000_, _03708_);
  and (_30002_, _05898_, _03707_);
  nor (_30003_, _30002_, _03394_);
  and (_30004_, _30003_, _30001_);
  and (_30005_, _10048_, _03394_);
  or (_30006_, _30005_, _03705_);
  nor (_30007_, _30006_, _30004_);
  nor (_30008_, _29787_, _10860_);
  and (_30010_, _10201_, _10860_);
  nor (_30011_, _30010_, _30008_);
  nor (_30012_, _30011_, _03706_);
  or (_30013_, _30012_, _30007_);
  and (_30014_, _30013_, _10887_);
  nor (_30015_, _29741_, _10887_);
  or (_30016_, _30015_, _30014_);
  nand (_30017_, _30016_, _03704_);
  and (_30018_, _29748_, _03703_);
  nor (_30019_, _30018_, _27375_);
  nand (_30021_, _30019_, _30017_);
  nor (_30022_, _29742_, _10894_);
  nor (_30023_, _30022_, _03833_);
  nand (_30024_, _30023_, _30021_);
  and (_30025_, _04446_, _03833_);
  nor (_30026_, _30025_, _03400_);
  and (_30027_, _30026_, _30024_);
  and (_30028_, _10048_, _03400_);
  or (_30029_, _30028_, _03384_);
  or (_30030_, _30029_, _30027_);
  nor (_30032_, _30011_, _03385_);
  nor (_30033_, _30032_, _10911_);
  nand (_30034_, _30033_, _30030_);
  nor (_30035_, _29742_, _10910_);
  nor (_30036_, _30035_, _03701_);
  nand (_30037_, _30036_, _30034_);
  and (_30038_, _29748_, _03701_);
  nor (_30039_, _30038_, _26323_);
  nand (_30040_, _30039_, _30037_);
  nor (_30041_, _29742_, _10917_);
  nor (_30043_, _30041_, _03841_);
  and (_30044_, _30043_, _30040_);
  or (_30045_, _30044_, _29745_);
  and (_30046_, _10048_, _03399_);
  nor (_30047_, _30046_, _10928_);
  and (_30048_, _30047_, _30045_);
  nor (_30049_, _30048_, _29743_);
  or (_30050_, _30049_, _42912_);
  or (_30051_, _42908_, \oc8051_golden_model_1.PC [12]);
  and (_30052_, _30051_, _41654_);
  and (_43283_, _30052_, _30050_);
  nor (_30054_, _09998_, \oc8051_golden_model_1.PC [13]);
  nor (_30055_, _30054_, _09999_);
  and (_30056_, _30055_, _10928_);
  or (_30057_, _30055_, _10008_);
  or (_30058_, _30055_, _10012_);
  or (_30059_, _10044_, _10016_);
  and (_30060_, _30059_, _10015_);
  or (_30061_, _30055_, _10027_);
  or (_30062_, _10044_, _10031_);
  and (_30064_, _30062_, _10030_);
  or (_30065_, _10046_, _10045_);
  not (_30066_, _30065_);
  nor (_30067_, _30066_, _10133_);
  and (_30068_, _30066_, _10133_);
  or (_30069_, _30068_, _30067_);
  or (_30070_, _30069_, _08783_);
  or (_30071_, _10044_, _10146_);
  and (_30072_, _30071_, _10145_);
  and (_30073_, _30072_, _30070_);
  or (_30075_, _10044_, _06305_);
  and (_30076_, _10195_, _07559_);
  or (_30077_, _30055_, _10488_);
  and (_30078_, _30055_, _10481_);
  or (_30079_, _10198_, _10197_);
  not (_30080_, _30079_);
  nor (_30081_, _30080_, _10295_);
  and (_30082_, _30080_, _10295_);
  or (_30083_, _30082_, _30081_);
  and (_30084_, _30083_, _10183_);
  and (_30086_, _10195_, _10181_);
  or (_30087_, _30086_, _30084_);
  and (_30088_, _30087_, _03854_);
  nand (_30089_, _10423_, _10196_);
  or (_30090_, _30083_, _10423_);
  and (_30091_, _30090_, _10425_);
  and (_30092_, _30091_, _30089_);
  and (_30093_, _10044_, _03750_);
  or (_30094_, _30083_, _26387_);
  nand (_30095_, _26387_, _10196_);
  and (_30097_, _30095_, _03757_);
  and (_30098_, _30097_, _30094_);
  and (_30099_, _30069_, _10324_);
  and (_30100_, _10326_, _10044_);
  or (_30101_, _30100_, _30099_);
  and (_30102_, _30101_, _10320_);
  or (_30103_, _30055_, _28144_);
  not (_30104_, _04112_);
  or (_30105_, _10044_, _30104_);
  nor (_30106_, _04615_, \oc8051_golden_model_1.PC [13]);
  nand (_30108_, _30106_, _04944_);
  and (_30109_, _30108_, _30105_);
  or (_30110_, _30109_, _04234_);
  and (_30111_, _30110_, _30103_);
  and (_30112_, _10044_, _04111_);
  and (_30113_, _30055_, _25715_);
  or (_30114_, _30113_, _30112_);
  or (_30115_, _30114_, _30111_);
  and (_30116_, _30115_, _06140_);
  or (_30117_, _30116_, _04624_);
  or (_30119_, _30117_, _30102_);
  and (_30120_, _30119_, _04630_);
  or (_30121_, _30120_, _10355_);
  or (_30122_, _30121_, _30098_);
  or (_30123_, _30055_, _10360_);
  and (_30124_, _30123_, _10359_);
  and (_30125_, _30124_, _30122_);
  and (_30126_, _10366_, _10044_);
  or (_30127_, _30126_, _10365_);
  or (_30128_, _30127_, _30125_);
  or (_30130_, _30055_, _10364_);
  and (_30131_, _30130_, _03751_);
  and (_30132_, _30131_, _30128_);
  or (_30133_, _30132_, _30093_);
  and (_30134_, _30133_, _10375_);
  and (_30135_, _30055_, _10377_);
  or (_30136_, _30135_, _10382_);
  or (_30137_, _30136_, _30134_);
  or (_30138_, _10381_, _10044_);
  and (_30139_, _30138_, _10388_);
  and (_30141_, _30139_, _30137_);
  or (_30142_, _30141_, _30092_);
  and (_30143_, _30142_, _03855_);
  or (_30144_, _30143_, _30088_);
  and (_30145_, _30144_, _10433_);
  or (_30146_, _30083_, _10446_);
  nand (_30147_, _10446_, _10196_);
  and (_30148_, _30147_, _03847_);
  and (_30149_, _30148_, _30146_);
  or (_30150_, _30083_, _10462_);
  nand (_30152_, _10462_, _10196_);
  and (_30153_, _30152_, _03773_);
  and (_30154_, _30153_, _30150_);
  or (_30155_, _30154_, _30149_);
  nand (_30156_, _30055_, _10431_);
  nand (_30157_, _30156_, _10470_);
  or (_30158_, _30157_, _30155_);
  or (_30159_, _30158_, _30145_);
  or (_30160_, _10470_, _10044_);
  and (_30161_, _30160_, _10477_);
  and (_30163_, _30161_, _30159_);
  or (_30164_, _30163_, _30078_);
  and (_30165_, _30164_, _10484_);
  and (_30166_, _10485_, _10044_);
  or (_30167_, _30166_, _10494_);
  or (_30168_, _30167_, _30165_);
  and (_30169_, _30168_, _30077_);
  or (_30170_, _30169_, _10493_);
  or (_30171_, _10044_, _10492_);
  and (_30172_, _30171_, _03422_);
  and (_30174_, _30172_, _30170_);
  nand (_30175_, _30055_, _03547_);
  nand (_30176_, _30175_, _10502_);
  or (_30177_, _30176_, _30174_);
  or (_30178_, _10502_, _10044_);
  and (_30179_, _30178_, _09806_);
  and (_30180_, _30179_, _30177_);
  nand (_30181_, _10195_, _03861_);
  nand (_30182_, _30181_, _10510_);
  or (_30183_, _30182_, _30180_);
  or (_30185_, _10510_, _10044_);
  and (_30186_, _30185_, _03415_);
  and (_30187_, _30186_, _30183_);
  or (_30188_, _30187_, _30076_);
  and (_30189_, _30188_, _10517_);
  and (_30190_, _30055_, _10521_);
  or (_30191_, _30190_, _10520_);
  or (_30192_, _30191_, _30189_);
  or (_30193_, _10519_, _10044_);
  and (_30194_, _30193_, _10526_);
  and (_30196_, _30194_, _30192_);
  and (_30197_, _30069_, _10525_);
  or (_30198_, _30197_, _06306_);
  or (_30199_, _30198_, _30196_);
  and (_30200_, _30199_, _30075_);
  or (_30201_, _30200_, _03839_);
  nand (_30202_, _10196_, _03839_);
  and (_30203_, _30202_, _08457_);
  and (_30204_, _30203_, _30201_);
  and (_30205_, _10044_, _08456_);
  or (_30207_, _30205_, _30204_);
  and (_30208_, _30207_, _10541_);
  or (_30209_, _10571_, \oc8051_golden_model_1.DPH [5]);
  nor (_30210_, _10572_, _10541_);
  and (_30211_, _30210_, _30209_);
  or (_30212_, _30211_, _10544_);
  or (_30213_, _30212_, _30208_);
  or (_30214_, _10543_, _10044_);
  and (_30215_, _30214_, _10580_);
  and (_30216_, _30215_, _30213_);
  or (_30218_, _30216_, _30073_);
  and (_30219_, _30218_, _10585_);
  and (_30220_, _30055_, _10587_);
  or (_30221_, _30220_, _10590_);
  or (_30222_, _30221_, _30219_);
  or (_30223_, _10589_, _10044_);
  and (_30224_, _30223_, _04703_);
  and (_30225_, _30224_, _30222_);
  nand (_30226_, _10195_, _03838_);
  nand (_30227_, _30226_, _10597_);
  or (_30229_, _30227_, _30225_);
  or (_30230_, _10597_, _10044_);
  and (_30231_, _30230_, _10602_);
  and (_30232_, _30231_, _30229_);
  or (_30233_, _30069_, _10146_);
  or (_30234_, _10044_, _08783_);
  and (_30235_, _30234_, _10601_);
  and (_30236_, _30235_, _30233_);
  or (_30237_, _30236_, _30232_);
  and (_30238_, _30237_, _10612_);
  and (_30240_, _30055_, _10616_);
  or (_30241_, _30240_, _10615_);
  or (_30242_, _30241_, _30238_);
  or (_30243_, _10044_, _10614_);
  and (_30244_, _30243_, _04708_);
  and (_30245_, _30244_, _30242_);
  nand (_30246_, _10195_, _03866_);
  nand (_30247_, _30246_, _10031_);
  or (_30248_, _30247_, _30245_);
  and (_30249_, _30248_, _30064_);
  or (_30251_, _30069_, \oc8051_golden_model_1.PSW [7]);
  or (_30252_, _10044_, _08059_);
  and (_30253_, _30252_, _10029_);
  and (_30254_, _30253_, _30251_);
  or (_30255_, _30254_, _10628_);
  or (_30256_, _30255_, _30249_);
  and (_30257_, _30256_, _30061_);
  or (_30258_, _30257_, _08528_);
  or (_30259_, _10044_, _08527_);
  and (_30260_, _30259_, _06532_);
  and (_30262_, _30260_, _30258_);
  nand (_30263_, _10195_, _03835_);
  nand (_30264_, _30263_, _10016_);
  or (_30265_, _30264_, _30262_);
  and (_30266_, _30265_, _30060_);
  or (_30267_, _30069_, _08059_);
  or (_30268_, _10044_, \oc8051_golden_model_1.PSW [7]);
  and (_30269_, _30268_, _10014_);
  and (_30270_, _30269_, _30267_);
  or (_30271_, _30270_, _10646_);
  or (_30273_, _30271_, _30266_);
  and (_30274_, _30273_, _30058_);
  or (_30275_, _30274_, _10011_);
  or (_30276_, _10044_, _10010_);
  and (_30277_, _30276_, _08007_);
  and (_30278_, _30277_, _30275_);
  and (_30279_, _30055_, _08006_);
  or (_30280_, _30279_, _03974_);
  or (_30281_, _30280_, _30278_);
  nand (_30282_, _05799_, _03974_);
  and (_30284_, _30282_, _30281_);
  or (_30285_, _30284_, _03474_);
  or (_30286_, _10044_, _06543_);
  and (_30287_, _30286_, _04386_);
  and (_30288_, _30287_, _30285_);
  or (_30289_, _30083_, _10861_);
  or (_30290_, _10195_, _10860_);
  and (_30291_, _30290_, _03831_);
  and (_30292_, _30291_, _30289_);
  or (_30293_, _30292_, _10669_);
  or (_30295_, _30293_, _30288_);
  and (_30296_, _30295_, _30057_);
  or (_30297_, _30296_, _09990_);
  or (_30298_, _10044_, _09989_);
  and (_30299_, _30298_, _10870_);
  and (_30300_, _30299_, _30297_);
  and (_30301_, _30055_, _07964_);
  or (_30302_, _30301_, _03707_);
  or (_30303_, _30302_, _30300_);
  nand (_30304_, _05799_, _03707_);
  and (_30305_, _30304_, _30303_);
  or (_30306_, _30305_, _03394_);
  or (_30307_, _10044_, _03395_);
  and (_30308_, _30307_, _03706_);
  and (_30309_, _30308_, _30306_);
  or (_30310_, _30083_, _10860_);
  nand (_30311_, _10196_, _10860_);
  and (_30312_, _30311_, _30310_);
  and (_30313_, _30312_, _03705_);
  or (_30314_, _30313_, _10888_);
  or (_30317_, _30314_, _30309_);
  or (_30318_, _30055_, _10887_);
  and (_30319_, _30318_, _03704_);
  and (_30320_, _30319_, _30317_);
  nand (_30321_, _10044_, _03703_);
  nand (_30322_, _30321_, _10894_);
  or (_30323_, _30322_, _30320_);
  or (_30324_, _30055_, _10894_);
  and (_30325_, _30324_, _06956_);
  and (_30326_, _30325_, _30323_);
  nor (_30328_, _04034_, _06956_);
  or (_30329_, _30328_, _03400_);
  or (_30330_, _30329_, _30326_);
  or (_30331_, _10044_, _10904_);
  and (_30332_, _30331_, _03385_);
  and (_30333_, _30332_, _30330_);
  and (_30334_, _30312_, _03384_);
  or (_30335_, _30334_, _10911_);
  or (_30336_, _30335_, _30333_);
  or (_30337_, _30055_, _10910_);
  and (_30339_, _30337_, _03702_);
  and (_30340_, _30339_, _30336_);
  nand (_30341_, _10044_, _03701_);
  nand (_30342_, _30341_, _10917_);
  or (_30343_, _30342_, _30340_);
  or (_30344_, _30055_, _10917_);
  and (_30345_, _30344_, _10921_);
  and (_30346_, _30345_, _30343_);
  nor (_30347_, _04034_, _10921_);
  or (_30348_, _30347_, _03399_);
  or (_30350_, _30348_, _30346_);
  or (_30351_, _10044_, _10930_);
  and (_30352_, _30351_, _10929_);
  and (_30353_, _30352_, _30350_);
  or (_30354_, _30353_, _30056_);
  or (_30355_, _30354_, _42912_);
  or (_30356_, _42908_, \oc8051_golden_model_1.PC [13]);
  and (_30357_, _30356_, _41654_);
  and (_43284_, _30357_, _30355_);
  nor (_30358_, _09999_, \oc8051_golden_model_1.PC [14]);
  nor (_30360_, _30358_, _10000_);
  nor (_30361_, _30360_, _10929_);
  nor (_30362_, _30360_, _10870_);
  not (_30363_, _10038_);
  nor (_30364_, _30363_, _10016_);
  nor (_30365_, _30363_, _10031_);
  nor (_30366_, _10597_, _30363_);
  nor (_30367_, _10543_, _30363_);
  nor (_30368_, _10470_, _10038_);
  nor (_30369_, _30360_, _10364_);
  not (_30371_, _30360_);
  nor (_30372_, _30371_, _10360_);
  or (_30373_, _10316_, _10189_);
  and (_30374_, _10297_, _10193_);
  nor (_30375_, _30374_, _10298_);
  not (_30376_, _30375_);
  or (_30377_, _30376_, _10314_);
  and (_30378_, _30377_, _30373_);
  or (_30379_, _30378_, _04630_);
  and (_30381_, _10135_, _10042_);
  nor (_30384_, _30381_, _10136_);
  and (_30386_, _30384_, _10324_);
  and (_30388_, _10326_, _10038_);
  nor (_30390_, _30388_, _30386_);
  nand (_30392_, _30390_, _10320_);
  or (_30394_, _04624_, _03757_);
  nor (_30396_, _30360_, _28144_);
  and (_30398_, _30363_, _04112_);
  nor (_30400_, _04615_, \oc8051_golden_model_1.PC [14]);
  and (_30402_, _30400_, _04944_);
  nor (_30404_, _30402_, _30398_);
  nor (_30405_, _30404_, _04234_);
  nor (_30406_, _30405_, _30396_);
  nor (_30407_, _30371_, _10344_);
  and (_30408_, _10038_, _04111_);
  nor (_30409_, _30408_, _10320_);
  not (_30410_, _30409_);
  nor (_30411_, _30410_, _30407_);
  not (_30412_, _30411_);
  nor (_30413_, _30412_, _30406_);
  nor (_30415_, _30413_, _30394_);
  nand (_30416_, _30415_, _30392_);
  nand (_30417_, _30416_, _30379_);
  and (_30418_, _30417_, _10354_);
  or (_30419_, _30418_, _30372_);
  nand (_30420_, _30419_, _10359_);
  nor (_30421_, _10359_, _30363_);
  nor (_30422_, _30421_, _10365_);
  and (_30423_, _30422_, _30420_);
  or (_30424_, _30423_, _30369_);
  nand (_30426_, _30424_, _03751_);
  nor (_30427_, _10038_, _03751_);
  nor (_30428_, _30427_, _10377_);
  and (_30429_, _30428_, _30426_);
  nor (_30430_, _30371_, _10375_);
  or (_30431_, _30430_, _30429_);
  nand (_30432_, _30431_, _10381_);
  nor (_30433_, _10381_, _30363_);
  nor (_30434_, _30433_, _10425_);
  nand (_30435_, _30434_, _30432_);
  and (_30437_, _10423_, _10188_);
  nor (_30438_, _30376_, _10423_);
  or (_30439_, _30438_, _10388_);
  nor (_30440_, _30439_, _30437_);
  nor (_30441_, _30440_, _03854_);
  nand (_30442_, _30441_, _30435_);
  nand (_30443_, _10188_, _10181_);
  or (_30444_, _30376_, _10181_);
  nand (_30445_, _30444_, _30443_);
  nand (_30446_, _30445_, _03854_);
  nand (_30448_, _30446_, _30442_);
  nand (_30449_, _30448_, _10433_);
  and (_30450_, _10446_, _10188_);
  and (_30451_, _30375_, _27160_);
  or (_30452_, _30451_, _30450_);
  and (_30453_, _30452_, _03847_);
  nor (_30454_, _30375_, _10462_);
  and (_30455_, _10462_, _10189_);
  or (_30456_, _30455_, _04216_);
  nor (_30457_, _30456_, _30454_);
  nor (_30459_, _30457_, _30453_);
  and (_30460_, _30360_, _10431_);
  not (_30461_, _30460_);
  and (_30462_, _30461_, _10470_);
  and (_30463_, _30462_, _30459_);
  and (_30464_, _30463_, _30449_);
  or (_30465_, _30464_, _30368_);
  nand (_30466_, _30465_, _10477_);
  nor (_30467_, _30360_, _10477_);
  nor (_30468_, _30467_, _10485_);
  nand (_30470_, _30468_, _30466_);
  nor (_30471_, _10484_, _30363_);
  nor (_30472_, _30471_, _10494_);
  nand (_30473_, _30472_, _30470_);
  nor (_30474_, _30360_, _10488_);
  nor (_30475_, _30474_, _10493_);
  and (_30476_, _30475_, _30473_);
  nor (_30477_, _30363_, _10492_);
  or (_30478_, _30477_, _03547_);
  or (_30479_, _30478_, _30476_);
  nor (_30481_, _30360_, _03422_);
  nor (_30482_, _30481_, _10503_);
  nand (_30483_, _30482_, _30479_);
  nor (_30484_, _10502_, _30363_);
  nor (_30485_, _30484_, _03861_);
  nand (_30486_, _30485_, _30483_);
  nor (_30487_, _10188_, _09806_);
  nor (_30488_, _30487_, _11528_);
  nand (_30489_, _30488_, _30486_);
  nor (_30490_, _10510_, _30363_);
  nor (_30492_, _30490_, _07559_);
  nand (_30493_, _30492_, _30489_);
  nor (_30494_, _10188_, _03415_);
  nor (_30495_, _30494_, _10521_);
  nand (_30496_, _30495_, _30493_);
  nor (_30497_, _30371_, _10517_);
  nor (_30498_, _30497_, _10520_);
  nand (_30499_, _30498_, _30496_);
  nor (_30500_, _10519_, _10038_);
  nor (_30501_, _30500_, _10525_);
  and (_30503_, _30501_, _30499_);
  and (_30504_, _30384_, _10525_);
  nor (_30505_, _30504_, _30503_);
  or (_30506_, _30505_, _06306_);
  or (_30507_, _30363_, _06305_);
  and (_30508_, _30507_, _04694_);
  nand (_30509_, _30508_, _30506_);
  nor (_30510_, _10188_, _04694_);
  nor (_30511_, _30510_, _08456_);
  nand (_30512_, _30511_, _30509_);
  and (_30513_, _10038_, _08456_);
  nor (_30514_, _30513_, _10540_);
  nand (_30515_, _30514_, _30512_);
  nor (_30516_, _10572_, \oc8051_golden_model_1.DPH [6]);
  nor (_30517_, _30516_, _10573_);
  nor (_30518_, _30517_, _10541_);
  nor (_30519_, _30518_, _10544_);
  and (_30520_, _30519_, _30515_);
  or (_30521_, _30520_, _30367_);
  nand (_30522_, _30521_, _10580_);
  nor (_30524_, _10038_, _10146_);
  nor (_30525_, _30384_, _08783_);
  or (_30526_, _30525_, _10580_);
  nor (_30527_, _30526_, _30524_);
  nor (_30528_, _30527_, _10587_);
  nand (_30529_, _30528_, _30522_);
  nor (_30530_, _30360_, _10585_);
  nor (_30531_, _30530_, _10590_);
  nand (_30532_, _30531_, _30529_);
  nor (_30533_, _10589_, _30363_);
  nor (_30535_, _30533_, _03838_);
  nand (_30536_, _30535_, _30532_);
  nor (_30537_, _10188_, _04703_);
  nor (_30538_, _30537_, _10598_);
  and (_30539_, _30538_, _30536_);
  or (_30540_, _30539_, _30366_);
  nand (_30541_, _30540_, _10602_);
  nor (_30542_, _10038_, _08783_);
  nor (_30543_, _30384_, _10146_);
  or (_30544_, _30543_, _10602_);
  or (_30546_, _30544_, _30542_);
  and (_30547_, _30546_, _10612_);
  nand (_30548_, _30547_, _30541_);
  nor (_30549_, _30360_, _10612_);
  nor (_30550_, _30549_, _10615_);
  nand (_30551_, _30550_, _30548_);
  nor (_30552_, _30363_, _10614_);
  nor (_30553_, _30552_, _03866_);
  nand (_30554_, _30553_, _30551_);
  nor (_30555_, _10188_, _04708_);
  nor (_30557_, _30555_, _10623_);
  and (_30558_, _30557_, _30554_);
  or (_30559_, _30558_, _30365_);
  nand (_30560_, _30559_, _10030_);
  nor (_30561_, _30384_, \oc8051_golden_model_1.PSW [7]);
  nor (_30562_, _10038_, _08059_);
  nor (_30563_, _30562_, _10030_);
  not (_30564_, _30563_);
  nor (_30565_, _30564_, _30561_);
  nor (_30566_, _30565_, _10628_);
  nand (_30568_, _30566_, _30560_);
  nor (_30569_, _30360_, _10027_);
  nor (_30570_, _30569_, _08528_);
  nand (_30571_, _30570_, _30568_);
  nor (_30572_, _30363_, _08527_);
  nor (_30573_, _30572_, _03835_);
  nand (_30574_, _30573_, _30571_);
  nor (_30575_, _10188_, _06532_);
  nor (_30576_, _30575_, _10640_);
  and (_30577_, _30576_, _30574_);
  or (_30579_, _30577_, _30364_);
  nand (_30580_, _30579_, _10015_);
  nand (_30581_, _10038_, _08059_);
  nand (_30582_, _30384_, \oc8051_golden_model_1.PSW [7]);
  and (_30583_, _30582_, _30581_);
  or (_30584_, _30583_, _10015_);
  and (_30585_, _30584_, _30580_);
  nand (_30586_, _30585_, _10012_);
  nor (_30587_, _30360_, _10012_);
  nor (_30588_, _30587_, _10011_);
  nand (_30590_, _30588_, _30586_);
  nor (_30591_, _30363_, _10010_);
  nor (_30592_, _30591_, _08006_);
  nand (_30593_, _30592_, _30590_);
  nor (_30594_, _30360_, _08007_);
  nor (_30595_, _30594_, _03974_);
  and (_30596_, _30595_, _30593_);
  nor (_30597_, _06013_, _11621_);
  or (_30598_, _30597_, _03474_);
  or (_30599_, _30598_, _30596_);
  nor (_30601_, _10038_, _06543_);
  nor (_30602_, _30601_, _03831_);
  nand (_30603_, _30602_, _30599_);
  nor (_30604_, _10188_, _10860_);
  and (_30605_, _30376_, _10860_);
  or (_30606_, _30605_, _04386_);
  or (_30607_, _30606_, _30604_);
  and (_30608_, _30607_, _10008_);
  nand (_30609_, _30608_, _30603_);
  nor (_30610_, _30360_, _10008_);
  nor (_30612_, _30610_, _09990_);
  nand (_30613_, _30612_, _30609_);
  nor (_30614_, _30363_, _09989_);
  nor (_30615_, _30614_, _07964_);
  and (_30616_, _30615_, _30613_);
  or (_30617_, _30616_, _30362_);
  nand (_30618_, _30617_, _03708_);
  and (_30619_, _06013_, _03707_);
  nor (_30620_, _30619_, _03394_);
  and (_30621_, _30620_, _30618_);
  and (_30623_, _10038_, _03394_);
  or (_30624_, _30623_, _03705_);
  nor (_30625_, _30624_, _30621_);
  and (_30626_, _10189_, _10860_);
  nor (_30627_, _30375_, _10860_);
  nor (_30628_, _30627_, _30626_);
  nor (_30629_, _30628_, _03706_);
  or (_30630_, _30629_, _30625_);
  and (_30631_, _30630_, _10887_);
  nor (_30632_, _30360_, _10887_);
  or (_30634_, _30632_, _30631_);
  nand (_30635_, _30634_, _03704_);
  and (_30636_, _30363_, _03703_);
  nor (_30637_, _30636_, _27375_);
  nand (_30638_, _30637_, _30635_);
  nor (_30639_, _30371_, _10894_);
  nor (_30640_, _30639_, _03833_);
  nand (_30641_, _30640_, _30638_);
  and (_30642_, _03833_, _03740_);
  nor (_30643_, _30642_, _03400_);
  and (_30645_, _30643_, _30641_);
  and (_30646_, _10038_, _03400_);
  or (_30647_, _30646_, _03384_);
  or (_30648_, _30647_, _30645_);
  nor (_30649_, _30628_, _03385_);
  nor (_30650_, _30649_, _10911_);
  nand (_30651_, _30650_, _30648_);
  nor (_30652_, _30371_, _10910_);
  nor (_30653_, _30652_, _03701_);
  nand (_30654_, _30653_, _30651_);
  and (_30656_, _30363_, _03701_);
  nor (_30657_, _30656_, _26323_);
  nand (_30658_, _30657_, _30654_);
  nor (_30659_, _30371_, _10917_);
  nor (_30660_, _30659_, _03841_);
  nand (_30661_, _30660_, _30658_);
  and (_30662_, _03841_, _03740_);
  nor (_30663_, _30662_, _03399_);
  nand (_30664_, _30663_, _30661_);
  and (_30665_, _10038_, _03399_);
  nor (_30667_, _30665_, _10928_);
  and (_30668_, _30667_, _30664_);
  nor (_30669_, _30668_, _30361_);
  or (_30670_, _30669_, _42912_);
  or (_30671_, _42908_, \oc8051_golden_model_1.PC [14]);
  and (_30672_, _30671_, _41654_);
  and (_43285_, _30672_, _30670_);
  nor (_30673_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_30674_, _30673_, _05330_);
  and (_30675_, _10943_, \oc8051_golden_model_1.P2 [0]);
  nand (_30677_, _11074_, _03558_);
  or (_30678_, _11074_, _03558_);
  and (_30679_, _30678_, _30677_);
  and (_30680_, _30679_, _05380_);
  or (_30681_, _30680_, _30675_);
  and (_30682_, _30681_, _03959_);
  and (_30683_, _05380_, _04608_);
  or (_30684_, _30683_, _30675_);
  or (_30685_, _30684_, _06994_);
  and (_30686_, _11074_, _05380_);
  or (_30688_, _30686_, _30675_);
  or (_30689_, _30688_, _04630_);
  and (_30690_, _05380_, \oc8051_golden_model_1.ACC [0]);
  or (_30691_, _30690_, _30675_);
  and (_30692_, _30691_, _04615_);
  and (_30693_, _04616_, \oc8051_golden_model_1.P2 [0]);
  or (_30694_, _30693_, _03757_);
  or (_30695_, _30694_, _30692_);
  and (_30696_, _30695_, _03697_);
  and (_30697_, _30696_, _30689_);
  not (_30699_, _06104_);
  and (_30700_, _30699_, \oc8051_golden_model_1.P2 [0]);
  and (_30701_, _06110_, \oc8051_golden_model_1.P0 [0]);
  and (_30702_, _06104_, \oc8051_golden_model_1.P2 [0]);
  or (_30703_, _30702_, _30701_);
  and (_30704_, _06112_, \oc8051_golden_model_1.P1 [0]);
  and (_30705_, _06106_, \oc8051_golden_model_1.P3 [0]);
  or (_30706_, _30705_, _30704_);
  nor (_30707_, _30706_, _30703_);
  and (_30708_, _30707_, _10768_);
  nand (_30710_, _30708_, _10765_);
  or (_30711_, _30710_, _05651_);
  or (_30712_, _30711_, _10753_);
  and (_30713_, _30712_, _06104_);
  or (_30714_, _30713_, _30700_);
  and (_30715_, _30714_, _03696_);
  or (_30716_, _30715_, _30697_);
  and (_30717_, _30716_, _04537_);
  and (_30718_, _30684_, _03755_);
  or (_30719_, _30718_, _03750_);
  or (_30721_, _30719_, _30717_);
  or (_30722_, _30691_, _03751_);
  and (_30723_, _30722_, _03692_);
  and (_30724_, _30723_, _30721_);
  and (_30725_, _30675_, _03691_);
  or (_30726_, _30725_, _03684_);
  or (_30727_, _30726_, _30724_);
  or (_30728_, _30688_, _03685_);
  and (_30729_, _30728_, _03680_);
  and (_30730_, _30729_, _30727_);
  or (_30732_, _30700_, _14175_);
  and (_30733_, _30732_, _03679_);
  and (_30734_, _30733_, _30714_);
  or (_30735_, _30734_, _07544_);
  or (_30736_, _30735_, _30730_);
  and (_30737_, _30736_, _30685_);
  or (_30738_, _30737_, _04678_);
  and (_30739_, _06935_, _05380_);
  or (_30740_, _30675_, _04679_);
  or (_30741_, _30740_, _30739_);
  and (_30743_, _30741_, _03415_);
  and (_30744_, _30743_, _30738_);
  and (_30745_, _06466_, \oc8051_golden_model_1.P0 [0]);
  and (_30746_, _06470_, \oc8051_golden_model_1.P1 [0]);
  and (_30747_, _06474_, \oc8051_golden_model_1.P2 [0]);
  and (_30748_, _06476_, \oc8051_golden_model_1.P3 [0]);
  or (_30749_, _30748_, _30747_);
  or (_30750_, _30749_, _30746_);
  nor (_30751_, _30750_, _30745_);
  and (_30752_, _30751_, _12114_);
  and (_30754_, _30752_, _12102_);
  nand (_30755_, _30754_, _12095_);
  or (_30756_, _30755_, _12074_);
  and (_30757_, _30756_, _05380_);
  or (_30758_, _30757_, _30675_);
  and (_30759_, _30758_, _07559_);
  or (_30760_, _30759_, _30744_);
  or (_30761_, _30760_, _08854_);
  nand (_30762_, _11074_, _04326_);
  nor (_30763_, _11074_, _04326_);
  not (_30765_, _30763_);
  and (_30766_, _30765_, _30762_);
  and (_30767_, _30766_, _05380_);
  or (_30768_, _30675_, _04703_);
  or (_30769_, _30768_, _30767_);
  and (_30770_, _05380_, _06428_);
  or (_30771_, _30770_, _30675_);
  or (_30772_, _30771_, _04694_);
  and (_30773_, _30772_, _04701_);
  and (_30774_, _30773_, _30769_);
  and (_30776_, _30774_, _30761_);
  or (_30777_, _30776_, _30682_);
  and (_30778_, _30777_, _04708_);
  nand (_30779_, _30771_, _03866_);
  nor (_30780_, _30779_, _30686_);
  or (_30781_, _30780_, _30778_);
  and (_30782_, _30781_, _04706_);
  not (_30783_, _11074_);
  or (_30784_, _30675_, _30783_);
  and (_30785_, _30691_, _03967_);
  and (_30787_, _30785_, _30784_);
  or (_30788_, _30787_, _03835_);
  or (_30789_, _30788_, _30782_);
  and (_30790_, _30762_, _05380_);
  or (_30791_, _30675_, _06532_);
  or (_30792_, _30791_, _30790_);
  and (_30793_, _30792_, _06537_);
  and (_30794_, _30793_, _30789_);
  and (_30795_, _30677_, _05380_);
  or (_30796_, _30795_, _30675_);
  and (_30797_, _30796_, _03954_);
  or (_30798_, _30797_, _03703_);
  or (_30799_, _30798_, _30794_);
  or (_30800_, _30688_, _03704_);
  and (_30801_, _30800_, _03385_);
  and (_30802_, _30801_, _30799_);
  and (_30803_, _30675_, _03384_);
  or (_30804_, _30803_, _03701_);
  or (_30805_, _30804_, _30802_);
  or (_30806_, _30688_, _03702_);
  and (_30809_, _30806_, _42908_);
  and (_30810_, _30809_, _30805_);
  or (_43288_, _30810_, _30674_);
  nor (_30811_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_30812_, _30811_, _05330_);
  or (_30813_, _05380_, \oc8051_golden_model_1.P2 [1]);
  and (_30814_, _11057_, _04515_);
  nor (_30815_, _11057_, _04515_);
  nor (_30816_, _30815_, _30814_);
  or (_30817_, _30816_, _10943_);
  and (_30819_, _30817_, _03838_);
  nand (_30820_, _05380_, _04515_);
  and (_30821_, _30820_, _03839_);
  or (_30822_, _30821_, _30819_);
  and (_30823_, _30822_, _30813_);
  nor (_30824_, _11195_, _11075_);
  and (_30825_, _30824_, _05380_);
  not (_30826_, _30825_);
  and (_30827_, _30826_, _30813_);
  or (_30828_, _30827_, _04630_);
  nand (_30830_, _05380_, _03491_);
  and (_30831_, _30830_, _30813_);
  and (_30832_, _30831_, _04615_);
  and (_30833_, _04616_, \oc8051_golden_model_1.P2 [1]);
  or (_30834_, _30833_, _03757_);
  or (_30835_, _30834_, _30832_);
  and (_30836_, _30835_, _03697_);
  and (_30837_, _30836_, _30828_);
  and (_30838_, _30699_, \oc8051_golden_model_1.P2 [1]);
  and (_30839_, _06110_, \oc8051_golden_model_1.P0 [1]);
  and (_30841_, _06104_, \oc8051_golden_model_1.P2 [1]);
  nor (_30842_, _30841_, _30839_);
  and (_30843_, _06112_, \oc8051_golden_model_1.P1 [1]);
  and (_30844_, _06106_, \oc8051_golden_model_1.P3 [1]);
  nor (_30845_, _30844_, _30843_);
  and (_30846_, _30845_, _30842_);
  and (_30847_, _30846_, _10713_);
  and (_30848_, _30847_, _10710_);
  and (_30849_, _30848_, _05601_);
  nand (_30850_, _30849_, _10699_);
  and (_30852_, _30850_, _06104_);
  or (_30853_, _30852_, _30838_);
  and (_30854_, _30853_, _03696_);
  or (_30855_, _30854_, _03755_);
  or (_30856_, _30855_, _30837_);
  and (_30857_, _10943_, \oc8051_golden_model_1.P2 [1]);
  and (_30858_, _05380_, _04813_);
  or (_30859_, _30858_, _30857_);
  or (_30860_, _30859_, _04537_);
  and (_30861_, _30860_, _30856_);
  or (_30863_, _30861_, _03750_);
  or (_30864_, _30831_, _03751_);
  and (_30865_, _30864_, _03692_);
  and (_30866_, _30865_, _30863_);
  nor (_30867_, _30849_, _10697_);
  and (_30868_, _30867_, _06104_);
  or (_30869_, _30868_, _30838_);
  and (_30870_, _30869_, _03691_);
  or (_30871_, _30870_, _03684_);
  or (_30872_, _30871_, _30866_);
  or (_30874_, _30849_, _10699_);
  and (_30875_, _30852_, _30874_);
  or (_30876_, _30838_, _03685_);
  or (_30877_, _30876_, _30875_);
  and (_30878_, _30877_, _30872_);
  and (_30879_, _30878_, _03680_);
  or (_30880_, _30867_, _12255_);
  and (_30881_, _30880_, _06104_);
  or (_30882_, _30838_, _30881_);
  and (_30883_, _30882_, _03679_);
  or (_30885_, _30883_, _07544_);
  or (_30886_, _30885_, _30879_);
  or (_30887_, _30859_, _06994_);
  and (_30888_, _30887_, _30886_);
  or (_30889_, _30888_, _04678_);
  and (_30890_, _06934_, _05380_);
  or (_30891_, _30857_, _04679_);
  or (_30892_, _30891_, _30890_);
  and (_30893_, _30892_, _03415_);
  and (_30894_, _30893_, _30889_);
  and (_30896_, _06466_, \oc8051_golden_model_1.P0 [1]);
  and (_30897_, _06470_, \oc8051_golden_model_1.P1 [1]);
  and (_30898_, _06474_, \oc8051_golden_model_1.P2 [1]);
  and (_30899_, _06476_, \oc8051_golden_model_1.P3 [1]);
  or (_30900_, _30899_, _30898_);
  or (_30901_, _30900_, _30897_);
  nor (_30902_, _30901_, _30896_);
  and (_30903_, _30902_, _12280_);
  and (_30904_, _30903_, _12294_);
  nand (_30905_, _30904_, _12310_);
  or (_30907_, _30905_, _12268_);
  and (_30908_, _30907_, _05380_);
  or (_30909_, _30908_, _30857_);
  and (_30910_, _30909_, _07559_);
  or (_30911_, _30910_, _30894_);
  and (_30912_, _30911_, _03840_);
  or (_30913_, _30912_, _30823_);
  and (_30914_, _30913_, _04701_);
  nand (_30915_, _11057_, _03491_);
  or (_30916_, _11057_, _03491_);
  and (_30918_, _30916_, _30915_);
  or (_30919_, _30918_, _10943_);
  and (_30920_, _30813_, _03959_);
  and (_30921_, _30920_, _30919_);
  or (_30922_, _30921_, _30914_);
  and (_30923_, _30922_, _04708_);
  or (_30924_, _30815_, _10943_);
  and (_30925_, _30813_, _03866_);
  and (_30926_, _30925_, _30924_);
  or (_30927_, _30926_, _30923_);
  and (_30929_, _30927_, _04706_);
  not (_30930_, _11057_);
  or (_30931_, _30857_, _30930_);
  and (_30932_, _30831_, _03967_);
  and (_30933_, _30932_, _30931_);
  or (_30934_, _30933_, _30929_);
  and (_30935_, _30934_, _03955_);
  or (_30936_, _30820_, _30930_);
  and (_30937_, _30813_, _03835_);
  and (_30938_, _30937_, _30936_);
  or (_30940_, _30915_, _10943_);
  and (_30941_, _30813_, _03954_);
  and (_30942_, _30941_, _30940_);
  or (_30943_, _30942_, _03703_);
  or (_30944_, _30943_, _30938_);
  or (_30945_, _30944_, _30935_);
  or (_30946_, _30827_, _03704_);
  and (_30947_, _30946_, _03385_);
  and (_30948_, _30947_, _30945_);
  and (_30949_, _30869_, _03384_);
  or (_30951_, _30949_, _03701_);
  or (_30952_, _30951_, _30948_);
  or (_30953_, _30857_, _03702_);
  or (_30954_, _30953_, _30825_);
  and (_30955_, _30954_, _42908_);
  and (_30956_, _30955_, _30952_);
  or (_43289_, _30956_, _30812_);
  and (_30957_, _10943_, \oc8051_golden_model_1.P2 [2]);
  nor (_30958_, _10943_, _05236_);
  or (_30959_, _30958_, _30957_);
  or (_30961_, _30959_, _06994_);
  or (_30962_, _30959_, _04537_);
  nor (_30963_, _11075_, _11046_);
  or (_30964_, _30963_, _11076_);
  and (_30965_, _30964_, _05380_);
  or (_30966_, _30965_, _30957_);
  or (_30967_, _30966_, _04630_);
  and (_30968_, _05380_, \oc8051_golden_model_1.ACC [2]);
  or (_30969_, _30968_, _30957_);
  and (_30970_, _30969_, _04615_);
  and (_30972_, _04616_, \oc8051_golden_model_1.P2 [2]);
  or (_30973_, _30972_, _03757_);
  or (_30974_, _30973_, _30970_);
  and (_30975_, _30974_, _03697_);
  and (_30976_, _30975_, _30967_);
  and (_30977_, _30699_, \oc8051_golden_model_1.P2 [2]);
  and (_30978_, _06112_, \oc8051_golden_model_1.P1 [2]);
  and (_30979_, _06106_, \oc8051_golden_model_1.P3 [2]);
  nor (_30980_, _30979_, _30978_);
  and (_30981_, _06110_, \oc8051_golden_model_1.P0 [2]);
  and (_30983_, _06104_, \oc8051_golden_model_1.P2 [2]);
  nor (_30984_, _30983_, _30981_);
  and (_30985_, _30984_, _30980_);
  and (_30986_, _30985_, _10683_);
  nand (_30987_, _30986_, _10675_);
  nor (_30988_, _30987_, _10684_);
  and (_30989_, _30988_, _05698_);
  nand (_30990_, _30989_, _10695_);
  and (_30991_, _30990_, _06104_);
  or (_30992_, _30991_, _30977_);
  and (_30994_, _30992_, _03696_);
  or (_30995_, _30994_, _03755_);
  or (_30996_, _30995_, _30976_);
  and (_30997_, _30996_, _30962_);
  or (_30998_, _30997_, _03750_);
  or (_30999_, _30969_, _03751_);
  and (_31000_, _30999_, _03692_);
  and (_31001_, _31000_, _30998_);
  nor (_31002_, _30989_, _10694_);
  and (_31003_, _31002_, _06104_);
  or (_31005_, _31003_, _30977_);
  and (_31006_, _31005_, _03691_);
  or (_31007_, _31006_, _03684_);
  or (_31008_, _31007_, _31001_);
  or (_31009_, _30989_, _10695_);
  and (_31010_, _30991_, _31009_);
  or (_31011_, _30977_, _03685_);
  or (_31012_, _31011_, _31010_);
  and (_31013_, _31012_, _03680_);
  and (_31014_, _31013_, _31008_);
  or (_31016_, _31002_, _12464_);
  and (_31017_, _31016_, _06104_);
  or (_31018_, _31017_, _30977_);
  and (_31019_, _31018_, _03679_);
  or (_31020_, _31019_, _07544_);
  or (_31021_, _31020_, _31014_);
  and (_31022_, _31021_, _30961_);
  or (_31023_, _31022_, _04678_);
  and (_31024_, _06938_, _05380_);
  or (_31025_, _30957_, _04679_);
  or (_31026_, _31025_, _31024_);
  and (_31027_, _31026_, _03415_);
  and (_31028_, _31027_, _31023_);
  and (_31029_, _06470_, \oc8051_golden_model_1.P1 [2]);
  and (_31030_, _06466_, \oc8051_golden_model_1.P0 [2]);
  and (_31031_, _06474_, \oc8051_golden_model_1.P2 [2]);
  and (_31032_, _06476_, \oc8051_golden_model_1.P3 [2]);
  or (_31033_, _31032_, _31031_);
  or (_31034_, _31033_, _31030_);
  nor (_31035_, _31034_, _31029_);
  and (_31038_, _31035_, _12489_);
  and (_31039_, _31038_, _12484_);
  nand (_31040_, _31039_, _12520_);
  or (_31041_, _31040_, _12477_);
  and (_31042_, _31041_, _05380_);
  or (_31043_, _30957_, _31042_);
  and (_31044_, _31043_, _07559_);
  or (_31045_, _31044_, _31028_);
  or (_31046_, _31045_, _08854_);
  nand (_31047_, _11046_, _04077_);
  or (_31049_, _11046_, _04077_);
  and (_31050_, _31049_, _31047_);
  and (_31051_, _31050_, _05380_);
  or (_31052_, _30957_, _04703_);
  or (_31053_, _31052_, _31051_);
  and (_31054_, _05380_, _06457_);
  or (_31055_, _31054_, _30957_);
  or (_31056_, _31055_, _04694_);
  and (_31057_, _31056_, _04701_);
  and (_31058_, _31057_, _31053_);
  and (_31060_, _31058_, _31046_);
  nand (_31061_, _11046_, _07740_);
  or (_31062_, _11046_, _07740_);
  and (_31063_, _31062_, _31061_);
  and (_31064_, _31063_, _05380_);
  or (_31065_, _31064_, _30957_);
  and (_31066_, _31065_, _03959_);
  or (_31067_, _31066_, _31060_);
  and (_31068_, _31067_, _04708_);
  or (_31069_, _30957_, _11194_);
  and (_31071_, _31055_, _03866_);
  and (_31072_, _31071_, _31069_);
  or (_31073_, _31072_, _31068_);
  and (_31074_, _31073_, _04706_);
  and (_31075_, _30969_, _03967_);
  and (_31076_, _31075_, _31069_);
  or (_31077_, _31076_, _03835_);
  or (_31078_, _31077_, _31074_);
  and (_31079_, _31047_, _05380_);
  or (_31080_, _30957_, _06532_);
  or (_31082_, _31080_, _31079_);
  and (_31083_, _31082_, _06537_);
  and (_31084_, _31083_, _31078_);
  and (_31085_, _31061_, _05380_);
  or (_31086_, _31085_, _30957_);
  and (_31087_, _31086_, _03954_);
  or (_31088_, _31087_, _03703_);
  or (_31089_, _31088_, _31084_);
  or (_31090_, _30966_, _03704_);
  and (_31091_, _31090_, _03385_);
  and (_31093_, _31091_, _31089_);
  and (_31094_, _31005_, _03384_);
  or (_31095_, _31094_, _03701_);
  or (_31096_, _31095_, _31093_);
  nor (_31097_, _11195_, _11194_);
  nor (_31098_, _31097_, _11196_);
  and (_31099_, _31098_, _05380_);
  or (_31100_, _30957_, _03702_);
  or (_31101_, _31100_, _31099_);
  and (_31102_, _31101_, _42908_);
  and (_31104_, _31102_, _31096_);
  nor (_31105_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_31106_, _31105_, _05330_);
  or (_43290_, _31106_, _31104_);
  and (_31107_, _10943_, \oc8051_golden_model_1.P2 [3]);
  nor (_31108_, _10943_, _05050_);
  or (_31109_, _31108_, _31107_);
  or (_31110_, _31109_, _06994_);
  nor (_31111_, _11076_, _11029_);
  or (_31112_, _31111_, _11077_);
  and (_31114_, _31112_, _05380_);
  or (_31115_, _31114_, _31107_);
  or (_31116_, _31115_, _04630_);
  and (_31117_, _05380_, \oc8051_golden_model_1.ACC [3]);
  or (_31118_, _31117_, _31107_);
  and (_31119_, _31118_, _04615_);
  and (_31120_, _04616_, \oc8051_golden_model_1.P2 [3]);
  or (_31121_, _31120_, _03757_);
  or (_31122_, _31121_, _31119_);
  and (_31123_, _31122_, _03697_);
  and (_31125_, _31123_, _31116_);
  and (_31126_, _30699_, \oc8051_golden_model_1.P2 [3]);
  and (_31127_, _06112_, \oc8051_golden_model_1.P1 [3]);
  and (_31128_, _06106_, \oc8051_golden_model_1.P3 [3]);
  nor (_31129_, _31128_, _31127_);
  and (_31130_, _06110_, \oc8051_golden_model_1.P0 [3]);
  and (_31131_, _06104_, \oc8051_golden_model_1.P2 [3]);
  nor (_31132_, _31131_, _31130_);
  and (_31133_, _31132_, _31129_);
  and (_31134_, _31133_, _10819_);
  and (_31136_, _31134_, _10816_);
  and (_31137_, _31136_, _05552_);
  nand (_31138_, _31137_, _10831_);
  and (_31139_, _31138_, _06104_);
  or (_31140_, _31139_, _31126_);
  and (_31141_, _31140_, _03696_);
  or (_31142_, _31141_, _03755_);
  or (_31143_, _31142_, _31125_);
  or (_31144_, _31109_, _04537_);
  and (_31145_, _31144_, _31143_);
  or (_31147_, _31145_, _03750_);
  or (_31148_, _31118_, _03751_);
  and (_31149_, _31148_, _03692_);
  and (_31150_, _31149_, _31147_);
  nor (_31151_, _31137_, _10830_);
  and (_31152_, _31151_, _06104_);
  or (_31153_, _31152_, _31126_);
  and (_31154_, _31153_, _03691_);
  or (_31155_, _31154_, _03684_);
  or (_31156_, _31155_, _31150_);
  or (_31158_, _31137_, _10831_);
  or (_31159_, _31126_, _31158_);
  and (_31160_, _31159_, _31140_);
  or (_31161_, _31160_, _03685_);
  and (_31162_, _31161_, _03680_);
  and (_31163_, _31162_, _31156_);
  or (_31164_, _31151_, _12664_);
  and (_31165_, _31164_, _06104_);
  or (_31166_, _31165_, _31126_);
  and (_31167_, _31166_, _03679_);
  or (_31169_, _31167_, _07544_);
  or (_31170_, _31169_, _31163_);
  and (_31171_, _31170_, _31110_);
  or (_31172_, _31171_, _04678_);
  and (_31173_, _06937_, _05380_);
  or (_31174_, _31107_, _04679_);
  or (_31175_, _31174_, _31173_);
  and (_31176_, _31175_, _03415_);
  and (_31177_, _31176_, _31172_);
  and (_31178_, _06470_, \oc8051_golden_model_1.P1 [3]);
  and (_31180_, _06466_, \oc8051_golden_model_1.P0 [3]);
  and (_31181_, _06474_, \oc8051_golden_model_1.P2 [3]);
  and (_31182_, _06476_, \oc8051_golden_model_1.P3 [3]);
  or (_31183_, _31182_, _31181_);
  or (_31184_, _31183_, _31180_);
  nor (_31185_, _31184_, _31178_);
  and (_31186_, _31185_, _12691_);
  and (_31187_, _31186_, _12701_);
  nand (_31188_, _31187_, _12721_);
  or (_31189_, _31188_, _12679_);
  and (_31191_, _31189_, _05380_);
  or (_31192_, _31107_, _31191_);
  and (_31193_, _31192_, _07559_);
  or (_31194_, _31193_, _31177_);
  or (_31195_, _31194_, _08854_);
  nand (_31196_, _11029_, _03946_);
  or (_31197_, _11029_, _03946_);
  and (_31198_, _31197_, _31196_);
  and (_31199_, _31198_, _05380_);
  or (_31200_, _31107_, _04703_);
  or (_31202_, _31200_, _31199_);
  and (_31203_, _05380_, _06415_);
  or (_31204_, _31203_, _31107_);
  or (_31205_, _31204_, _04694_);
  and (_31206_, _31205_, _04701_);
  and (_31207_, _31206_, _31202_);
  and (_31208_, _31207_, _31195_);
  nand (_31209_, _11029_, _07734_);
  or (_31210_, _11029_, _07734_);
  and (_31211_, _31210_, _31209_);
  and (_31213_, _31211_, _05380_);
  or (_31214_, _31213_, _31107_);
  and (_31215_, _31214_, _03959_);
  or (_31216_, _31215_, _31208_);
  and (_31217_, _31216_, _04708_);
  or (_31218_, _31107_, _11193_);
  and (_31219_, _31204_, _03866_);
  and (_31220_, _31219_, _31218_);
  or (_31221_, _31220_, _31217_);
  and (_31222_, _31221_, _04706_);
  and (_31224_, _31118_, _03967_);
  and (_31225_, _31224_, _31218_);
  or (_31226_, _31225_, _03835_);
  or (_31227_, _31226_, _31222_);
  and (_31228_, _31196_, _05380_);
  or (_31229_, _31107_, _06532_);
  or (_31230_, _31229_, _31228_);
  and (_31231_, _31230_, _06537_);
  and (_31232_, _31231_, _31227_);
  and (_31233_, _31209_, _05380_);
  or (_31235_, _31233_, _31107_);
  and (_31236_, _31235_, _03954_);
  or (_31237_, _31236_, _03703_);
  or (_31238_, _31237_, _31232_);
  or (_31239_, _31115_, _03704_);
  and (_31240_, _31239_, _03385_);
  and (_31241_, _31240_, _31238_);
  and (_31242_, _31153_, _03384_);
  or (_31243_, _31242_, _03701_);
  or (_31244_, _31243_, _31241_);
  nor (_31245_, _11196_, _11193_);
  nor (_31246_, _31245_, _11197_);
  and (_31247_, _31246_, _05380_);
  or (_31248_, _31107_, _03702_);
  or (_31249_, _31248_, _31247_);
  and (_31250_, _31249_, _42908_);
  and (_31251_, _31250_, _31244_);
  nor (_31252_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_31253_, _31252_, _05330_);
  or (_43291_, _31253_, _31251_);
  nor (_31255_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_31256_, _31255_, _05330_);
  and (_31257_, _10943_, \oc8051_golden_model_1.P2 [4]);
  nor (_31258_, _05898_, _10943_);
  or (_31259_, _31258_, _31257_);
  or (_31260_, _31259_, _06994_);
  and (_31261_, _30699_, \oc8051_golden_model_1.P2 [4]);
  and (_31262_, _06106_, \oc8051_golden_model_1.P3 [4]);
  nor (_31263_, _31262_, _10733_);
  and (_31264_, _31263_, _10740_);
  and (_31266_, _06112_, \oc8051_golden_model_1.P1 [4]);
  and (_31267_, _06104_, \oc8051_golden_model_1.P2 [4]);
  and (_31268_, _06110_, \oc8051_golden_model_1.P0 [4]);
  or (_31269_, _31268_, _31267_);
  nor (_31270_, _31269_, _31266_);
  and (_31271_, _31270_, _31264_);
  and (_31272_, _31271_, _10732_);
  and (_31273_, _31272_, _05899_);
  nor (_31274_, _31273_, _10748_);
  and (_31275_, _31274_, _06104_);
  or (_31277_, _31275_, _31261_);
  and (_31278_, _31277_, _03691_);
  nor (_31279_, _11077_, _11011_);
  or (_31280_, _31279_, _11078_);
  and (_31281_, _31280_, _05380_);
  or (_31282_, _31281_, _31257_);
  or (_31283_, _31282_, _04630_);
  and (_31284_, _05380_, \oc8051_golden_model_1.ACC [4]);
  or (_31285_, _31284_, _31257_);
  and (_31286_, _31285_, _04615_);
  and (_31288_, _04616_, \oc8051_golden_model_1.P2 [4]);
  or (_31289_, _31288_, _03757_);
  or (_31290_, _31289_, _31286_);
  and (_31291_, _31290_, _03697_);
  and (_31292_, _31291_, _31283_);
  nand (_31293_, _31273_, _10749_);
  and (_31294_, _31293_, _06104_);
  or (_31295_, _31294_, _31261_);
  and (_31296_, _31295_, _03696_);
  or (_31297_, _31296_, _03755_);
  or (_31299_, _31297_, _31292_);
  or (_31300_, _31259_, _04537_);
  and (_31301_, _31300_, _31299_);
  or (_31302_, _31301_, _03750_);
  or (_31303_, _31285_, _03751_);
  and (_31304_, _31303_, _03692_);
  and (_31305_, _31304_, _31302_);
  or (_31306_, _31305_, _31278_);
  and (_31307_, _31306_, _03685_);
  or (_31308_, _31273_, _10749_);
  or (_31310_, _31261_, _31308_);
  and (_31311_, _31310_, _03684_);
  and (_31312_, _31311_, _31295_);
  or (_31313_, _31312_, _31307_);
  and (_31314_, _31313_, _03680_);
  or (_31315_, _31274_, _12809_);
  and (_31316_, _31315_, _06104_);
  or (_31317_, _31316_, _31261_);
  and (_31318_, _31317_, _03679_);
  or (_31319_, _31318_, _07544_);
  or (_31321_, _31319_, _31314_);
  and (_31322_, _31321_, _31260_);
  or (_31323_, _31322_, _04678_);
  and (_31324_, _06942_, _05380_);
  or (_31325_, _31257_, _04679_);
  or (_31326_, _31325_, _31324_);
  and (_31327_, _31326_, _03415_);
  and (_31328_, _31327_, _31323_);
  and (_31329_, _06466_, \oc8051_golden_model_1.P0 [4]);
  and (_31330_, _06470_, \oc8051_golden_model_1.P1 [4]);
  and (_31332_, _06474_, \oc8051_golden_model_1.P2 [4]);
  and (_31333_, _06476_, \oc8051_golden_model_1.P3 [4]);
  or (_31334_, _31333_, _31332_);
  or (_31335_, _31334_, _31330_);
  nor (_31336_, _31335_, _31329_);
  and (_31337_, _31336_, _12886_);
  and (_31338_, _31337_, _12881_);
  nand (_31339_, _31338_, _12916_);
  or (_31340_, _31339_, _12874_);
  and (_31341_, _31340_, _05380_);
  or (_31343_, _31341_, _31257_);
  and (_31344_, _31343_, _07559_);
  or (_31345_, _31344_, _08854_);
  or (_31346_, _31345_, _31328_);
  nand (_31347_, _11011_, _06339_);
  or (_31348_, _11011_, _06339_);
  and (_31349_, _31348_, _31347_);
  and (_31350_, _31349_, _05380_);
  or (_31351_, _31257_, _04703_);
  or (_31352_, _31351_, _31350_);
  and (_31354_, _06422_, _05380_);
  or (_31355_, _31354_, _31257_);
  or (_31356_, _31355_, _04694_);
  and (_31357_, _31356_, _04701_);
  and (_31358_, _31357_, _31352_);
  and (_31359_, _31358_, _31346_);
  nand (_31360_, _11011_, _07640_);
  or (_31361_, _11011_, _07640_);
  and (_31362_, _31361_, _31360_);
  and (_31363_, _31362_, _05380_);
  or (_31365_, _31363_, _31257_);
  and (_31366_, _31365_, _03959_);
  or (_31367_, _31366_, _31359_);
  and (_31368_, _31367_, _04708_);
  or (_31369_, _31257_, _11192_);
  and (_31370_, _31355_, _03866_);
  and (_31371_, _31370_, _31369_);
  or (_31372_, _31371_, _31368_);
  and (_31373_, _31372_, _04706_);
  and (_31374_, _31285_, _03967_);
  and (_31376_, _31374_, _31369_);
  or (_31377_, _31376_, _03835_);
  or (_31378_, _31377_, _31373_);
  and (_31379_, _31347_, _05380_);
  or (_31380_, _31257_, _06532_);
  or (_31381_, _31380_, _31379_);
  and (_31382_, _31381_, _06537_);
  and (_31383_, _31382_, _31378_);
  and (_31384_, _31360_, _05380_);
  or (_31385_, _31384_, _31257_);
  and (_31387_, _31385_, _03954_);
  or (_31388_, _31387_, _03703_);
  or (_31389_, _31388_, _31383_);
  or (_31390_, _31282_, _03704_);
  and (_31391_, _31390_, _03385_);
  and (_31392_, _31391_, _31389_);
  and (_31393_, _31277_, _03384_);
  or (_31394_, _31393_, _03701_);
  or (_31395_, _31394_, _31392_);
  nor (_31396_, _11197_, _11192_);
  nor (_31398_, _31396_, _11198_);
  and (_31399_, _31398_, _05380_);
  or (_31400_, _31257_, _03702_);
  or (_31401_, _31400_, _31399_);
  and (_31402_, _31401_, _42908_);
  and (_31403_, _31402_, _31395_);
  or (_43292_, _31403_, _31256_);
  nor (_31404_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_31405_, _31404_, _05330_);
  and (_31406_, _10943_, \oc8051_golden_model_1.P2 [5]);
  nor (_31408_, _11078_, _11000_);
  or (_31409_, _31408_, _11079_);
  and (_31410_, _31409_, _05380_);
  or (_31411_, _31410_, _31406_);
  or (_31412_, _31411_, _04630_);
  and (_31413_, _05380_, \oc8051_golden_model_1.ACC [5]);
  or (_31414_, _31413_, _31406_);
  and (_31415_, _31414_, _04615_);
  and (_31416_, _04616_, \oc8051_golden_model_1.P2 [5]);
  or (_31417_, _31416_, _03757_);
  or (_31419_, _31417_, _31415_);
  and (_31420_, _31419_, _03697_);
  and (_31421_, _31420_, _31412_);
  and (_31422_, _30699_, \oc8051_golden_model_1.P2 [5]);
  and (_31423_, _06106_, \oc8051_golden_model_1.P3 [5]);
  nor (_31424_, _31423_, _10846_);
  and (_31425_, _31424_, _10838_);
  and (_31426_, _06112_, \oc8051_golden_model_1.P1 [5]);
  and (_31427_, _06104_, \oc8051_golden_model_1.P2 [5]);
  and (_31428_, _06110_, \oc8051_golden_model_1.P0 [5]);
  or (_31430_, _31428_, _31427_);
  nor (_31431_, _31430_, _31426_);
  and (_31432_, _31431_, _10845_);
  and (_31433_, _31432_, _31425_);
  and (_31434_, _31433_, _05800_);
  nand (_31435_, _31434_, _10856_);
  and (_31436_, _31435_, _06104_);
  or (_31437_, _31436_, _31422_);
  and (_31438_, _31437_, _03696_);
  or (_31439_, _31438_, _03755_);
  or (_31441_, _31439_, _31421_);
  nor (_31442_, _05799_, _10943_);
  or (_31443_, _31442_, _31406_);
  or (_31444_, _31443_, _04537_);
  and (_31445_, _31444_, _31441_);
  or (_31446_, _31445_, _03750_);
  or (_31447_, _31414_, _03751_);
  and (_31448_, _31447_, _03692_);
  and (_31449_, _31448_, _31446_);
  nor (_31450_, _31434_, _10855_);
  and (_31452_, _31450_, _06104_);
  or (_31453_, _31452_, _31422_);
  and (_31454_, _31453_, _03691_);
  or (_31455_, _31454_, _03684_);
  or (_31456_, _31455_, _31449_);
  or (_31457_, _31434_, _10856_);
  or (_31458_, _31422_, _31457_);
  and (_31459_, _31458_, _31437_);
  or (_31460_, _31459_, _03685_);
  and (_31461_, _31460_, _03680_);
  and (_31463_, _31461_, _31456_);
  or (_31464_, _31450_, _13008_);
  and (_31465_, _31464_, _06104_);
  or (_31466_, _31465_, _31422_);
  and (_31467_, _31466_, _03679_);
  or (_31468_, _31467_, _07544_);
  or (_31469_, _31468_, _31463_);
  or (_31470_, _31443_, _06994_);
  and (_31471_, _31470_, _31469_);
  or (_31472_, _31471_, _04678_);
  and (_31474_, _06941_, _05380_);
  or (_31475_, _31406_, _04679_);
  or (_31476_, _31475_, _31474_);
  and (_31477_, _31476_, _03415_);
  and (_31478_, _31477_, _31472_);
  and (_31479_, _06470_, \oc8051_golden_model_1.P1 [5]);
  and (_31480_, _06466_, \oc8051_golden_model_1.P0 [5]);
  and (_31481_, _06474_, \oc8051_golden_model_1.P2 [5]);
  and (_31482_, _06476_, \oc8051_golden_model_1.P3 [5]);
  or (_31483_, _31482_, _31481_);
  or (_31485_, _31483_, _31480_);
  nor (_31486_, _31485_, _31479_);
  and (_31487_, _31486_, _13084_);
  and (_31488_, _31487_, _13078_);
  nand (_31489_, _31488_, _13115_);
  or (_31490_, _31489_, _13071_);
  and (_31491_, _31490_, _05380_);
  or (_31492_, _31491_, _31406_);
  and (_31493_, _31492_, _07559_);
  or (_31494_, _31493_, _08854_);
  or (_31496_, _31494_, _31478_);
  nand (_31497_, _11000_, _06370_);
  or (_31498_, _11000_, _06370_);
  and (_31499_, _31498_, _31497_);
  and (_31500_, _31499_, _05380_);
  or (_31501_, _31406_, _04703_);
  or (_31502_, _31501_, _31500_);
  and (_31503_, _06371_, _05380_);
  or (_31504_, _31503_, _31406_);
  or (_31505_, _31504_, _04694_);
  and (_31507_, _31505_, _04701_);
  and (_31508_, _31507_, _31502_);
  and (_31509_, _31508_, _31496_);
  nand (_31510_, _11000_, _07634_);
  or (_31511_, _11000_, _07634_);
  and (_31512_, _31511_, _31510_);
  and (_31513_, _31512_, _05380_);
  or (_31514_, _31513_, _31406_);
  and (_31515_, _31514_, _03959_);
  or (_31516_, _31515_, _31509_);
  and (_31518_, _31516_, _04708_);
  or (_31519_, _31406_, _11191_);
  and (_31520_, _31504_, _03866_);
  and (_31521_, _31520_, _31519_);
  or (_31522_, _31521_, _31518_);
  and (_31523_, _31522_, _04706_);
  and (_31524_, _31414_, _03967_);
  and (_31525_, _31524_, _31519_);
  or (_31526_, _31525_, _03835_);
  or (_31527_, _31526_, _31523_);
  and (_31529_, _31497_, _05380_);
  or (_31530_, _31406_, _06532_);
  or (_31531_, _31530_, _31529_);
  and (_31532_, _31531_, _06537_);
  and (_31533_, _31532_, _31527_);
  and (_31534_, _31510_, _05380_);
  or (_31535_, _31534_, _31406_);
  and (_31536_, _31535_, _03954_);
  or (_31537_, _31536_, _03703_);
  or (_31538_, _31537_, _31533_);
  or (_31540_, _31411_, _03704_);
  and (_31541_, _31540_, _03385_);
  and (_31542_, _31541_, _31538_);
  and (_31543_, _31453_, _03384_);
  or (_31544_, _31543_, _03701_);
  or (_31545_, _31544_, _31542_);
  nor (_31546_, _11198_, _11191_);
  nor (_31547_, _31546_, _11199_);
  and (_31548_, _31547_, _05380_);
  or (_31549_, _31406_, _03702_);
  or (_31551_, _31549_, _31548_);
  and (_31552_, _31551_, _42908_);
  and (_31553_, _31552_, _31545_);
  or (_43293_, _31553_, _31405_);
  and (_31554_, _10943_, \oc8051_golden_model_1.P2 [6]);
  nor (_31555_, _06013_, _10943_);
  or (_31556_, _31555_, _31554_);
  or (_31557_, _31556_, _06994_);
  and (_31558_, _30699_, \oc8051_golden_model_1.P2 [6]);
  and (_31559_, _06110_, \oc8051_golden_model_1.P0 [6]);
  and (_31561_, _06104_, \oc8051_golden_model_1.P2 [6]);
  nor (_31562_, _31561_, _31559_);
  and (_31563_, _06112_, \oc8051_golden_model_1.P1 [6]);
  and (_31564_, _06106_, \oc8051_golden_model_1.P3 [6]);
  nor (_31565_, _31564_, _31563_);
  and (_31566_, _31565_, _31562_);
  and (_31567_, _31566_, _10792_);
  and (_31568_, _31567_, _10789_);
  and (_31569_, _31568_, _06014_);
  nor (_31570_, _31569_, _10803_);
  and (_31572_, _31570_, _06104_);
  or (_31573_, _31572_, _31558_);
  and (_31574_, _31573_, _03691_);
  nor (_31575_, _11079_, _10984_);
  or (_31576_, _31575_, _11080_);
  and (_31577_, _31576_, _05380_);
  or (_31578_, _31577_, _31554_);
  or (_31579_, _31578_, _04630_);
  and (_31580_, _05380_, \oc8051_golden_model_1.ACC [6]);
  or (_31581_, _31580_, _31554_);
  and (_31583_, _31581_, _04615_);
  and (_31584_, _04616_, \oc8051_golden_model_1.P2 [6]);
  or (_31585_, _31584_, _03757_);
  or (_31586_, _31585_, _31583_);
  and (_31587_, _31586_, _03697_);
  and (_31588_, _31587_, _31579_);
  nand (_31589_, _31569_, _10804_);
  and (_31590_, _31589_, _06104_);
  or (_31591_, _31590_, _31558_);
  and (_31592_, _31591_, _03696_);
  or (_31594_, _31592_, _03755_);
  or (_31595_, _31594_, _31588_);
  or (_31596_, _31556_, _04537_);
  and (_31597_, _31596_, _31595_);
  or (_31598_, _31597_, _03750_);
  or (_31599_, _31581_, _03751_);
  and (_31600_, _31599_, _03692_);
  and (_31601_, _31600_, _31598_);
  or (_31602_, _31601_, _31574_);
  and (_31603_, _31602_, _03685_);
  or (_31604_, _31569_, _10804_);
  or (_31605_, _31558_, _31604_);
  and (_31606_, _31605_, _03684_);
  and (_31607_, _31606_, _31591_);
  or (_31608_, _31607_, _31603_);
  and (_31609_, _31608_, _03680_);
  or (_31610_, _31570_, _13219_);
  and (_31611_, _31610_, _06104_);
  or (_31612_, _31611_, _31558_);
  and (_31613_, _31612_, _03679_);
  or (_31616_, _31613_, _07544_);
  or (_31617_, _31616_, _31609_);
  and (_31618_, _31617_, _31557_);
  or (_31619_, _31618_, _04678_);
  and (_31620_, _06933_, _05380_);
  or (_31621_, _31554_, _04679_);
  or (_31622_, _31621_, _31620_);
  and (_31623_, _31622_, _03415_);
  and (_31624_, _31623_, _31619_);
  and (_31625_, _06474_, \oc8051_golden_model_1.P2 [6]);
  and (_31627_, _06470_, \oc8051_golden_model_1.P1 [6]);
  and (_31628_, _06466_, \oc8051_golden_model_1.P0 [6]);
  nor (_31629_, _31628_, _31627_);
  nand (_31630_, _31629_, _13287_);
  or (_31631_, _31630_, _31625_);
  not (_31632_, _13292_);
  and (_31633_, _13311_, _31632_);
  nand (_31634_, _31633_, _13307_);
  not (_31635_, _13288_);
  nand (_31636_, _13314_, _31635_);
  or (_31638_, _13316_, _13318_);
  and (_31639_, _06476_, \oc8051_golden_model_1.P3 [6]);
  or (_31640_, _31639_, _13289_);
  or (_31641_, _31640_, _31638_);
  or (_31642_, _31641_, _13291_);
  or (_31643_, _31642_, _31636_);
  or (_31644_, _31643_, _31634_);
  or (_31645_, _31644_, _31631_);
  or (_31646_, _31645_, _13280_);
  and (_31647_, _31646_, _05380_);
  or (_31649_, _31647_, _31554_);
  and (_31650_, _31649_, _07559_);
  or (_31651_, _31650_, _08854_);
  or (_31652_, _31651_, _31624_);
  nand (_31653_, _10984_, _06406_);
  or (_31654_, _10984_, _06406_);
  and (_31655_, _31654_, _31653_);
  and (_31656_, _31655_, _05380_);
  or (_31657_, _31554_, _04703_);
  or (_31658_, _31657_, _31656_);
  and (_31660_, _13333_, _05380_);
  or (_31661_, _31660_, _31554_);
  or (_31662_, _31661_, _04694_);
  and (_31663_, _31662_, _04701_);
  and (_31664_, _31663_, _31658_);
  and (_31665_, _31664_, _31652_);
  nand (_31666_, _10984_, _07586_);
  or (_31667_, _10984_, _07586_);
  and (_31668_, _31667_, _31666_);
  and (_31669_, _31668_, _05380_);
  or (_31671_, _31669_, _31554_);
  and (_31672_, _31671_, _03959_);
  or (_31673_, _31672_, _31665_);
  and (_31674_, _31673_, _04708_);
  or (_31675_, _31554_, _11190_);
  and (_31676_, _31661_, _03866_);
  and (_31677_, _31676_, _31675_);
  or (_31678_, _31677_, _31674_);
  and (_31679_, _31678_, _04706_);
  and (_31680_, _31581_, _03967_);
  and (_31682_, _31680_, _31675_);
  or (_31683_, _31682_, _03835_);
  or (_31684_, _31683_, _31679_);
  and (_31685_, _31653_, _05380_);
  or (_31686_, _31554_, _06532_);
  or (_31687_, _31686_, _31685_);
  and (_31688_, _31687_, _06537_);
  and (_31689_, _31688_, _31684_);
  and (_31690_, _31666_, _05380_);
  or (_31691_, _31690_, _31554_);
  and (_31693_, _31691_, _03954_);
  or (_31694_, _31693_, _03703_);
  or (_31695_, _31694_, _31689_);
  or (_31696_, _31578_, _03704_);
  and (_31697_, _31696_, _03385_);
  and (_31698_, _31697_, _31695_);
  and (_31699_, _31573_, _03384_);
  or (_31700_, _31699_, _03701_);
  or (_31701_, _31700_, _31698_);
  or (_31702_, _11199_, _11190_);
  and (_31704_, _31702_, _11200_);
  and (_31705_, _31704_, _05380_);
  or (_31706_, _31554_, _03702_);
  or (_31707_, _31706_, _31705_);
  and (_31708_, _31707_, _42908_);
  and (_31709_, _31708_, _31701_);
  nor (_31710_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_31711_, _31710_, _05330_);
  or (_43294_, _31711_, _31709_);
  nor (_31712_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_31714_, _31712_, _05330_);
  and (_31715_, _11209_, \oc8051_golden_model_1.P3 [0]);
  and (_31716_, _30679_, _05382_);
  or (_31717_, _31716_, _31715_);
  and (_31718_, _31717_, _03959_);
  and (_31719_, _05382_, _04608_);
  or (_31720_, _31719_, _31715_);
  or (_31721_, _31720_, _06994_);
  and (_31722_, _11074_, _05382_);
  or (_31723_, _31722_, _31715_);
  or (_31725_, _31723_, _04630_);
  and (_31726_, _05382_, \oc8051_golden_model_1.ACC [0]);
  or (_31727_, _31726_, _31715_);
  and (_31728_, _31727_, _04615_);
  and (_31729_, _04616_, \oc8051_golden_model_1.P3 [0]);
  or (_31730_, _31729_, _03757_);
  or (_31731_, _31730_, _31728_);
  and (_31732_, _31731_, _03697_);
  and (_31733_, _31732_, _31725_);
  and (_31734_, _11214_, \oc8051_golden_model_1.P3 [0]);
  and (_31736_, _30712_, _06106_);
  or (_31737_, _31736_, _31734_);
  and (_31738_, _31737_, _03696_);
  or (_31739_, _31738_, _31733_);
  and (_31740_, _31739_, _04537_);
  and (_31741_, _31720_, _03755_);
  or (_31742_, _31741_, _03750_);
  or (_31743_, _31742_, _31740_);
  or (_31744_, _31727_, _03751_);
  and (_31745_, _31744_, _03692_);
  and (_31747_, _31745_, _31743_);
  and (_31748_, _31715_, _03691_);
  or (_31749_, _31748_, _03684_);
  or (_31750_, _31749_, _31747_);
  or (_31751_, _31723_, _03685_);
  and (_31752_, _31751_, _03680_);
  and (_31753_, _31752_, _31750_);
  or (_31754_, _31734_, _14175_);
  and (_31755_, _31754_, _03679_);
  and (_31756_, _31755_, _31737_);
  or (_31758_, _31756_, _07544_);
  or (_31759_, _31758_, _31753_);
  and (_31760_, _31759_, _31721_);
  or (_31761_, _31760_, _04678_);
  and (_31762_, _06935_, _05382_);
  or (_31763_, _31715_, _04679_);
  or (_31764_, _31763_, _31762_);
  and (_31765_, _31764_, _03415_);
  and (_31766_, _31765_, _31761_);
  and (_31767_, _30756_, _05382_);
  or (_31769_, _31767_, _31715_);
  and (_31770_, _31769_, _07559_);
  or (_31771_, _31770_, _31766_);
  or (_31772_, _31771_, _08854_);
  and (_31773_, _30766_, _05382_);
  or (_31774_, _31715_, _04703_);
  or (_31775_, _31774_, _31773_);
  and (_31776_, _05382_, _06428_);
  or (_31777_, _31776_, _31715_);
  or (_31778_, _31777_, _04694_);
  and (_31780_, _31778_, _04701_);
  and (_31781_, _31780_, _31775_);
  and (_31782_, _31781_, _31772_);
  or (_31783_, _31782_, _31718_);
  and (_31784_, _31783_, _04708_);
  nand (_31785_, _31777_, _03866_);
  nor (_31786_, _31785_, _31722_);
  or (_31787_, _31786_, _31784_);
  and (_31788_, _31787_, _04706_);
  or (_31789_, _31715_, _30783_);
  and (_31791_, _31727_, _03967_);
  and (_31792_, _31791_, _31789_);
  or (_31793_, _31792_, _03835_);
  or (_31794_, _31793_, _31788_);
  and (_31795_, _30762_, _05382_);
  or (_31796_, _31715_, _06532_);
  or (_31797_, _31796_, _31795_);
  and (_31798_, _31797_, _06537_);
  and (_31799_, _31798_, _31794_);
  and (_31800_, _30677_, _05382_);
  or (_31802_, _31800_, _31715_);
  and (_31803_, _31802_, _03954_);
  or (_31804_, _31803_, _03703_);
  or (_31805_, _31804_, _31799_);
  or (_31806_, _31723_, _03704_);
  and (_31807_, _31806_, _03385_);
  and (_31808_, _31807_, _31805_);
  and (_31809_, _31715_, _03384_);
  or (_31810_, _31809_, _03701_);
  or (_31811_, _31810_, _31808_);
  or (_31813_, _31723_, _03702_);
  and (_31814_, _31813_, _42908_);
  and (_31815_, _31814_, _31811_);
  or (_43295_, _31815_, _31714_);
  or (_31816_, _05382_, \oc8051_golden_model_1.P3 [1]);
  and (_31817_, _30824_, _05382_);
  not (_31818_, _31817_);
  and (_31819_, _31818_, _31816_);
  or (_31820_, _31819_, _04630_);
  nand (_31821_, _05382_, _03491_);
  and (_31823_, _31821_, _31816_);
  and (_31824_, _31823_, _04615_);
  and (_31825_, _04616_, \oc8051_golden_model_1.P3 [1]);
  or (_31826_, _31825_, _03757_);
  or (_31827_, _31826_, _31824_);
  and (_31828_, _31827_, _03697_);
  and (_31829_, _31828_, _31820_);
  and (_31830_, _11214_, \oc8051_golden_model_1.P3 [1]);
  and (_31831_, _30850_, _06106_);
  or (_31832_, _31831_, _31830_);
  and (_31834_, _31832_, _03696_);
  or (_31835_, _31834_, _03755_);
  or (_31836_, _31835_, _31829_);
  and (_31837_, _11209_, \oc8051_golden_model_1.P3 [1]);
  and (_31838_, _05382_, _04813_);
  or (_31839_, _31838_, _31837_);
  or (_31840_, _31839_, _04537_);
  and (_31841_, _31840_, _31836_);
  or (_31842_, _31841_, _03750_);
  or (_31843_, _31823_, _03751_);
  and (_31845_, _31843_, _03692_);
  and (_31846_, _31845_, _31842_);
  and (_31847_, _30867_, _06106_);
  or (_31848_, _31847_, _31830_);
  and (_31849_, _31848_, _03691_);
  or (_31850_, _31849_, _03684_);
  or (_31851_, _31850_, _31846_);
  and (_31852_, _31831_, _30874_);
  or (_31853_, _31830_, _03685_);
  or (_31854_, _31853_, _31852_);
  and (_31856_, _31854_, _31851_);
  and (_31857_, _31856_, _03680_);
  and (_31858_, _30880_, _06106_);
  or (_31859_, _31830_, _31858_);
  and (_31860_, _31859_, _03679_);
  or (_31861_, _31860_, _07544_);
  or (_31862_, _31861_, _31857_);
  or (_31863_, _31839_, _06994_);
  and (_31864_, _31863_, _31862_);
  or (_31865_, _31864_, _04678_);
  and (_31867_, _06934_, _05382_);
  or (_31868_, _31837_, _04679_);
  or (_31869_, _31868_, _31867_);
  and (_31870_, _31869_, _03415_);
  and (_31871_, _31870_, _31865_);
  and (_31872_, _30907_, _05382_);
  or (_31873_, _31872_, _31837_);
  and (_31874_, _31873_, _07559_);
  or (_31875_, _31874_, _31871_);
  and (_31876_, _31875_, _03840_);
  or (_31878_, _30816_, _11209_);
  and (_31879_, _31878_, _03838_);
  nand (_31880_, _05382_, _04515_);
  and (_31881_, _31880_, _03839_);
  or (_31882_, _31881_, _31879_);
  and (_31883_, _31882_, _31816_);
  or (_31884_, _31883_, _31876_);
  and (_31885_, _31884_, _04701_);
  or (_31886_, _30918_, _11209_);
  and (_31887_, _31816_, _03959_);
  and (_31889_, _31887_, _31886_);
  or (_31890_, _31889_, _31885_);
  and (_31891_, _31890_, _04708_);
  or (_31892_, _30815_, _11209_);
  and (_31893_, _31816_, _03866_);
  and (_31894_, _31893_, _31892_);
  or (_31895_, _31894_, _31891_);
  and (_31896_, _31895_, _04706_);
  or (_31897_, _31837_, _30930_);
  and (_31898_, _31823_, _03967_);
  and (_31900_, _31898_, _31897_);
  or (_31901_, _31900_, _31896_);
  and (_31902_, _31901_, _03955_);
  or (_31903_, _31821_, _30930_);
  and (_31904_, _31816_, _03954_);
  and (_31905_, _31904_, _31903_);
  or (_31906_, _31905_, _03703_);
  or (_31907_, _31880_, _30930_);
  and (_31908_, _31816_, _03835_);
  and (_31909_, _31908_, _31907_);
  or (_31911_, _31909_, _31906_);
  or (_31912_, _31911_, _31902_);
  or (_31913_, _31819_, _03704_);
  and (_31914_, _31913_, _03385_);
  and (_31915_, _31914_, _31912_);
  and (_31916_, _31848_, _03384_);
  or (_31917_, _31916_, _03701_);
  or (_31918_, _31917_, _31915_);
  or (_31919_, _31837_, _03702_);
  or (_31920_, _31919_, _31817_);
  and (_31922_, _31920_, _42908_);
  and (_31923_, _31922_, _31918_);
  nor (_31924_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_31925_, _31924_, _05330_);
  or (_43296_, _31925_, _31923_);
  and (_31926_, _11209_, \oc8051_golden_model_1.P3 [2]);
  nor (_31927_, _11209_, _05236_);
  or (_31928_, _31927_, _31926_);
  or (_31929_, _31928_, _06994_);
  or (_31930_, _31928_, _04537_);
  and (_31932_, _30964_, _05382_);
  or (_31933_, _31932_, _31926_);
  or (_31934_, _31933_, _04630_);
  and (_31935_, _05382_, \oc8051_golden_model_1.ACC [2]);
  or (_31936_, _31935_, _31926_);
  and (_31937_, _31936_, _04615_);
  and (_31938_, _04616_, \oc8051_golden_model_1.P3 [2]);
  or (_31939_, _31938_, _03757_);
  or (_31940_, _31939_, _31937_);
  and (_31941_, _31940_, _03697_);
  and (_31942_, _31941_, _31934_);
  and (_31943_, _11214_, \oc8051_golden_model_1.P3 [2]);
  and (_31944_, _30990_, _06106_);
  or (_31945_, _31944_, _31943_);
  and (_31946_, _31945_, _03696_);
  or (_31947_, _31946_, _03755_);
  or (_31948_, _31947_, _31942_);
  and (_31949_, _31948_, _31930_);
  or (_31950_, _31949_, _03750_);
  or (_31951_, _31936_, _03751_);
  and (_31953_, _31951_, _03692_);
  and (_31954_, _31953_, _31950_);
  and (_31955_, _31002_, _06106_);
  or (_31956_, _31955_, _31943_);
  and (_31957_, _31956_, _03691_);
  or (_31958_, _31957_, _03684_);
  or (_31959_, _31958_, _31954_);
  and (_31960_, _31944_, _31009_);
  or (_31961_, _31943_, _03685_);
  or (_31962_, _31961_, _31960_);
  and (_31964_, _31962_, _03680_);
  and (_31965_, _31964_, _31959_);
  and (_31966_, _31016_, _06106_);
  or (_31967_, _31966_, _31943_);
  and (_31968_, _31967_, _03679_);
  or (_31969_, _31968_, _07544_);
  or (_31970_, _31969_, _31965_);
  and (_31971_, _31970_, _31929_);
  or (_31972_, _31971_, _04678_);
  and (_31973_, _06938_, _05382_);
  or (_31975_, _31926_, _04679_);
  or (_31976_, _31975_, _31973_);
  and (_31977_, _31976_, _03415_);
  and (_31978_, _31977_, _31972_);
  and (_31979_, _31041_, _05382_);
  or (_31980_, _31926_, _31979_);
  and (_31981_, _31980_, _07559_);
  or (_31982_, _31981_, _31978_);
  or (_31983_, _31982_, _08854_);
  and (_31984_, _31050_, _05382_);
  or (_31986_, _31926_, _04703_);
  or (_31987_, _31986_, _31984_);
  and (_31988_, _05382_, _06457_);
  or (_31989_, _31988_, _31926_);
  or (_31990_, _31989_, _04694_);
  and (_31991_, _31990_, _04701_);
  and (_31992_, _31991_, _31987_);
  and (_31993_, _31992_, _31983_);
  and (_31994_, _31063_, _05382_);
  or (_31995_, _31994_, _31926_);
  and (_31997_, _31995_, _03959_);
  or (_31998_, _31997_, _31993_);
  and (_31999_, _31998_, _04708_);
  or (_32000_, _31926_, _11194_);
  and (_32001_, _31989_, _03866_);
  and (_32002_, _32001_, _32000_);
  or (_32003_, _32002_, _31999_);
  and (_32004_, _32003_, _04706_);
  and (_32005_, _31936_, _03967_);
  and (_32006_, _32005_, _32000_);
  or (_32008_, _32006_, _03835_);
  or (_32009_, _32008_, _32004_);
  and (_32010_, _31047_, _05382_);
  or (_32011_, _31926_, _06532_);
  or (_32012_, _32011_, _32010_);
  and (_32013_, _32012_, _06537_);
  and (_32014_, _32013_, _32009_);
  and (_32015_, _31061_, _05382_);
  or (_32016_, _32015_, _31926_);
  and (_32017_, _32016_, _03954_);
  or (_32019_, _32017_, _03703_);
  or (_32020_, _32019_, _32014_);
  or (_32021_, _31933_, _03704_);
  and (_32022_, _32021_, _03385_);
  and (_32023_, _32022_, _32020_);
  and (_32024_, _31956_, _03384_);
  or (_32025_, _32024_, _03701_);
  or (_32026_, _32025_, _32023_);
  and (_32027_, _31098_, _05382_);
  or (_32028_, _31926_, _03702_);
  or (_32030_, _32028_, _32027_);
  and (_32031_, _32030_, _42908_);
  and (_32032_, _32031_, _32026_);
  nor (_32033_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_32034_, _32033_, _05330_);
  or (_43297_, _32034_, _32032_);
  and (_32035_, _11209_, \oc8051_golden_model_1.P3 [3]);
  nor (_32036_, _11209_, _05050_);
  or (_32037_, _32036_, _32035_);
  or (_32038_, _32037_, _06994_);
  and (_32040_, _31112_, _05382_);
  or (_32041_, _32040_, _32035_);
  or (_32042_, _32041_, _04630_);
  and (_32043_, _05382_, \oc8051_golden_model_1.ACC [3]);
  or (_32044_, _32043_, _32035_);
  and (_32045_, _32044_, _04615_);
  and (_32046_, _04616_, \oc8051_golden_model_1.P3 [3]);
  or (_32047_, _32046_, _03757_);
  or (_32048_, _32047_, _32045_);
  and (_32049_, _32048_, _03697_);
  and (_32051_, _32049_, _32042_);
  and (_32052_, _11214_, \oc8051_golden_model_1.P3 [3]);
  and (_32053_, _31138_, _06106_);
  or (_32054_, _32053_, _32052_);
  and (_32055_, _32054_, _03696_);
  or (_32056_, _32055_, _03755_);
  or (_32057_, _32056_, _32051_);
  or (_32058_, _32037_, _04537_);
  and (_32059_, _32058_, _32057_);
  or (_32060_, _32059_, _03750_);
  or (_32062_, _32044_, _03751_);
  and (_32063_, _32062_, _03692_);
  and (_32064_, _32063_, _32060_);
  and (_32065_, _31151_, _06106_);
  or (_32066_, _32065_, _32052_);
  and (_32067_, _32066_, _03691_);
  or (_32068_, _32067_, _03684_);
  or (_32069_, _32068_, _32064_);
  or (_32070_, _32052_, _31158_);
  and (_32071_, _32070_, _32054_);
  or (_32073_, _32071_, _03685_);
  and (_32074_, _32073_, _03680_);
  and (_32075_, _32074_, _32069_);
  and (_32076_, _31164_, _06106_);
  or (_32077_, _32076_, _32052_);
  and (_32078_, _32077_, _03679_);
  or (_32079_, _32078_, _07544_);
  or (_32080_, _32079_, _32075_);
  and (_32081_, _32080_, _32038_);
  or (_32082_, _32081_, _04678_);
  and (_32084_, _06937_, _05382_);
  or (_32085_, _32035_, _04679_);
  or (_32086_, _32085_, _32084_);
  and (_32087_, _32086_, _03415_);
  and (_32088_, _32087_, _32082_);
  and (_32089_, _31189_, _05382_);
  or (_32090_, _32035_, _32089_);
  and (_32091_, _32090_, _07559_);
  or (_32092_, _32091_, _32088_);
  or (_32093_, _32092_, _08854_);
  and (_32095_, _31198_, _05382_);
  or (_32096_, _32035_, _04703_);
  or (_32097_, _32096_, _32095_);
  and (_32098_, _05382_, _06415_);
  or (_32099_, _32098_, _32035_);
  or (_32100_, _32099_, _04694_);
  and (_32101_, _32100_, _04701_);
  and (_32102_, _32101_, _32097_);
  and (_32103_, _32102_, _32093_);
  and (_32104_, _31211_, _05382_);
  or (_32106_, _32104_, _32035_);
  and (_32107_, _32106_, _03959_);
  or (_32108_, _32107_, _32103_);
  and (_32109_, _32108_, _04708_);
  or (_32110_, _32035_, _11193_);
  and (_32111_, _32099_, _03866_);
  and (_32112_, _32111_, _32110_);
  or (_32113_, _32112_, _32109_);
  and (_32114_, _32113_, _04706_);
  and (_32115_, _32044_, _03967_);
  and (_32117_, _32115_, _32110_);
  or (_32118_, _32117_, _03835_);
  or (_32119_, _32118_, _32114_);
  and (_32120_, _31196_, _05382_);
  or (_32121_, _32035_, _06532_);
  or (_32122_, _32121_, _32120_);
  and (_32123_, _32122_, _06537_);
  and (_32124_, _32123_, _32119_);
  and (_32125_, _31209_, _05382_);
  or (_32126_, _32125_, _32035_);
  and (_32128_, _32126_, _03954_);
  or (_32129_, _32128_, _03703_);
  or (_32130_, _32129_, _32124_);
  or (_32131_, _32041_, _03704_);
  and (_32132_, _32131_, _03385_);
  and (_32133_, _32132_, _32130_);
  and (_32134_, _32066_, _03384_);
  or (_32135_, _32134_, _03701_);
  or (_32136_, _32135_, _32133_);
  and (_32137_, _31246_, _05382_);
  or (_32139_, _32035_, _03702_);
  or (_32140_, _32139_, _32137_);
  and (_32141_, _32140_, _42908_);
  and (_32142_, _32141_, _32136_);
  nor (_32143_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_32144_, _32143_, _05330_);
  or (_43298_, _32144_, _32142_);
  and (_32145_, _11209_, \oc8051_golden_model_1.P3 [4]);
  nor (_32146_, _05898_, _11209_);
  or (_32147_, _32146_, _32145_);
  or (_32149_, _32147_, _06994_);
  and (_32150_, _11214_, \oc8051_golden_model_1.P3 [4]);
  and (_32151_, _31274_, _06106_);
  or (_32152_, _32151_, _32150_);
  and (_32153_, _32152_, _03691_);
  and (_32154_, _31280_, _05382_);
  or (_32155_, _32154_, _32145_);
  or (_32156_, _32155_, _04630_);
  and (_32157_, _05382_, \oc8051_golden_model_1.ACC [4]);
  or (_32158_, _32157_, _32145_);
  and (_32160_, _32158_, _04615_);
  and (_32161_, _04616_, \oc8051_golden_model_1.P3 [4]);
  or (_32162_, _32161_, _03757_);
  or (_32163_, _32162_, _32160_);
  and (_32164_, _32163_, _03697_);
  and (_32165_, _32164_, _32156_);
  and (_32166_, _31293_, _06106_);
  or (_32167_, _32166_, _32150_);
  and (_32168_, _32167_, _03696_);
  or (_32169_, _32168_, _03755_);
  or (_32171_, _32169_, _32165_);
  or (_32172_, _32147_, _04537_);
  and (_32173_, _32172_, _32171_);
  or (_32174_, _32173_, _03750_);
  or (_32175_, _32158_, _03751_);
  and (_32176_, _32175_, _03692_);
  and (_32177_, _32176_, _32174_);
  or (_32178_, _32177_, _32153_);
  and (_32179_, _32178_, _03685_);
  or (_32180_, _32150_, _31308_);
  and (_32182_, _32180_, _03684_);
  and (_32183_, _32182_, _32167_);
  or (_32184_, _32183_, _32179_);
  and (_32185_, _32184_, _03680_);
  and (_32186_, _31315_, _06106_);
  or (_32187_, _32186_, _32150_);
  and (_32188_, _32187_, _03679_);
  or (_32189_, _32188_, _07544_);
  or (_32190_, _32189_, _32185_);
  and (_32191_, _32190_, _32149_);
  or (_32193_, _32191_, _04678_);
  and (_32194_, _06942_, _05382_);
  or (_32195_, _32145_, _04679_);
  or (_32196_, _32195_, _32194_);
  and (_32197_, _32196_, _03415_);
  and (_32198_, _32197_, _32193_);
  and (_32199_, _31340_, _05382_);
  or (_32200_, _32199_, _32145_);
  and (_32201_, _32200_, _07559_);
  or (_32202_, _32201_, _08854_);
  or (_32204_, _32202_, _32198_);
  and (_32205_, _31349_, _05382_);
  or (_32206_, _32145_, _04703_);
  or (_32207_, _32206_, _32205_);
  and (_32208_, _06422_, _05382_);
  or (_32209_, _32208_, _32145_);
  or (_32210_, _32209_, _04694_);
  and (_32211_, _32210_, _04701_);
  and (_32212_, _32211_, _32207_);
  and (_32213_, _32212_, _32204_);
  and (_32215_, _31362_, _05382_);
  or (_32216_, _32215_, _32145_);
  and (_32217_, _32216_, _03959_);
  or (_32218_, _32217_, _32213_);
  and (_32219_, _32218_, _04708_);
  or (_32220_, _32145_, _11192_);
  and (_32221_, _32209_, _03866_);
  and (_32222_, _32221_, _32220_);
  or (_32223_, _32222_, _32219_);
  and (_32224_, _32223_, _04706_);
  and (_32226_, _32158_, _03967_);
  and (_32227_, _32226_, _32220_);
  or (_32228_, _32227_, _03835_);
  or (_32229_, _32228_, _32224_);
  and (_32230_, _31347_, _05382_);
  or (_32231_, _32145_, _06532_);
  or (_32232_, _32231_, _32230_);
  and (_32233_, _32232_, _06537_);
  and (_32234_, _32233_, _32229_);
  and (_32235_, _31360_, _05382_);
  or (_32236_, _32235_, _32145_);
  and (_32237_, _32236_, _03954_);
  or (_32238_, _32237_, _03703_);
  or (_32239_, _32238_, _32234_);
  or (_32240_, _32155_, _03704_);
  and (_32241_, _32240_, _03385_);
  and (_32242_, _32241_, _32239_);
  and (_32243_, _32152_, _03384_);
  or (_32244_, _32243_, _03701_);
  or (_32245_, _32244_, _32242_);
  and (_32248_, _31398_, _05382_);
  or (_32249_, _32145_, _03702_);
  or (_32250_, _32249_, _32248_);
  and (_32251_, _32250_, _42908_);
  and (_32252_, _32251_, _32245_);
  nor (_32253_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_32254_, _32253_, _05330_);
  or (_43299_, _32254_, _32252_);
  nor (_32255_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_32256_, _32255_, _05330_);
  and (_32258_, _11209_, \oc8051_golden_model_1.P3 [5]);
  and (_32259_, _31409_, _05382_);
  or (_32260_, _32259_, _32258_);
  or (_32261_, _32260_, _04630_);
  and (_32262_, _05382_, \oc8051_golden_model_1.ACC [5]);
  or (_32263_, _32262_, _32258_);
  and (_32264_, _32263_, _04615_);
  and (_32265_, _04616_, \oc8051_golden_model_1.P3 [5]);
  or (_32266_, _32265_, _03757_);
  or (_32267_, _32266_, _32264_);
  and (_32269_, _32267_, _03697_);
  and (_32270_, _32269_, _32261_);
  and (_32271_, _11214_, \oc8051_golden_model_1.P3 [5]);
  and (_32272_, _31435_, _06106_);
  or (_32273_, _32272_, _32271_);
  and (_32274_, _32273_, _03696_);
  or (_32275_, _32274_, _03755_);
  or (_32276_, _32275_, _32270_);
  nor (_32277_, _05799_, _11209_);
  or (_32278_, _32277_, _32258_);
  or (_32280_, _32278_, _04537_);
  and (_32281_, _32280_, _32276_);
  or (_32282_, _32281_, _03750_);
  or (_32283_, _32263_, _03751_);
  and (_32284_, _32283_, _03692_);
  and (_32285_, _32284_, _32282_);
  and (_32286_, _31450_, _06106_);
  or (_32287_, _32286_, _32271_);
  and (_32288_, _32287_, _03691_);
  or (_32289_, _32288_, _03684_);
  or (_32291_, _32289_, _32285_);
  or (_32292_, _32271_, _31457_);
  and (_32293_, _32292_, _32273_);
  or (_32294_, _32293_, _03685_);
  and (_32295_, _32294_, _03680_);
  and (_32296_, _32295_, _32291_);
  and (_32297_, _31464_, _06106_);
  or (_32298_, _32297_, _32271_);
  and (_32299_, _32298_, _03679_);
  or (_32300_, _32299_, _07544_);
  or (_32302_, _32300_, _32296_);
  or (_32303_, _32278_, _06994_);
  and (_32304_, _32303_, _32302_);
  or (_32305_, _32304_, _04678_);
  and (_32306_, _06941_, _05382_);
  or (_32307_, _32258_, _04679_);
  or (_32308_, _32307_, _32306_);
  and (_32309_, _32308_, _03415_);
  and (_32310_, _32309_, _32305_);
  and (_32311_, _31490_, _05382_);
  or (_32313_, _32311_, _32258_);
  and (_32314_, _32313_, _07559_);
  or (_32315_, _32314_, _08854_);
  or (_32316_, _32315_, _32310_);
  and (_32317_, _31499_, _05382_);
  or (_32318_, _32258_, _04703_);
  or (_32319_, _32318_, _32317_);
  and (_32320_, _06371_, _05382_);
  or (_32321_, _32320_, _32258_);
  or (_32322_, _32321_, _04694_);
  and (_32324_, _32322_, _04701_);
  and (_32325_, _32324_, _32319_);
  and (_32326_, _32325_, _32316_);
  and (_32327_, _31512_, _05382_);
  or (_32328_, _32327_, _32258_);
  and (_32329_, _32328_, _03959_);
  or (_32330_, _32329_, _32326_);
  and (_32331_, _32330_, _04708_);
  or (_32332_, _32258_, _11191_);
  and (_32333_, _32321_, _03866_);
  and (_32335_, _32333_, _32332_);
  or (_32336_, _32335_, _32331_);
  and (_32337_, _32336_, _04706_);
  and (_32338_, _32263_, _03967_);
  and (_32339_, _32338_, _32332_);
  or (_32340_, _32339_, _03835_);
  or (_32341_, _32340_, _32337_);
  and (_32342_, _31497_, _05382_);
  or (_32343_, _32258_, _06532_);
  or (_32344_, _32343_, _32342_);
  and (_32346_, _32344_, _06537_);
  and (_32347_, _32346_, _32341_);
  and (_32348_, _31510_, _05382_);
  or (_32349_, _32348_, _32258_);
  and (_32350_, _32349_, _03954_);
  or (_32351_, _32350_, _03703_);
  or (_32352_, _32351_, _32347_);
  or (_32353_, _32260_, _03704_);
  and (_32354_, _32353_, _03385_);
  and (_32355_, _32354_, _32352_);
  and (_32357_, _32287_, _03384_);
  or (_32358_, _32357_, _03701_);
  or (_32359_, _32358_, _32355_);
  and (_32360_, _31547_, _05382_);
  or (_32361_, _32258_, _03702_);
  or (_32362_, _32361_, _32360_);
  and (_32363_, _32362_, _42908_);
  and (_32364_, _32363_, _32359_);
  or (_43302_, _32364_, _32256_);
  nor (_32365_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_32367_, _32365_, _05330_);
  and (_32368_, _11209_, \oc8051_golden_model_1.P3 [6]);
  nor (_32369_, _06013_, _11209_);
  or (_32370_, _32369_, _32368_);
  or (_32371_, _32370_, _06994_);
  and (_32372_, _11214_, \oc8051_golden_model_1.P3 [6]);
  and (_32373_, _31570_, _06106_);
  or (_32374_, _32373_, _32372_);
  and (_32375_, _32374_, _03691_);
  and (_32376_, _31576_, _05382_);
  or (_32378_, _32376_, _32368_);
  or (_32379_, _32378_, _04630_);
  and (_32380_, _05382_, \oc8051_golden_model_1.ACC [6]);
  or (_32381_, _32380_, _32368_);
  and (_32382_, _32381_, _04615_);
  and (_32383_, _04616_, \oc8051_golden_model_1.P3 [6]);
  or (_32384_, _32383_, _03757_);
  or (_32385_, _32384_, _32382_);
  and (_32386_, _32385_, _03697_);
  and (_32387_, _32386_, _32379_);
  and (_32389_, _31589_, _06106_);
  or (_32390_, _32389_, _32372_);
  and (_32391_, _32390_, _03696_);
  or (_32392_, _32391_, _03755_);
  or (_32393_, _32392_, _32387_);
  or (_32394_, _32370_, _04537_);
  and (_32395_, _32394_, _32393_);
  or (_32396_, _32395_, _03750_);
  or (_32397_, _32381_, _03751_);
  and (_32398_, _32397_, _03692_);
  and (_32400_, _32398_, _32396_);
  or (_32401_, _32400_, _32375_);
  and (_32402_, _32401_, _03685_);
  or (_32403_, _32372_, _31604_);
  and (_32404_, _32403_, _03684_);
  and (_32405_, _32404_, _32390_);
  or (_32406_, _32405_, _32402_);
  and (_32407_, _32406_, _03680_);
  and (_32408_, _31610_, _06106_);
  or (_32409_, _32408_, _32372_);
  and (_32411_, _32409_, _03679_);
  or (_32412_, _32411_, _07544_);
  or (_32413_, _32412_, _32407_);
  and (_32414_, _32413_, _32371_);
  or (_32415_, _32414_, _04678_);
  and (_32416_, _06933_, _05382_);
  or (_32417_, _32368_, _04679_);
  or (_32418_, _32417_, _32416_);
  and (_32419_, _32418_, _03415_);
  and (_32420_, _32419_, _32415_);
  and (_32422_, _31646_, _05382_);
  or (_32423_, _32422_, _32368_);
  and (_32424_, _32423_, _07559_);
  or (_32425_, _32424_, _08854_);
  or (_32426_, _32425_, _32420_);
  and (_32427_, _31655_, _05382_);
  or (_32428_, _32368_, _04703_);
  or (_32429_, _32428_, _32427_);
  and (_32430_, _13333_, _05382_);
  or (_32431_, _32430_, _32368_);
  or (_32433_, _32431_, _04694_);
  and (_32434_, _32433_, _04701_);
  and (_32435_, _32434_, _32429_);
  and (_32436_, _32435_, _32426_);
  and (_32437_, _31668_, _05382_);
  or (_32438_, _32437_, _32368_);
  and (_32439_, _32438_, _03959_);
  or (_32440_, _32439_, _32436_);
  and (_32441_, _32440_, _04708_);
  or (_32442_, _32368_, _11190_);
  and (_32444_, _32431_, _03866_);
  and (_32445_, _32444_, _32442_);
  or (_32446_, _32445_, _32441_);
  and (_32447_, _32446_, _04706_);
  and (_32448_, _32381_, _03967_);
  and (_32449_, _32448_, _32442_);
  or (_32450_, _32449_, _03835_);
  or (_32451_, _32450_, _32447_);
  and (_32452_, _31653_, _05382_);
  or (_32453_, _32368_, _06532_);
  or (_32455_, _32453_, _32452_);
  and (_32456_, _32455_, _06537_);
  and (_32457_, _32456_, _32451_);
  and (_32458_, _31666_, _05382_);
  or (_32459_, _32458_, _32368_);
  and (_32460_, _32459_, _03954_);
  or (_32461_, _32460_, _03703_);
  or (_32462_, _32461_, _32457_);
  or (_32463_, _32378_, _03704_);
  and (_32464_, _32463_, _03385_);
  and (_32466_, _32464_, _32462_);
  and (_32467_, _32374_, _03384_);
  or (_32468_, _32467_, _03701_);
  or (_32469_, _32468_, _32466_);
  and (_32470_, _31704_, _05382_);
  or (_32471_, _32368_, _03702_);
  or (_32472_, _32471_, _32470_);
  and (_32473_, _32472_, _42908_);
  and (_32474_, _32473_, _32469_);
  or (_43303_, _32474_, _32367_);
  nor (_32476_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_32477_, _32476_, _05330_);
  and (_32478_, _11311_, \oc8051_golden_model_1.P0 [0]);
  and (_32479_, _30679_, _05372_);
  or (_32480_, _32479_, _32478_);
  and (_32481_, _32480_, _03959_);
  and (_32482_, _05372_, _04608_);
  or (_32483_, _32482_, _32478_);
  or (_32484_, _32483_, _06994_);
  and (_32485_, _11074_, _05372_);
  or (_32487_, _32485_, _32478_);
  or (_32488_, _32487_, _04630_);
  and (_32489_, _05372_, \oc8051_golden_model_1.ACC [0]);
  or (_32490_, _32489_, _32478_);
  and (_32491_, _32490_, _04615_);
  and (_32492_, _04616_, \oc8051_golden_model_1.P0 [0]);
  or (_32493_, _32492_, _03757_);
  or (_32494_, _32493_, _32491_);
  and (_32495_, _32494_, _03697_);
  and (_32496_, _32495_, _32488_);
  and (_32498_, _11316_, \oc8051_golden_model_1.P0 [0]);
  and (_32499_, _30712_, _06110_);
  or (_32500_, _32499_, _32498_);
  and (_32501_, _32500_, _03696_);
  or (_32502_, _32501_, _32496_);
  and (_32503_, _32502_, _04537_);
  and (_32504_, _32483_, _03755_);
  or (_32505_, _32504_, _03750_);
  or (_32506_, _32505_, _32503_);
  or (_32507_, _32490_, _03751_);
  and (_32509_, _32507_, _03692_);
  and (_32510_, _32509_, _32506_);
  and (_32511_, _32478_, _03691_);
  or (_32512_, _32511_, _03684_);
  or (_32513_, _32512_, _32510_);
  or (_32514_, _32487_, _03685_);
  and (_32515_, _32514_, _03680_);
  and (_32516_, _32515_, _32513_);
  or (_32517_, _32498_, _14175_);
  and (_32518_, _32517_, _03679_);
  and (_32520_, _32518_, _32500_);
  or (_32521_, _32520_, _07544_);
  or (_32522_, _32521_, _32516_);
  and (_32523_, _32522_, _32484_);
  or (_32524_, _32523_, _04678_);
  and (_32525_, _06935_, _05372_);
  or (_32526_, _32478_, _04679_);
  or (_32527_, _32526_, _32525_);
  and (_32528_, _32527_, _03415_);
  and (_32529_, _32528_, _32524_);
  and (_32531_, _30756_, _05372_);
  or (_32532_, _32531_, _32478_);
  and (_32533_, _32532_, _07559_);
  or (_32534_, _32533_, _32529_);
  or (_32535_, _32534_, _08854_);
  and (_32536_, _30766_, _05372_);
  or (_32537_, _32478_, _04703_);
  or (_32538_, _32537_, _32536_);
  and (_32539_, _05372_, _06428_);
  or (_32540_, _32539_, _32478_);
  or (_32541_, _32540_, _04694_);
  and (_32542_, _32541_, _04701_);
  and (_32543_, _32542_, _32538_);
  and (_32544_, _32543_, _32535_);
  or (_32545_, _32544_, _32481_);
  and (_32546_, _32545_, _04708_);
  nand (_32547_, _32540_, _03866_);
  nor (_32548_, _32547_, _32485_);
  or (_32549_, _32548_, _32546_);
  and (_32550_, _32549_, _04706_);
  or (_32553_, _32478_, _30783_);
  and (_32554_, _32490_, _03967_);
  and (_32555_, _32554_, _32553_);
  or (_32556_, _32555_, _03835_);
  or (_32557_, _32556_, _32550_);
  and (_32558_, _30762_, _05372_);
  or (_32559_, _32478_, _06532_);
  or (_32560_, _32559_, _32558_);
  and (_32561_, _32560_, _06537_);
  and (_32562_, _32561_, _32557_);
  and (_32564_, _30677_, _05372_);
  or (_32565_, _32564_, _32478_);
  and (_32566_, _32565_, _03954_);
  or (_32567_, _32566_, _03703_);
  or (_32568_, _32567_, _32562_);
  or (_32569_, _32487_, _03704_);
  and (_32570_, _32569_, _03385_);
  and (_32571_, _32570_, _32568_);
  and (_32572_, _32478_, _03384_);
  or (_32573_, _32572_, _03701_);
  or (_32575_, _32573_, _32571_);
  or (_32576_, _32487_, _03702_);
  and (_32577_, _32576_, _42908_);
  and (_32578_, _32577_, _32575_);
  or (_43304_, _32578_, _32477_);
  nor (_32579_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_32580_, _32579_, _05330_);
  or (_32581_, _05372_, \oc8051_golden_model_1.P0 [1]);
  and (_32582_, _30824_, _05372_);
  not (_32583_, _32582_);
  and (_32585_, _32583_, _32581_);
  or (_32586_, _32585_, _04630_);
  nand (_32587_, _05372_, _03491_);
  and (_32588_, _32587_, _32581_);
  and (_32589_, _32588_, _04615_);
  and (_32590_, _04616_, \oc8051_golden_model_1.P0 [1]);
  or (_32591_, _32590_, _03757_);
  or (_32592_, _32591_, _32589_);
  and (_32593_, _32592_, _03697_);
  and (_32594_, _32593_, _32586_);
  and (_32596_, _11316_, \oc8051_golden_model_1.P0 [1]);
  and (_32597_, _30850_, _06110_);
  or (_32598_, _32597_, _32596_);
  and (_32599_, _32598_, _03696_);
  or (_32600_, _32599_, _03755_);
  or (_32601_, _32600_, _32594_);
  and (_32602_, _11311_, \oc8051_golden_model_1.P0 [1]);
  and (_32603_, _05372_, _04813_);
  or (_32604_, _32603_, _32602_);
  or (_32605_, _32604_, _04537_);
  and (_32607_, _32605_, _32601_);
  or (_32608_, _32607_, _03750_);
  or (_32609_, _32588_, _03751_);
  and (_32610_, _32609_, _03692_);
  and (_32611_, _32610_, _32608_);
  and (_32612_, _30867_, _06110_);
  or (_32613_, _32612_, _32596_);
  and (_32614_, _32613_, _03691_);
  or (_32615_, _32614_, _03684_);
  or (_32616_, _32615_, _32611_);
  and (_32618_, _32597_, _30874_);
  or (_32619_, _32596_, _03685_);
  or (_32620_, _32619_, _32618_);
  and (_32621_, _32620_, _32616_);
  and (_32622_, _32621_, _03680_);
  and (_32623_, _30880_, _06110_);
  or (_32624_, _32596_, _32623_);
  and (_32625_, _32624_, _03679_);
  or (_32626_, _32625_, _07544_);
  or (_32627_, _32626_, _32622_);
  or (_32629_, _32604_, _06994_);
  and (_32630_, _32629_, _32627_);
  or (_32631_, _32630_, _04678_);
  and (_32632_, _06934_, _05372_);
  or (_32633_, _32602_, _04679_);
  or (_32634_, _32633_, _32632_);
  and (_32635_, _32634_, _03415_);
  and (_32636_, _32635_, _32631_);
  and (_32637_, _30907_, _05372_);
  or (_32638_, _32637_, _32602_);
  and (_32640_, _32638_, _07559_);
  or (_32641_, _32640_, _32636_);
  and (_32642_, _32641_, _03840_);
  or (_32643_, _30816_, _11311_);
  and (_32644_, _32643_, _03838_);
  nand (_32645_, _05372_, _04515_);
  and (_32646_, _32645_, _03839_);
  or (_32647_, _32646_, _32644_);
  and (_32648_, _32647_, _32581_);
  or (_32649_, _32648_, _32642_);
  and (_32651_, _32649_, _04701_);
  or (_32652_, _30918_, _11311_);
  and (_32653_, _32581_, _03959_);
  and (_32654_, _32653_, _32652_);
  or (_32655_, _32654_, _32651_);
  and (_32656_, _32655_, _04708_);
  or (_32657_, _30815_, _11311_);
  and (_32658_, _32581_, _03866_);
  and (_32659_, _32658_, _32657_);
  or (_32660_, _32659_, _32656_);
  and (_32662_, _32660_, _04706_);
  or (_32663_, _32602_, _30930_);
  and (_32664_, _32588_, _03967_);
  and (_32665_, _32664_, _32663_);
  or (_32666_, _32665_, _32662_);
  and (_32667_, _32666_, _03955_);
  or (_32668_, _30915_, _11311_);
  and (_32669_, _32581_, _03954_);
  and (_32670_, _32669_, _32668_);
  or (_32671_, _32670_, _03703_);
  or (_32673_, _32645_, _30930_);
  and (_32674_, _32581_, _03835_);
  and (_32675_, _32674_, _32673_);
  or (_32676_, _32675_, _32671_);
  or (_32677_, _32676_, _32667_);
  or (_32678_, _32585_, _03704_);
  and (_32679_, _32678_, _03385_);
  and (_32680_, _32679_, _32677_);
  and (_32681_, _32613_, _03384_);
  or (_32682_, _32681_, _03701_);
  or (_32684_, _32682_, _32680_);
  or (_32685_, _32602_, _03702_);
  or (_32686_, _32685_, _32582_);
  and (_32687_, _32686_, _42908_);
  and (_32688_, _32687_, _32684_);
  or (_43307_, _32688_, _32580_);
  and (_32689_, _11311_, \oc8051_golden_model_1.P0 [2]);
  nor (_32690_, _11311_, _05236_);
  or (_32691_, _32690_, _32689_);
  or (_32692_, _32691_, _06994_);
  or (_32694_, _32691_, _04537_);
  and (_32695_, _30964_, _05372_);
  or (_32696_, _32695_, _32689_);
  or (_32697_, _32696_, _04630_);
  and (_32698_, _05372_, \oc8051_golden_model_1.ACC [2]);
  or (_32699_, _32698_, _32689_);
  and (_32700_, _32699_, _04615_);
  and (_32701_, _04616_, \oc8051_golden_model_1.P0 [2]);
  or (_32702_, _32701_, _03757_);
  or (_32703_, _32702_, _32700_);
  and (_32705_, _32703_, _03697_);
  and (_32706_, _32705_, _32697_);
  and (_32707_, _11316_, \oc8051_golden_model_1.P0 [2]);
  and (_32708_, _30990_, _06110_);
  or (_32709_, _32708_, _32707_);
  and (_32710_, _32709_, _03696_);
  or (_32711_, _32710_, _03755_);
  or (_32712_, _32711_, _32706_);
  and (_32713_, _32712_, _32694_);
  or (_32714_, _32713_, _03750_);
  or (_32716_, _32699_, _03751_);
  and (_32717_, _32716_, _03692_);
  and (_32718_, _32717_, _32714_);
  and (_32719_, _31002_, _06110_);
  or (_32720_, _32719_, _32707_);
  and (_32721_, _32720_, _03691_);
  or (_32722_, _32721_, _03684_);
  or (_32723_, _32722_, _32718_);
  and (_32724_, _32708_, _31009_);
  or (_32725_, _32707_, _03685_);
  or (_32726_, _32725_, _32724_);
  and (_32727_, _32726_, _03680_);
  and (_32728_, _32727_, _32723_);
  and (_32729_, _31016_, _06110_);
  or (_32730_, _32729_, _32707_);
  and (_32731_, _32730_, _03679_);
  or (_32732_, _32731_, _07544_);
  or (_32733_, _32732_, _32728_);
  and (_32734_, _32733_, _32692_);
  or (_32735_, _32734_, _04678_);
  and (_32737_, _06938_, _05372_);
  or (_32738_, _32689_, _04679_);
  or (_32739_, _32738_, _32737_);
  and (_32740_, _32739_, _03415_);
  and (_32741_, _32740_, _32735_);
  and (_32742_, _31041_, _05372_);
  or (_32743_, _32689_, _32742_);
  and (_32744_, _32743_, _07559_);
  or (_32745_, _32744_, _32741_);
  or (_32746_, _32745_, _08854_);
  and (_32748_, _31050_, _05372_);
  or (_32749_, _32689_, _04703_);
  or (_32750_, _32749_, _32748_);
  and (_32751_, _05372_, _06457_);
  or (_32752_, _32751_, _32689_);
  or (_32753_, _32752_, _04694_);
  and (_32754_, _32753_, _04701_);
  and (_32755_, _32754_, _32750_);
  and (_32756_, _32755_, _32746_);
  and (_32757_, _31063_, _05372_);
  or (_32759_, _32757_, _32689_);
  and (_32760_, _32759_, _03959_);
  or (_32761_, _32760_, _32756_);
  and (_32762_, _32761_, _04708_);
  or (_32763_, _32689_, _11194_);
  and (_32764_, _32752_, _03866_);
  and (_32765_, _32764_, _32763_);
  or (_32766_, _32765_, _32762_);
  and (_32767_, _32766_, _04706_);
  and (_32768_, _32699_, _03967_);
  and (_32770_, _32768_, _32763_);
  or (_32771_, _32770_, _03835_);
  or (_32772_, _32771_, _32767_);
  and (_32773_, _31047_, _05372_);
  or (_32774_, _32689_, _06532_);
  or (_32775_, _32774_, _32773_);
  and (_32776_, _32775_, _06537_);
  and (_32777_, _32776_, _32772_);
  and (_32778_, _31061_, _05372_);
  or (_32779_, _32778_, _32689_);
  and (_32781_, _32779_, _03954_);
  or (_32782_, _32781_, _03703_);
  or (_32783_, _32782_, _32777_);
  or (_32784_, _32696_, _03704_);
  and (_32785_, _32784_, _03385_);
  and (_32786_, _32785_, _32783_);
  and (_32787_, _32720_, _03384_);
  or (_32788_, _32787_, _03701_);
  or (_32789_, _32788_, _32786_);
  and (_32790_, _31098_, _05372_);
  or (_32792_, _32689_, _03702_);
  or (_32793_, _32792_, _32790_);
  and (_32794_, _32793_, _42908_);
  and (_32795_, _32794_, _32789_);
  nor (_32796_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_32797_, _32796_, _05330_);
  or (_43308_, _32797_, _32795_);
  and (_32798_, _11311_, \oc8051_golden_model_1.P0 [3]);
  nor (_32799_, _11311_, _05050_);
  or (_32800_, _32799_, _32798_);
  or (_32802_, _32800_, _06994_);
  and (_32803_, _31112_, _05372_);
  or (_32804_, _32803_, _32798_);
  or (_32805_, _32804_, _04630_);
  and (_32806_, _05372_, \oc8051_golden_model_1.ACC [3]);
  or (_32807_, _32806_, _32798_);
  and (_32808_, _32807_, _04615_);
  and (_32809_, _04616_, \oc8051_golden_model_1.P0 [3]);
  or (_32810_, _32809_, _03757_);
  or (_32811_, _32810_, _32808_);
  and (_32813_, _32811_, _03697_);
  and (_32814_, _32813_, _32805_);
  and (_32815_, _11316_, \oc8051_golden_model_1.P0 [3]);
  and (_32816_, _31138_, _06110_);
  or (_32817_, _32816_, _32815_);
  and (_32818_, _32817_, _03696_);
  or (_32819_, _32818_, _03755_);
  or (_32820_, _32819_, _32814_);
  or (_32821_, _32800_, _04537_);
  and (_32822_, _32821_, _32820_);
  or (_32824_, _32822_, _03750_);
  or (_32825_, _32807_, _03751_);
  and (_32826_, _32825_, _03692_);
  and (_32827_, _32826_, _32824_);
  and (_32828_, _31151_, _06110_);
  or (_32829_, _32828_, _32815_);
  and (_32830_, _32829_, _03691_);
  or (_32831_, _32830_, _03684_);
  or (_32832_, _32831_, _32827_);
  or (_32833_, _32815_, _31158_);
  and (_32835_, _32833_, _32817_);
  or (_32836_, _32835_, _03685_);
  and (_32837_, _32836_, _03680_);
  and (_32838_, _32837_, _32832_);
  and (_32839_, _31164_, _06110_);
  or (_32840_, _32839_, _32815_);
  and (_32841_, _32840_, _03679_);
  or (_32842_, _32841_, _07544_);
  or (_32843_, _32842_, _32838_);
  and (_32844_, _32843_, _32802_);
  or (_32846_, _32844_, _04678_);
  and (_32847_, _06937_, _05372_);
  or (_32848_, _32798_, _04679_);
  or (_32849_, _32848_, _32847_);
  and (_32850_, _32849_, _03415_);
  and (_32851_, _32850_, _32846_);
  and (_32852_, _31189_, _05372_);
  or (_32853_, _32798_, _32852_);
  and (_32854_, _32853_, _07559_);
  or (_32855_, _32854_, _32851_);
  or (_32857_, _32855_, _08854_);
  and (_32858_, _31198_, _05372_);
  or (_32859_, _32798_, _04703_);
  or (_32860_, _32859_, _32858_);
  and (_32861_, _05372_, _06415_);
  or (_32862_, _32861_, _32798_);
  or (_32863_, _32862_, _04694_);
  and (_32864_, _32863_, _04701_);
  and (_32865_, _32864_, _32860_);
  and (_32866_, _32865_, _32857_);
  and (_32868_, _31211_, _05372_);
  or (_32869_, _32868_, _32798_);
  and (_32870_, _32869_, _03959_);
  or (_32871_, _32870_, _32866_);
  and (_32872_, _32871_, _04708_);
  or (_32873_, _32798_, _11193_);
  and (_32874_, _32862_, _03866_);
  and (_32875_, _32874_, _32873_);
  or (_32876_, _32875_, _32872_);
  and (_32877_, _32876_, _04706_);
  and (_32879_, _32807_, _03967_);
  and (_32880_, _32879_, _32873_);
  or (_32881_, _32880_, _03835_);
  or (_32882_, _32881_, _32877_);
  and (_32883_, _31196_, _05372_);
  or (_32884_, _32798_, _06532_);
  or (_32885_, _32884_, _32883_);
  and (_32886_, _32885_, _06537_);
  and (_32887_, _32886_, _32882_);
  and (_32888_, _31209_, _05372_);
  or (_32889_, _32888_, _32798_);
  and (_32890_, _32889_, _03954_);
  or (_32891_, _32890_, _03703_);
  or (_32892_, _32891_, _32887_);
  or (_32893_, _32804_, _03704_);
  and (_32894_, _32893_, _03385_);
  and (_32895_, _32894_, _32892_);
  and (_32896_, _32829_, _03384_);
  or (_32897_, _32896_, _03701_);
  or (_32898_, _32897_, _32895_);
  and (_32901_, _31246_, _05372_);
  or (_32902_, _32798_, _03702_);
  or (_32903_, _32902_, _32901_);
  and (_32904_, _32903_, _42908_);
  and (_32905_, _32904_, _32898_);
  nor (_32906_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_32907_, _32906_, _05330_);
  or (_43309_, _32907_, _32905_);
  and (_32908_, _11311_, \oc8051_golden_model_1.P0 [4]);
  nor (_32909_, _05898_, _11311_);
  or (_32911_, _32909_, _32908_);
  or (_32912_, _32911_, _06994_);
  and (_32913_, _11316_, \oc8051_golden_model_1.P0 [4]);
  and (_32914_, _31274_, _06110_);
  or (_32915_, _32914_, _32913_);
  and (_32916_, _32915_, _03691_);
  and (_32917_, _31280_, _05372_);
  or (_32918_, _32917_, _32908_);
  or (_32919_, _32918_, _04630_);
  and (_32920_, _05372_, \oc8051_golden_model_1.ACC [4]);
  or (_32922_, _32920_, _32908_);
  and (_32923_, _32922_, _04615_);
  and (_32924_, _04616_, \oc8051_golden_model_1.P0 [4]);
  or (_32925_, _32924_, _03757_);
  or (_32926_, _32925_, _32923_);
  and (_32927_, _32926_, _03697_);
  and (_32928_, _32927_, _32919_);
  and (_32929_, _31293_, _06110_);
  or (_32930_, _32929_, _32913_);
  and (_32931_, _32930_, _03696_);
  or (_32933_, _32931_, _03755_);
  or (_32934_, _32933_, _32928_);
  or (_32935_, _32911_, _04537_);
  and (_32936_, _32935_, _32934_);
  or (_32937_, _32936_, _03750_);
  or (_32938_, _32922_, _03751_);
  and (_32939_, _32938_, _03692_);
  and (_32940_, _32939_, _32937_);
  or (_32941_, _32940_, _32916_);
  and (_32942_, _32941_, _03685_);
  or (_32944_, _32913_, _31308_);
  and (_32945_, _32930_, _03684_);
  and (_32946_, _32945_, _32944_);
  or (_32947_, _32946_, _32942_);
  and (_32948_, _32947_, _03680_);
  and (_32949_, _31315_, _06110_);
  or (_32950_, _32949_, _32913_);
  and (_32951_, _32950_, _03679_);
  or (_32952_, _32951_, _07544_);
  or (_32953_, _32952_, _32948_);
  and (_32955_, _32953_, _32912_);
  or (_32956_, _32955_, _04678_);
  and (_32957_, _06942_, _05372_);
  or (_32958_, _32908_, _04679_);
  or (_32959_, _32958_, _32957_);
  and (_32960_, _32959_, _03415_);
  and (_32961_, _32960_, _32956_);
  and (_32962_, _31340_, _05372_);
  or (_32963_, _32962_, _32908_);
  and (_32964_, _32963_, _07559_);
  or (_32966_, _32964_, _08854_);
  or (_32967_, _32966_, _32961_);
  and (_32968_, _31349_, _05372_);
  or (_32969_, _32908_, _04703_);
  or (_32970_, _32969_, _32968_);
  and (_32971_, _06422_, _05372_);
  or (_32972_, _32971_, _32908_);
  or (_32973_, _32972_, _04694_);
  and (_32974_, _32973_, _04701_);
  and (_32975_, _32974_, _32970_);
  and (_32977_, _32975_, _32967_);
  and (_32978_, _31362_, _05372_);
  or (_32979_, _32978_, _32908_);
  and (_32980_, _32979_, _03959_);
  or (_32981_, _32980_, _32977_);
  and (_32982_, _32981_, _04708_);
  or (_32983_, _32908_, _11192_);
  and (_32984_, _32972_, _03866_);
  and (_32985_, _32984_, _32983_);
  or (_32986_, _32985_, _32982_);
  and (_32988_, _32986_, _04706_);
  and (_32989_, _32922_, _03967_);
  and (_32990_, _32989_, _32983_);
  or (_32991_, _32990_, _03835_);
  or (_32992_, _32991_, _32988_);
  and (_32993_, _31347_, _05372_);
  or (_32994_, _32908_, _06532_);
  or (_32995_, _32994_, _32993_);
  and (_32996_, _32995_, _06537_);
  and (_32997_, _32996_, _32992_);
  and (_32999_, _31360_, _05372_);
  or (_33000_, _32999_, _32908_);
  and (_33001_, _33000_, _03954_);
  or (_33002_, _33001_, _03703_);
  or (_33003_, _33002_, _32997_);
  or (_33004_, _32918_, _03704_);
  and (_33005_, _33004_, _03385_);
  and (_33006_, _33005_, _33003_);
  and (_33007_, _32915_, _03384_);
  or (_33008_, _33007_, _03701_);
  or (_33010_, _33008_, _33006_);
  and (_33011_, _31398_, _05372_);
  or (_33012_, _32908_, _03702_);
  or (_33013_, _33012_, _33011_);
  and (_33014_, _33013_, _42908_);
  and (_33015_, _33014_, _33010_);
  nor (_33016_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_33017_, _33016_, _05330_);
  or (_43310_, _33017_, _33015_);
  and (_33018_, _11311_, \oc8051_golden_model_1.P0 [5]);
  and (_33020_, _31409_, _05372_);
  or (_33021_, _33020_, _33018_);
  or (_33022_, _33021_, _04630_);
  and (_33023_, _05372_, \oc8051_golden_model_1.ACC [5]);
  or (_33024_, _33023_, _33018_);
  and (_33025_, _33024_, _04615_);
  and (_33026_, _04616_, \oc8051_golden_model_1.P0 [5]);
  or (_33027_, _33026_, _03757_);
  or (_33028_, _33027_, _33025_);
  and (_33029_, _33028_, _03697_);
  and (_33031_, _33029_, _33022_);
  and (_33032_, _11316_, \oc8051_golden_model_1.P0 [5]);
  and (_33033_, _31435_, _06110_);
  or (_33034_, _33033_, _33032_);
  and (_33035_, _33034_, _03696_);
  or (_33036_, _33035_, _03755_);
  or (_33037_, _33036_, _33031_);
  nor (_33038_, _05799_, _11311_);
  or (_33039_, _33038_, _33018_);
  or (_33040_, _33039_, _04537_);
  and (_33042_, _33040_, _33037_);
  or (_33043_, _33042_, _03750_);
  or (_33044_, _33024_, _03751_);
  and (_33045_, _33044_, _03692_);
  and (_33046_, _33045_, _33043_);
  and (_33047_, _31450_, _06110_);
  or (_33048_, _33047_, _33032_);
  and (_33049_, _33048_, _03691_);
  or (_33050_, _33049_, _03684_);
  or (_33051_, _33050_, _33046_);
  or (_33053_, _33032_, _31457_);
  and (_33054_, _33053_, _33034_);
  or (_33055_, _33054_, _03685_);
  and (_33056_, _33055_, _03680_);
  and (_33057_, _33056_, _33051_);
  and (_33058_, _31464_, _06110_);
  or (_33059_, _33058_, _33032_);
  and (_33060_, _33059_, _03679_);
  or (_33061_, _33060_, _07544_);
  or (_33062_, _33061_, _33057_);
  or (_33064_, _33039_, _06994_);
  and (_33065_, _33064_, _33062_);
  or (_33066_, _33065_, _04678_);
  and (_33067_, _06941_, _05372_);
  or (_33068_, _33018_, _04679_);
  or (_33069_, _33068_, _33067_);
  and (_33070_, _33069_, _03415_);
  and (_33071_, _33070_, _33066_);
  and (_33072_, _31490_, _05372_);
  or (_33073_, _33072_, _33018_);
  and (_33075_, _33073_, _07559_);
  or (_33076_, _33075_, _08854_);
  or (_33077_, _33076_, _33071_);
  and (_33078_, _31499_, _05372_);
  or (_33079_, _33018_, _04703_);
  or (_33080_, _33079_, _33078_);
  and (_33081_, _06371_, _05372_);
  or (_33082_, _33081_, _33018_);
  or (_33083_, _33082_, _04694_);
  and (_33084_, _33083_, _04701_);
  and (_33086_, _33084_, _33080_);
  and (_33087_, _33086_, _33077_);
  and (_33088_, _31512_, _05372_);
  or (_33089_, _33088_, _33018_);
  and (_33090_, _33089_, _03959_);
  or (_33091_, _33090_, _33087_);
  and (_33092_, _33091_, _04708_);
  or (_33093_, _33018_, _11191_);
  and (_33094_, _33082_, _03866_);
  and (_33095_, _33094_, _33093_);
  or (_33097_, _33095_, _33092_);
  and (_33098_, _33097_, _04706_);
  and (_33099_, _33024_, _03967_);
  and (_33100_, _33099_, _33093_);
  or (_33101_, _33100_, _03835_);
  or (_33102_, _33101_, _33098_);
  and (_33103_, _31497_, _05372_);
  or (_33104_, _33018_, _06532_);
  or (_33105_, _33104_, _33103_);
  and (_33106_, _33105_, _06537_);
  and (_33108_, _33106_, _33102_);
  and (_33109_, _31510_, _05372_);
  or (_33110_, _33109_, _33018_);
  and (_33111_, _33110_, _03954_);
  or (_33112_, _33111_, _03703_);
  or (_33113_, _33112_, _33108_);
  or (_33114_, _33021_, _03704_);
  and (_33115_, _33114_, _03385_);
  and (_33116_, _33115_, _33113_);
  and (_33117_, _33048_, _03384_);
  or (_33119_, _33117_, _03701_);
  or (_33120_, _33119_, _33116_);
  and (_33121_, _31547_, _05372_);
  or (_33122_, _33018_, _03702_);
  or (_33123_, _33122_, _33121_);
  and (_33124_, _33123_, _42908_);
  and (_33125_, _33124_, _33120_);
  nor (_33126_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_33127_, _33126_, _05330_);
  or (_43311_, _33127_, _33125_);
  nor (_33129_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_33130_, _33129_, _05330_);
  and (_33131_, _11311_, \oc8051_golden_model_1.P0 [6]);
  nor (_33132_, _06013_, _11311_);
  or (_33133_, _33132_, _33131_);
  or (_33134_, _33133_, _06994_);
  and (_33135_, _11316_, \oc8051_golden_model_1.P0 [6]);
  and (_33136_, _31570_, _06110_);
  or (_33137_, _33136_, _33135_);
  and (_33138_, _33137_, _03691_);
  and (_33140_, _31576_, _05372_);
  or (_33141_, _33140_, _33131_);
  or (_33142_, _33141_, _04630_);
  and (_33143_, _05372_, \oc8051_golden_model_1.ACC [6]);
  or (_33144_, _33143_, _33131_);
  and (_33145_, _33144_, _04615_);
  and (_33146_, _04616_, \oc8051_golden_model_1.P0 [6]);
  or (_33147_, _33146_, _03757_);
  or (_33148_, _33147_, _33145_);
  and (_33149_, _33148_, _03697_);
  and (_33151_, _33149_, _33142_);
  and (_33152_, _31589_, _06110_);
  or (_33153_, _33152_, _33135_);
  and (_33154_, _33153_, _03696_);
  or (_33155_, _33154_, _03755_);
  or (_33156_, _33155_, _33151_);
  or (_33157_, _33133_, _04537_);
  and (_33158_, _33157_, _33156_);
  or (_33159_, _33158_, _03750_);
  or (_33160_, _33144_, _03751_);
  and (_33162_, _33160_, _03692_);
  and (_33163_, _33162_, _33159_);
  or (_33164_, _33163_, _33138_);
  and (_33165_, _33164_, _03685_);
  or (_33166_, _33135_, _31604_);
  and (_33167_, _33166_, _03684_);
  and (_33168_, _33167_, _33153_);
  or (_33169_, _33168_, _33165_);
  and (_33170_, _33169_, _03680_);
  and (_33171_, _31610_, _06110_);
  or (_33173_, _33171_, _33135_);
  and (_33174_, _33173_, _03679_);
  or (_33175_, _33174_, _07544_);
  or (_33176_, _33175_, _33170_);
  and (_33177_, _33176_, _33134_);
  or (_33178_, _33177_, _04678_);
  and (_33179_, _06933_, _05372_);
  or (_33180_, _33131_, _04679_);
  or (_33181_, _33180_, _33179_);
  and (_33182_, _33181_, _03415_);
  and (_33184_, _33182_, _33178_);
  and (_33185_, _31646_, _05372_);
  or (_33186_, _33185_, _33131_);
  and (_33187_, _33186_, _07559_);
  or (_33188_, _33187_, _08854_);
  or (_33189_, _33188_, _33184_);
  and (_33190_, _31655_, _05372_);
  or (_33191_, _33131_, _04703_);
  or (_33192_, _33191_, _33190_);
  and (_33193_, _13333_, _05372_);
  or (_33195_, _33193_, _33131_);
  or (_33196_, _33195_, _04694_);
  and (_33197_, _33196_, _04701_);
  and (_33198_, _33197_, _33192_);
  and (_33199_, _33198_, _33189_);
  and (_33200_, _31668_, _05372_);
  or (_33201_, _33200_, _33131_);
  and (_33202_, _33201_, _03959_);
  or (_33203_, _33202_, _33199_);
  and (_33204_, _33203_, _04708_);
  or (_33206_, _33131_, _11190_);
  and (_33207_, _33195_, _03866_);
  and (_33208_, _33207_, _33206_);
  or (_33209_, _33208_, _33204_);
  and (_33210_, _33209_, _04706_);
  and (_33211_, _33144_, _03967_);
  and (_33212_, _33211_, _33206_);
  or (_33213_, _33212_, _03835_);
  or (_33214_, _33213_, _33210_);
  and (_33215_, _31653_, _05372_);
  or (_33217_, _33131_, _06532_);
  or (_33218_, _33217_, _33215_);
  and (_33219_, _33218_, _06537_);
  and (_33220_, _33219_, _33214_);
  and (_33221_, _31666_, _05372_);
  or (_33222_, _33221_, _33131_);
  and (_33223_, _33222_, _03954_);
  or (_33224_, _33223_, _03703_);
  or (_33225_, _33224_, _33220_);
  or (_33226_, _33141_, _03704_);
  and (_33228_, _33226_, _03385_);
  and (_33229_, _33228_, _33225_);
  and (_33230_, _33137_, _03384_);
  or (_33231_, _33230_, _03701_);
  or (_33232_, _33231_, _33229_);
  and (_33233_, _31704_, _05372_);
  or (_33234_, _33131_, _03702_);
  or (_33235_, _33234_, _33233_);
  and (_33236_, _33235_, _42908_);
  and (_33237_, _33236_, _33232_);
  or (_43312_, _33237_, _33130_);
  and (_33239_, _11413_, \oc8051_golden_model_1.P1 [0]);
  and (_33240_, _30679_, _05376_);
  or (_33241_, _33240_, _33239_);
  and (_33242_, _33241_, _03959_);
  and (_33243_, _11418_, \oc8051_golden_model_1.P1 [0]);
  and (_33244_, _30712_, _06112_);
  or (_33245_, _33244_, _33243_);
  or (_33246_, _33245_, _03697_);
  and (_33247_, _11074_, _05376_);
  or (_33249_, _33247_, _33239_);
  and (_33250_, _33249_, _03757_);
  and (_33251_, _04616_, \oc8051_golden_model_1.P1 [0]);
  and (_33252_, _05376_, \oc8051_golden_model_1.ACC [0]);
  or (_33253_, _33252_, _33239_);
  and (_33254_, _33253_, _04615_);
  or (_33255_, _33254_, _33251_);
  and (_33256_, _33255_, _04630_);
  or (_33257_, _33256_, _03696_);
  or (_33258_, _33257_, _33250_);
  and (_33259_, _33258_, _33246_);
  and (_33260_, _33259_, _04537_);
  and (_33261_, _05376_, _04608_);
  or (_33262_, _33261_, _33239_);
  and (_33263_, _33262_, _03755_);
  or (_33264_, _33263_, _03750_);
  or (_33265_, _33264_, _33260_);
  or (_33266_, _33253_, _03751_);
  and (_33267_, _33266_, _03692_);
  and (_33268_, _33267_, _33265_);
  and (_33271_, _33239_, _03691_);
  or (_33272_, _33271_, _03684_);
  or (_33273_, _33272_, _33268_);
  or (_33274_, _33249_, _03685_);
  and (_33275_, _33274_, _03680_);
  and (_33276_, _33275_, _33273_);
  or (_33277_, _33243_, _14175_);
  and (_33278_, _33277_, _03679_);
  and (_33279_, _33278_, _33245_);
  or (_33280_, _33279_, _07544_);
  or (_33282_, _33280_, _33276_);
  or (_33283_, _33262_, _06994_);
  and (_33284_, _33283_, _33282_);
  or (_33285_, _33284_, _04678_);
  and (_33286_, _06935_, _05376_);
  or (_33287_, _33239_, _04679_);
  or (_33288_, _33287_, _33286_);
  and (_33289_, _33288_, _03415_);
  and (_33290_, _33289_, _33285_);
  and (_33291_, _30756_, _05376_);
  or (_33293_, _33291_, _33239_);
  and (_33294_, _33293_, _07559_);
  or (_33295_, _33294_, _33290_);
  or (_33296_, _33295_, _08854_);
  and (_33297_, _30766_, _05376_);
  or (_33298_, _33239_, _04703_);
  or (_33299_, _33298_, _33297_);
  and (_33300_, _05376_, _06428_);
  or (_33301_, _33300_, _33239_);
  or (_33302_, _33301_, _04694_);
  and (_33304_, _33302_, _04701_);
  and (_33305_, _33304_, _33299_);
  and (_33306_, _33305_, _33296_);
  or (_33307_, _33306_, _33242_);
  and (_33308_, _33307_, _04708_);
  nand (_33309_, _33301_, _03866_);
  nor (_33310_, _33309_, _33247_);
  or (_33311_, _33310_, _33308_);
  and (_33312_, _33311_, _04706_);
  or (_33313_, _33239_, _30783_);
  and (_33315_, _33253_, _03967_);
  and (_33316_, _33315_, _33313_);
  or (_33317_, _33316_, _03835_);
  or (_33318_, _33317_, _33312_);
  and (_33319_, _30762_, _05376_);
  or (_33320_, _33239_, _06532_);
  or (_33321_, _33320_, _33319_);
  and (_33322_, _33321_, _06537_);
  and (_33323_, _33322_, _33318_);
  and (_33324_, _30677_, _05376_);
  or (_33326_, _33324_, _33239_);
  and (_33327_, _33326_, _03954_);
  or (_33328_, _33327_, _03703_);
  or (_33329_, _33328_, _33323_);
  or (_33330_, _33249_, _03704_);
  and (_33331_, _33330_, _03385_);
  and (_33332_, _33331_, _33329_);
  and (_33333_, _33239_, _03384_);
  or (_33334_, _33333_, _03701_);
  or (_33335_, _33334_, _33332_);
  or (_33337_, _33249_, _03702_);
  and (_33338_, _33337_, _42908_);
  and (_33339_, _33338_, _33335_);
  nor (_33340_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_33341_, _33340_, _05330_);
  or (_43313_, _33341_, _33339_);
  or (_33342_, _05376_, \oc8051_golden_model_1.P1 [1]);
  and (_33343_, _30824_, _05376_);
  not (_33344_, _33343_);
  and (_33345_, _33344_, _33342_);
  or (_33347_, _33345_, _04630_);
  nand (_33348_, _05376_, _03491_);
  and (_33349_, _33348_, _33342_);
  and (_33350_, _33349_, _04615_);
  and (_33351_, _04616_, \oc8051_golden_model_1.P1 [1]);
  or (_33352_, _33351_, _03757_);
  or (_33353_, _33352_, _33350_);
  and (_33354_, _33353_, _03697_);
  and (_33355_, _33354_, _33347_);
  and (_33356_, _11418_, \oc8051_golden_model_1.P1 [1]);
  and (_33358_, _30850_, _06112_);
  or (_33359_, _33358_, _33356_);
  and (_33360_, _33359_, _03696_);
  or (_33361_, _33360_, _03755_);
  or (_33362_, _33361_, _33355_);
  and (_33363_, _11413_, \oc8051_golden_model_1.P1 [1]);
  and (_33364_, _05376_, _04813_);
  or (_33365_, _33364_, _33363_);
  or (_33366_, _33365_, _04537_);
  and (_33367_, _33366_, _33362_);
  or (_33369_, _33367_, _03750_);
  or (_33370_, _33349_, _03751_);
  and (_33371_, _33370_, _03692_);
  and (_33372_, _33371_, _33369_);
  and (_33373_, _30867_, _06112_);
  or (_33374_, _33373_, _33356_);
  and (_33375_, _33374_, _03691_);
  or (_33376_, _33375_, _03684_);
  or (_33377_, _33376_, _33372_);
  and (_33378_, _33358_, _30874_);
  or (_33380_, _33356_, _03685_);
  or (_33381_, _33380_, _33378_);
  and (_33382_, _33381_, _33377_);
  and (_33383_, _33382_, _03680_);
  and (_33384_, _30880_, _06112_);
  or (_33385_, _33356_, _33384_);
  and (_33386_, _33385_, _03679_);
  or (_33387_, _33386_, _07544_);
  or (_33388_, _33387_, _33383_);
  or (_33389_, _33365_, _06994_);
  and (_33391_, _33389_, _33388_);
  or (_33392_, _33391_, _04678_);
  and (_33393_, _06934_, _05376_);
  or (_33394_, _33363_, _04679_);
  or (_33395_, _33394_, _33393_);
  and (_33396_, _33395_, _03415_);
  and (_33397_, _33396_, _33392_);
  and (_33398_, _30907_, _05376_);
  or (_33399_, _33398_, _33363_);
  and (_33400_, _33399_, _07559_);
  or (_33402_, _33400_, _33397_);
  and (_33403_, _33402_, _03840_);
  or (_33404_, _30816_, _11413_);
  and (_33405_, _33404_, _03838_);
  nand (_33406_, _05376_, _04515_);
  and (_33407_, _33406_, _03839_);
  or (_33408_, _33407_, _33405_);
  and (_33409_, _33408_, _33342_);
  or (_33410_, _33409_, _33403_);
  and (_33411_, _33410_, _04701_);
  or (_33413_, _30918_, _11413_);
  and (_33414_, _33342_, _03959_);
  and (_33415_, _33414_, _33413_);
  or (_33416_, _33415_, _33411_);
  and (_33417_, _33416_, _04708_);
  or (_33418_, _30815_, _11413_);
  and (_33419_, _33342_, _03866_);
  and (_33420_, _33419_, _33418_);
  or (_33421_, _33420_, _33417_);
  and (_33422_, _33421_, _04706_);
  or (_33424_, _33363_, _30930_);
  and (_33425_, _33349_, _03967_);
  and (_33426_, _33425_, _33424_);
  or (_33427_, _33426_, _33422_);
  and (_33428_, _33427_, _03955_);
  or (_33429_, _33406_, _30930_);
  and (_33430_, _33342_, _03835_);
  and (_33431_, _33430_, _33429_);
  or (_33432_, _33348_, _30930_);
  and (_33433_, _33342_, _03954_);
  and (_33435_, _33433_, _33432_);
  or (_33436_, _33435_, _03703_);
  or (_33437_, _33436_, _33431_);
  or (_33438_, _33437_, _33428_);
  or (_33439_, _33345_, _03704_);
  and (_33440_, _33439_, _03385_);
  and (_33441_, _33440_, _33438_);
  and (_33442_, _33374_, _03384_);
  or (_33443_, _33442_, _03701_);
  or (_33444_, _33443_, _33441_);
  or (_33446_, _33363_, _03702_);
  or (_33447_, _33446_, _33343_);
  and (_33448_, _33447_, _42908_);
  and (_33449_, _33448_, _33444_);
  nor (_33450_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_33451_, _33450_, _05330_);
  or (_43314_, _33451_, _33449_);
  and (_33452_, _11413_, \oc8051_golden_model_1.P1 [2]);
  nor (_33453_, _11413_, _05236_);
  or (_33454_, _33453_, _33452_);
  or (_33456_, _33454_, _06994_);
  or (_33457_, _33454_, _04537_);
  and (_33458_, _30964_, _05376_);
  or (_33459_, _33458_, _33452_);
  or (_33460_, _33459_, _04630_);
  and (_33461_, _05376_, \oc8051_golden_model_1.ACC [2]);
  or (_33462_, _33461_, _33452_);
  and (_33463_, _33462_, _04615_);
  and (_33464_, _04616_, \oc8051_golden_model_1.P1 [2]);
  or (_33465_, _33464_, _03757_);
  or (_33467_, _33465_, _33463_);
  and (_33468_, _33467_, _03697_);
  and (_33469_, _33468_, _33460_);
  and (_33470_, _11418_, \oc8051_golden_model_1.P1 [2]);
  and (_33471_, _30990_, _06112_);
  or (_33472_, _33471_, _33470_);
  and (_33473_, _33472_, _03696_);
  or (_33474_, _33473_, _03755_);
  or (_33475_, _33474_, _33469_);
  and (_33476_, _33475_, _33457_);
  or (_33478_, _33476_, _03750_);
  or (_33479_, _33462_, _03751_);
  and (_33480_, _33479_, _03692_);
  and (_33481_, _33480_, _33478_);
  and (_33482_, _31002_, _06112_);
  or (_33483_, _33482_, _33470_);
  and (_33484_, _33483_, _03691_);
  or (_33485_, _33484_, _03684_);
  or (_33486_, _33485_, _33481_);
  and (_33487_, _33471_, _31009_);
  or (_33488_, _33470_, _03685_);
  or (_33489_, _33488_, _33487_);
  and (_33490_, _33489_, _03680_);
  and (_33491_, _33490_, _33486_);
  and (_33492_, _31016_, _06112_);
  or (_33493_, _33492_, _33470_);
  and (_33494_, _33493_, _03679_);
  or (_33495_, _33494_, _07544_);
  or (_33496_, _33495_, _33491_);
  and (_33497_, _33496_, _33456_);
  or (_33499_, _33497_, _04678_);
  and (_33500_, _06938_, _05376_);
  or (_33501_, _33452_, _04679_);
  or (_33502_, _33501_, _33500_);
  and (_33503_, _33502_, _03415_);
  and (_33504_, _33503_, _33499_);
  and (_33505_, _31041_, _05376_);
  or (_33506_, _33452_, _33505_);
  and (_33507_, _33506_, _07559_);
  or (_33508_, _33507_, _33504_);
  or (_33510_, _33508_, _08854_);
  and (_33511_, _31050_, _05376_);
  or (_33512_, _33452_, _04703_);
  or (_33513_, _33512_, _33511_);
  and (_33514_, _05376_, _06457_);
  or (_33515_, _33514_, _33452_);
  or (_33516_, _33515_, _04694_);
  and (_33517_, _33516_, _04701_);
  and (_33518_, _33517_, _33513_);
  and (_33519_, _33518_, _33510_);
  and (_33521_, _31063_, _05376_);
  or (_33522_, _33521_, _33452_);
  and (_33523_, _33522_, _03959_);
  or (_33524_, _33523_, _33519_);
  and (_33525_, _33524_, _04708_);
  or (_33526_, _33452_, _11194_);
  and (_33527_, _33515_, _03866_);
  and (_33528_, _33527_, _33526_);
  or (_33529_, _33528_, _33525_);
  and (_33530_, _33529_, _04706_);
  and (_33532_, _33462_, _03967_);
  and (_33533_, _33532_, _33526_);
  or (_33534_, _33533_, _03835_);
  or (_33535_, _33534_, _33530_);
  and (_33536_, _31047_, _05376_);
  or (_33537_, _33452_, _06532_);
  or (_33538_, _33537_, _33536_);
  and (_33539_, _33538_, _06537_);
  and (_33540_, _33539_, _33535_);
  and (_33541_, _31061_, _05376_);
  or (_33543_, _33541_, _33452_);
  and (_33544_, _33543_, _03954_);
  or (_33545_, _33544_, _03703_);
  or (_33546_, _33545_, _33540_);
  or (_33547_, _33459_, _03704_);
  and (_33548_, _33547_, _03385_);
  and (_33549_, _33548_, _33546_);
  and (_33550_, _33483_, _03384_);
  or (_33551_, _33550_, _03701_);
  or (_33552_, _33551_, _33549_);
  and (_33554_, _31098_, _05376_);
  or (_33555_, _33452_, _03702_);
  or (_33556_, _33555_, _33554_);
  and (_33557_, _33556_, _42908_);
  and (_33558_, _33557_, _33552_);
  nor (_33559_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_33560_, _33559_, _05330_);
  or (_43315_, _33560_, _33558_);
  nor (_33561_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_33562_, _33561_, _05330_);
  and (_33564_, _11413_, \oc8051_golden_model_1.P1 [3]);
  nor (_33565_, _11413_, _05050_);
  or (_33566_, _33565_, _33564_);
  or (_33567_, _33566_, _06994_);
  and (_33568_, _31112_, _05376_);
  or (_33569_, _33568_, _33564_);
  or (_33570_, _33569_, _04630_);
  and (_33571_, _05376_, \oc8051_golden_model_1.ACC [3]);
  or (_33572_, _33571_, _33564_);
  and (_33573_, _33572_, _04615_);
  and (_33575_, _04616_, \oc8051_golden_model_1.P1 [3]);
  or (_33576_, _33575_, _03757_);
  or (_33577_, _33576_, _33573_);
  and (_33578_, _33577_, _03697_);
  and (_33579_, _33578_, _33570_);
  and (_33580_, _11418_, \oc8051_golden_model_1.P1 [3]);
  and (_33581_, _31138_, _06112_);
  or (_33582_, _33581_, _33580_);
  and (_33583_, _33582_, _03696_);
  or (_33584_, _33583_, _03755_);
  or (_33586_, _33584_, _33579_);
  or (_33587_, _33566_, _04537_);
  and (_33588_, _33587_, _33586_);
  or (_33589_, _33588_, _03750_);
  or (_33590_, _33572_, _03751_);
  and (_33591_, _33590_, _03692_);
  and (_33592_, _33591_, _33589_);
  and (_33593_, _31151_, _06112_);
  or (_33594_, _33593_, _33580_);
  and (_33595_, _33594_, _03691_);
  or (_33597_, _33595_, _03684_);
  or (_33598_, _33597_, _33592_);
  or (_33599_, _33580_, _31158_);
  and (_33600_, _33599_, _33582_);
  or (_33601_, _33600_, _03685_);
  and (_33602_, _33601_, _03680_);
  and (_33603_, _33602_, _33598_);
  and (_33604_, _31164_, _06112_);
  or (_33605_, _33604_, _33580_);
  and (_33606_, _33605_, _03679_);
  or (_33608_, _33606_, _07544_);
  or (_33609_, _33608_, _33603_);
  and (_33610_, _33609_, _33567_);
  or (_33611_, _33610_, _04678_);
  and (_33612_, _06937_, _05376_);
  or (_33613_, _33564_, _04679_);
  or (_33614_, _33613_, _33612_);
  and (_33615_, _33614_, _03415_);
  and (_33616_, _33615_, _33611_);
  and (_33617_, _31189_, _05376_);
  or (_33619_, _33564_, _33617_);
  and (_33620_, _33619_, _07559_);
  or (_33621_, _33620_, _33616_);
  or (_33622_, _33621_, _08854_);
  and (_33623_, _31198_, _05376_);
  or (_33624_, _33564_, _04703_);
  or (_33625_, _33624_, _33623_);
  and (_33626_, _05376_, _06415_);
  or (_33627_, _33626_, _33564_);
  or (_33628_, _33627_, _04694_);
  and (_33630_, _33628_, _04701_);
  and (_33631_, _33630_, _33625_);
  and (_33632_, _33631_, _33622_);
  and (_33633_, _31211_, _05376_);
  or (_33634_, _33633_, _33564_);
  and (_33635_, _33634_, _03959_);
  or (_33636_, _33635_, _33632_);
  and (_33637_, _33636_, _04708_);
  or (_33638_, _33564_, _11193_);
  and (_33639_, _33627_, _03866_);
  and (_33641_, _33639_, _33638_);
  or (_33642_, _33641_, _33637_);
  and (_33643_, _33642_, _04706_);
  and (_33644_, _33572_, _03967_);
  and (_33645_, _33644_, _33638_);
  or (_33646_, _33645_, _03835_);
  or (_33647_, _33646_, _33643_);
  and (_33648_, _31196_, _05376_);
  or (_33649_, _33564_, _06532_);
  or (_33650_, _33649_, _33648_);
  and (_33652_, _33650_, _06537_);
  and (_33653_, _33652_, _33647_);
  and (_33654_, _31209_, _05376_);
  or (_33655_, _33654_, _33564_);
  and (_33656_, _33655_, _03954_);
  or (_33657_, _33656_, _03703_);
  or (_33658_, _33657_, _33653_);
  or (_33659_, _33569_, _03704_);
  and (_33660_, _33659_, _03385_);
  and (_33661_, _33660_, _33658_);
  and (_33663_, _33594_, _03384_);
  or (_33664_, _33663_, _03701_);
  or (_33665_, _33664_, _33661_);
  and (_33666_, _31246_, _05376_);
  or (_33667_, _33564_, _03702_);
  or (_33668_, _33667_, _33666_);
  and (_33669_, _33668_, _42908_);
  and (_33670_, _33669_, _33665_);
  or (_43316_, _33670_, _33562_);
  nor (_33671_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_33673_, _33671_, _05330_);
  and (_33674_, _11413_, \oc8051_golden_model_1.P1 [4]);
  nor (_33675_, _05898_, _11413_);
  or (_33676_, _33675_, _33674_);
  or (_33677_, _33676_, _06994_);
  and (_33678_, _11418_, \oc8051_golden_model_1.P1 [4]);
  and (_33679_, _31274_, _06112_);
  or (_33680_, _33679_, _33678_);
  and (_33681_, _33680_, _03691_);
  and (_33682_, _31280_, _05376_);
  or (_33684_, _33682_, _33674_);
  or (_33685_, _33684_, _04630_);
  and (_33686_, _05376_, \oc8051_golden_model_1.ACC [4]);
  or (_33687_, _33686_, _33674_);
  and (_33688_, _33687_, _04615_);
  and (_33689_, _04616_, \oc8051_golden_model_1.P1 [4]);
  or (_33690_, _33689_, _03757_);
  or (_33691_, _33690_, _33688_);
  and (_33692_, _33691_, _03697_);
  and (_33693_, _33692_, _33685_);
  and (_33695_, _31293_, _06112_);
  or (_33696_, _33695_, _33678_);
  and (_33697_, _33696_, _03696_);
  or (_33698_, _33697_, _03755_);
  or (_33699_, _33698_, _33693_);
  or (_33700_, _33676_, _04537_);
  and (_33701_, _33700_, _33699_);
  or (_33702_, _33701_, _03750_);
  or (_33703_, _33687_, _03751_);
  and (_33704_, _33703_, _03692_);
  and (_33706_, _33704_, _33702_);
  or (_33707_, _33706_, _33681_);
  and (_33708_, _33707_, _03685_);
  or (_33709_, _33678_, _31308_);
  and (_33710_, _33696_, _03684_);
  and (_33711_, _33710_, _33709_);
  or (_33712_, _33711_, _33708_);
  and (_33713_, _33712_, _03680_);
  and (_33714_, _31315_, _06112_);
  or (_33715_, _33714_, _33678_);
  and (_33717_, _33715_, _03679_);
  or (_33718_, _33717_, _07544_);
  or (_33719_, _33718_, _33713_);
  and (_33720_, _33719_, _33677_);
  or (_33721_, _33720_, _04678_);
  and (_33722_, _06942_, _05376_);
  or (_33723_, _33674_, _04679_);
  or (_33724_, _33723_, _33722_);
  and (_33725_, _33724_, _03415_);
  and (_33726_, _33725_, _33721_);
  and (_33728_, _31340_, _05376_);
  or (_33729_, _33728_, _33674_);
  and (_33730_, _33729_, _07559_);
  or (_33731_, _33730_, _08854_);
  or (_33732_, _33731_, _33726_);
  and (_33733_, _31349_, _05376_);
  or (_33734_, _33674_, _04703_);
  or (_33735_, _33734_, _33733_);
  and (_33736_, _06422_, _05376_);
  or (_33737_, _33736_, _33674_);
  or (_33739_, _33737_, _04694_);
  and (_33740_, _33739_, _04701_);
  and (_33741_, _33740_, _33735_);
  and (_33742_, _33741_, _33732_);
  and (_33743_, _31362_, _05376_);
  or (_33744_, _33743_, _33674_);
  and (_33745_, _33744_, _03959_);
  or (_33746_, _33745_, _33742_);
  and (_33747_, _33746_, _04708_);
  or (_33748_, _33674_, _11192_);
  and (_33750_, _33737_, _03866_);
  and (_33751_, _33750_, _33748_);
  or (_33752_, _33751_, _33747_);
  and (_33753_, _33752_, _04706_);
  and (_33754_, _33687_, _03967_);
  and (_33755_, _33754_, _33748_);
  or (_33756_, _33755_, _03835_);
  or (_33757_, _33756_, _33753_);
  and (_33758_, _31347_, _05376_);
  or (_33759_, _33674_, _06532_);
  or (_33761_, _33759_, _33758_);
  and (_33762_, _33761_, _06537_);
  and (_33763_, _33762_, _33757_);
  and (_33764_, _31360_, _05376_);
  or (_33765_, _33764_, _33674_);
  and (_33766_, _33765_, _03954_);
  or (_33767_, _33766_, _03703_);
  or (_33768_, _33767_, _33763_);
  or (_33769_, _33684_, _03704_);
  and (_33770_, _33769_, _03385_);
  and (_33772_, _33770_, _33768_);
  and (_33773_, _33680_, _03384_);
  or (_33774_, _33773_, _03701_);
  or (_33775_, _33774_, _33772_);
  and (_33776_, _31398_, _05376_);
  or (_33777_, _33674_, _03702_);
  or (_33778_, _33777_, _33776_);
  and (_33779_, _33778_, _42908_);
  and (_33780_, _33779_, _33775_);
  or (_43317_, _33780_, _33673_);
  and (_33781_, _11413_, \oc8051_golden_model_1.P1 [5]);
  and (_33782_, _31409_, _05376_);
  or (_33783_, _33782_, _33781_);
  or (_33784_, _33783_, _04630_);
  and (_33785_, _05376_, \oc8051_golden_model_1.ACC [5]);
  or (_33786_, _33785_, _33781_);
  and (_33787_, _33786_, _04615_);
  and (_33788_, _04616_, \oc8051_golden_model_1.P1 [5]);
  or (_33789_, _33788_, _03757_);
  or (_33790_, _33789_, _33787_);
  and (_33793_, _33790_, _03697_);
  and (_33794_, _33793_, _33784_);
  and (_33795_, _11418_, \oc8051_golden_model_1.P1 [5]);
  and (_33796_, _31435_, _06112_);
  or (_33797_, _33796_, _33795_);
  and (_33798_, _33797_, _03696_);
  or (_33799_, _33798_, _03755_);
  or (_33800_, _33799_, _33794_);
  nor (_33801_, _05799_, _11413_);
  or (_33802_, _33801_, _33781_);
  or (_33804_, _33802_, _04537_);
  and (_33805_, _33804_, _33800_);
  or (_33806_, _33805_, _03750_);
  or (_33807_, _33786_, _03751_);
  and (_33808_, _33807_, _03692_);
  and (_33809_, _33808_, _33806_);
  and (_33810_, _31450_, _06112_);
  or (_33811_, _33810_, _33795_);
  and (_33812_, _33811_, _03691_);
  or (_33813_, _33812_, _03684_);
  or (_33815_, _33813_, _33809_);
  or (_33816_, _33795_, _31457_);
  and (_33817_, _33816_, _33797_);
  or (_33818_, _33817_, _03685_);
  and (_33819_, _33818_, _03680_);
  and (_33820_, _33819_, _33815_);
  and (_33821_, _31464_, _06112_);
  or (_33822_, _33821_, _33795_);
  and (_33823_, _33822_, _03679_);
  or (_33824_, _33823_, _07544_);
  or (_33826_, _33824_, _33820_);
  or (_33827_, _33802_, _06994_);
  and (_33828_, _33827_, _33826_);
  or (_33829_, _33828_, _04678_);
  and (_33830_, _06941_, _05376_);
  or (_33831_, _33781_, _04679_);
  or (_33832_, _33831_, _33830_);
  and (_33833_, _33832_, _03415_);
  and (_33834_, _33833_, _33829_);
  and (_33835_, _31490_, _05376_);
  or (_33837_, _33835_, _33781_);
  and (_33838_, _33837_, _07559_);
  or (_33839_, _33838_, _08854_);
  or (_33840_, _33839_, _33834_);
  and (_33841_, _31499_, _05376_);
  or (_33842_, _33781_, _04703_);
  or (_33843_, _33842_, _33841_);
  and (_33844_, _06371_, _05376_);
  or (_33845_, _33844_, _33781_);
  or (_33846_, _33845_, _04694_);
  and (_33848_, _33846_, _04701_);
  and (_33849_, _33848_, _33843_);
  and (_33850_, _33849_, _33840_);
  and (_33851_, _31512_, _05376_);
  or (_33852_, _33851_, _33781_);
  and (_33853_, _33852_, _03959_);
  or (_33854_, _33853_, _33850_);
  and (_33855_, _33854_, _04708_);
  or (_33856_, _33781_, _11191_);
  and (_33857_, _33845_, _03866_);
  and (_33859_, _33857_, _33856_);
  or (_33860_, _33859_, _33855_);
  and (_33861_, _33860_, _04706_);
  and (_33862_, _33786_, _03967_);
  and (_33863_, _33862_, _33856_);
  or (_33864_, _33863_, _03835_);
  or (_33865_, _33864_, _33861_);
  and (_33866_, _31497_, _05376_);
  or (_33867_, _33781_, _06532_);
  or (_33868_, _33867_, _33866_);
  and (_33870_, _33868_, _06537_);
  and (_33871_, _33870_, _33865_);
  and (_33872_, _31510_, _05376_);
  or (_33873_, _33872_, _33781_);
  and (_33874_, _33873_, _03954_);
  or (_33875_, _33874_, _03703_);
  or (_33876_, _33875_, _33871_);
  or (_33877_, _33783_, _03704_);
  and (_33878_, _33877_, _03385_);
  and (_33879_, _33878_, _33876_);
  and (_33881_, _33811_, _03384_);
  or (_33882_, _33881_, _03701_);
  or (_33883_, _33882_, _33879_);
  and (_33884_, _31547_, _05376_);
  or (_33885_, _33781_, _03702_);
  or (_33886_, _33885_, _33884_);
  and (_33887_, _33886_, _42908_);
  and (_33888_, _33887_, _33883_);
  nor (_33889_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_33890_, _33889_, _05330_);
  or (_43318_, _33890_, _33888_);
  and (_33892_, _11413_, \oc8051_golden_model_1.P1 [6]);
  nor (_33893_, _06013_, _11413_);
  or (_33894_, _33893_, _33892_);
  or (_33895_, _33894_, _06994_);
  and (_33896_, _11418_, \oc8051_golden_model_1.P1 [6]);
  and (_33897_, _31570_, _06112_);
  or (_33898_, _33897_, _33896_);
  and (_33899_, _33898_, _03691_);
  and (_33900_, _31576_, _05376_);
  or (_33902_, _33900_, _33892_);
  or (_33903_, _33902_, _04630_);
  and (_33904_, _05376_, \oc8051_golden_model_1.ACC [6]);
  or (_33905_, _33904_, _33892_);
  and (_33906_, _33905_, _04615_);
  and (_33907_, _04616_, \oc8051_golden_model_1.P1 [6]);
  or (_33908_, _33907_, _03757_);
  or (_33909_, _33908_, _33906_);
  and (_33910_, _33909_, _03697_);
  and (_33911_, _33910_, _33903_);
  and (_33913_, _31589_, _06112_);
  or (_33914_, _33913_, _33896_);
  and (_33915_, _33914_, _03696_);
  or (_33916_, _33915_, _03755_);
  or (_33917_, _33916_, _33911_);
  or (_33918_, _33894_, _04537_);
  and (_33919_, _33918_, _33917_);
  or (_33920_, _33919_, _03750_);
  or (_33921_, _33905_, _03751_);
  and (_33922_, _33921_, _03692_);
  and (_33924_, _33922_, _33920_);
  or (_33925_, _33924_, _33899_);
  and (_33926_, _33925_, _03685_);
  or (_33927_, _33896_, _31604_);
  and (_33928_, _33914_, _03684_);
  and (_33929_, _33928_, _33927_);
  or (_33930_, _33929_, _33926_);
  and (_33931_, _33930_, _03680_);
  and (_33932_, _31610_, _06112_);
  or (_33933_, _33932_, _33896_);
  and (_33935_, _33933_, _03679_);
  or (_33936_, _33935_, _07544_);
  or (_33937_, _33936_, _33931_);
  and (_33938_, _33937_, _33895_);
  or (_33939_, _33938_, _04678_);
  and (_33940_, _06933_, _05376_);
  or (_33941_, _33892_, _04679_);
  or (_33942_, _33941_, _33940_);
  and (_33943_, _33942_, _03415_);
  and (_33944_, _33943_, _33939_);
  and (_33946_, _31646_, _05376_);
  or (_33947_, _33946_, _33892_);
  and (_33948_, _33947_, _07559_);
  or (_33949_, _33948_, _08854_);
  or (_33950_, _33949_, _33944_);
  and (_33951_, _31655_, _05376_);
  or (_33952_, _33892_, _04703_);
  or (_33953_, _33952_, _33951_);
  and (_33954_, _13333_, _05376_);
  or (_33955_, _33954_, _33892_);
  or (_33957_, _33955_, _04694_);
  and (_33958_, _33957_, _04701_);
  and (_33959_, _33958_, _33953_);
  and (_33960_, _33959_, _33950_);
  and (_33961_, _31668_, _05376_);
  or (_33962_, _33961_, _33892_);
  and (_33963_, _33962_, _03959_);
  or (_33964_, _33963_, _33960_);
  and (_33965_, _33964_, _04708_);
  or (_33966_, _33892_, _11190_);
  and (_33968_, _33955_, _03866_);
  and (_33969_, _33968_, _33966_);
  or (_33970_, _33969_, _33965_);
  and (_33971_, _33970_, _04706_);
  and (_33972_, _33905_, _03967_);
  and (_33973_, _33972_, _33966_);
  or (_33974_, _33973_, _03835_);
  or (_33975_, _33974_, _33971_);
  and (_33976_, _31653_, _05376_);
  or (_33977_, _33892_, _06532_);
  or (_33979_, _33977_, _33976_);
  and (_33980_, _33979_, _06537_);
  and (_33981_, _33980_, _33975_);
  and (_33982_, _31666_, _05376_);
  or (_33983_, _33982_, _33892_);
  and (_33984_, _33983_, _03954_);
  or (_33985_, _33984_, _03703_);
  or (_33986_, _33985_, _33981_);
  or (_33987_, _33902_, _03704_);
  and (_33988_, _33987_, _03385_);
  and (_33990_, _33988_, _33986_);
  and (_33991_, _33898_, _03384_);
  or (_33992_, _33991_, _03701_);
  or (_33993_, _33992_, _33990_);
  and (_33994_, _31704_, _05376_);
  or (_33995_, _33892_, _03702_);
  or (_33996_, _33995_, _33994_);
  and (_33997_, _33996_, _42908_);
  and (_33998_, _33997_, _33993_);
  nor (_33999_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_34001_, _33999_, _05330_);
  or (_43319_, _34001_, _33998_);
  nor (_34002_, _05434_, _03674_);
  nor (_34003_, _05652_, _11529_);
  or (_34004_, _34003_, _34002_);
  or (_34005_, _34004_, _04630_);
  and (_34006_, _05434_, \oc8051_golden_model_1.ACC [0]);
  or (_34007_, _34006_, _34002_);
  and (_34008_, _34007_, _04615_);
  nor (_34009_, _04615_, _03674_);
  or (_34011_, _34009_, _03757_);
  or (_34012_, _34011_, _34008_);
  and (_34013_, _34012_, _04537_);
  and (_34014_, _34013_, _34005_);
  or (_34015_, _34014_, _04246_);
  or (_34016_, _34007_, _03751_);
  and (_34017_, _34016_, _04759_);
  and (_34018_, _34017_, _34015_);
  nand (_34019_, _06994_, _04655_);
  or (_34020_, _34019_, _34018_);
  and (_34022_, _05434_, _04608_);
  or (_34023_, _34002_, _06994_);
  or (_34024_, _34023_, _34022_);
  and (_34025_, _34024_, _34020_);
  or (_34026_, _34025_, _04678_);
  and (_34027_, _06935_, _05434_);
  or (_34028_, _34002_, _04679_);
  or (_34029_, _34028_, _34027_);
  and (_34030_, _34029_, _34026_);
  or (_34031_, _34030_, _07559_);
  nor (_34033_, _12119_, _11529_);
  or (_34034_, _34002_, _03415_);
  or (_34035_, _34034_, _34033_);
  and (_34036_, _34035_, _04694_);
  and (_34037_, _34036_, _34031_);
  and (_34038_, _05434_, _06428_);
  or (_34039_, _34038_, _34002_);
  and (_34040_, _34039_, _03839_);
  or (_34041_, _34040_, _03838_);
  or (_34042_, _34041_, _34037_);
  and (_34044_, _12133_, _05434_);
  or (_34045_, _34002_, _04703_);
  or (_34046_, _34045_, _34044_);
  and (_34047_, _34046_, _04701_);
  and (_34048_, _34047_, _34042_);
  nor (_34049_, _10458_, _11529_);
  or (_34050_, _34049_, _34002_);
  nand (_34051_, _08712_, _05434_);
  and (_34052_, _34051_, _03959_);
  and (_34053_, _34052_, _34050_);
  or (_34054_, _34053_, _34048_);
  and (_34055_, _34054_, _04708_);
  nand (_34056_, _34039_, _03866_);
  nor (_34057_, _34056_, _34003_);
  or (_34058_, _34057_, _03967_);
  or (_34059_, _34058_, _34055_);
  nor (_34060_, _34002_, _04706_);
  nand (_34061_, _34060_, _34051_);
  and (_34062_, _34061_, _34059_);
  or (_34063_, _34062_, _03835_);
  nor (_34066_, _12132_, _11529_);
  or (_34067_, _34002_, _06532_);
  or (_34068_, _34067_, _34066_);
  and (_34069_, _34068_, _06537_);
  and (_34070_, _34069_, _34063_);
  and (_34071_, _34050_, _03954_);
  or (_34072_, _34071_, _17066_);
  or (_34073_, _34072_, _34070_);
  or (_34074_, _34004_, _04170_);
  and (_34075_, _34074_, _42908_);
  and (_34077_, _34075_, _34073_);
  nor (_34078_, _42908_, _03674_);
  or (_34079_, _34078_, rst);
  or (_43322_, _34079_, _34077_);
  nor (_34080_, _05434_, _04536_);
  and (_34081_, _12225_, _05434_);
  or (_34082_, _34081_, _34080_);
  and (_34083_, _34082_, _03701_);
  nand (_34084_, _03974_, \oc8051_golden_model_1.SP [1]);
  nand (_34085_, _04755_, _03755_);
  not (_34087_, _34081_);
  or (_34088_, _05434_, \oc8051_golden_model_1.SP [1]);
  and (_34089_, _34088_, _34087_);
  or (_34090_, _34089_, _04630_);
  nand (_34091_, _04111_, \oc8051_golden_model_1.SP [1]);
  and (_34092_, _05434_, \oc8051_golden_model_1.ACC [1]);
  or (_34093_, _34092_, _34080_);
  and (_34094_, _34093_, _04615_);
  nor (_34095_, _04615_, _04536_);
  or (_34096_, _34095_, _04111_);
  or (_34098_, _34096_, _34094_);
  and (_34099_, _34098_, _34091_);
  or (_34100_, _34099_, _03757_);
  and (_34101_, _34100_, _03445_);
  and (_34102_, _34101_, _34090_);
  nor (_34103_, _03445_, \oc8051_golden_model_1.SP [1]);
  or (_34104_, _34103_, _03755_);
  or (_34105_, _34104_, _34102_);
  and (_34106_, _34105_, _34085_);
  or (_34107_, _34106_, _03750_);
  or (_34109_, _34093_, _03751_);
  and (_34110_, _34109_, _04759_);
  and (_34111_, _34110_, _34107_);
  not (_34112_, _04968_);
  or (_34113_, _34112_, _04851_);
  or (_34114_, _34113_, _34111_);
  or (_34115_, _04968_, _04536_);
  and (_34116_, _34115_, _06994_);
  and (_34117_, _34116_, _34114_);
  or (_34118_, _11529_, _04813_);
  and (_34120_, _34088_, _07544_);
  and (_34121_, _34120_, _34118_);
  or (_34122_, _34121_, _04678_);
  or (_34123_, _34122_, _34117_);
  and (_34124_, _06934_, _05434_);
  or (_34125_, _34080_, _04679_);
  or (_34126_, _34125_, _34124_);
  and (_34127_, _34126_, _03415_);
  and (_34128_, _34127_, _34123_);
  nor (_34129_, _12313_, _11529_);
  or (_34131_, _34129_, _34080_);
  and (_34132_, _34131_, _07559_);
  or (_34133_, _34132_, _34128_);
  and (_34134_, _34133_, _04694_);
  nand (_34135_, _05434_, _04515_);
  and (_34136_, _34088_, _03839_);
  and (_34137_, _34136_, _34135_);
  or (_34138_, _34137_, _03483_);
  or (_34139_, _34138_, _34134_);
  and (_34140_, _03483_, \oc8051_golden_model_1.SP [1]);
  nor (_34142_, _34140_, _03838_);
  and (_34143_, _34142_, _34139_);
  or (_34144_, _12207_, _11529_);
  and (_34145_, _34088_, _03838_);
  and (_34146_, _34145_, _34144_);
  or (_34147_, _34146_, _03959_);
  or (_34148_, _34147_, _34143_);
  nor (_34149_, _08710_, _11529_);
  or (_34150_, _34149_, _34080_);
  nand (_34151_, _08709_, _05434_);
  and (_34153_, _34151_, _34150_);
  or (_34154_, _34153_, _04701_);
  and (_34155_, _34154_, _04708_);
  and (_34156_, _34155_, _34148_);
  or (_34157_, _12206_, _11529_);
  and (_34158_, _34088_, _03866_);
  and (_34159_, _34158_, _34157_);
  or (_34160_, _34159_, _03967_);
  or (_34161_, _34160_, _34156_);
  nor (_34162_, _34080_, _04706_);
  nand (_34164_, _34162_, _34151_);
  and (_34165_, _34164_, _34161_);
  or (_34166_, _34165_, _03477_);
  and (_34167_, _03477_, \oc8051_golden_model_1.SP [1]);
  nor (_34168_, _34167_, _03835_);
  and (_34169_, _34168_, _34166_);
  or (_34170_, _34135_, _05603_);
  and (_34171_, _34088_, _03835_);
  and (_34172_, _34171_, _34170_);
  or (_34173_, _34172_, _34169_);
  and (_34175_, _34173_, _06537_);
  and (_34176_, _34150_, _03954_);
  or (_34177_, _34176_, _03974_);
  or (_34178_, _34177_, _34175_);
  nand (_34179_, _34178_, _34084_);
  nor (_34180_, _03707_, _03474_);
  nand (_34181_, _34180_, _34179_);
  or (_34182_, _34180_, _04536_);
  and (_34183_, _34182_, _03704_);
  and (_34184_, _34183_, _34181_);
  and (_34186_, _34089_, _03703_);
  or (_34187_, _34186_, _05156_);
  or (_34188_, _34187_, _34184_);
  or (_34189_, _04735_, _04536_);
  and (_34190_, _34189_, _03702_);
  and (_34191_, _34190_, _34188_);
  or (_34192_, _34191_, _34083_);
  and (_34193_, _34192_, _42908_);
  nor (_34194_, \oc8051_golden_model_1.SP [1], rst);
  nor (_34195_, _34194_, _00000_);
  or (_43323_, _34195_, _34193_);
  nor (_34197_, \oc8051_golden_model_1.SP [2], rst);
  nor (_34198_, _34197_, _00000_);
  nor (_34199_, _11529_, _05236_);
  nor (_34200_, _05434_, _04125_);
  or (_34201_, _34200_, _06994_);
  or (_34202_, _34201_, _34199_);
  or (_34203_, _05268_, _05105_);
  nand (_34204_, _06168_, _03755_);
  nor (_34205_, _12427_, _11529_);
  or (_34207_, _34205_, _34200_);
  or (_34208_, _34207_, _04630_);
  and (_34209_, _05434_, \oc8051_golden_model_1.ACC [2]);
  or (_34210_, _34209_, _34200_);
  or (_34211_, _34210_, _04616_);
  or (_34212_, _04615_, \oc8051_golden_model_1.SP [2]);
  and (_34213_, _34212_, _04948_);
  and (_34214_, _34213_, _34211_);
  and (_34215_, _05326_, _04111_);
  or (_34216_, _34215_, _03757_);
  or (_34217_, _34216_, _34214_);
  and (_34218_, _34217_, _03445_);
  and (_34219_, _34218_, _34208_);
  nor (_34220_, _13785_, _03445_);
  or (_34221_, _34220_, _03755_);
  or (_34222_, _34221_, _34219_);
  and (_34223_, _34222_, _34204_);
  or (_34224_, _34223_, _03750_);
  or (_34225_, _34210_, _03751_);
  and (_34226_, _34225_, _04759_);
  and (_34228_, _34226_, _34224_);
  or (_34229_, _34228_, _34203_);
  or (_34230_, _05326_, _03442_);
  and (_34231_, _34230_, _03418_);
  and (_34232_, _34231_, _34229_);
  or (_34233_, _13785_, _03418_);
  nand (_34234_, _34233_, _06994_);
  or (_34235_, _34234_, _34232_);
  and (_34236_, _34235_, _34202_);
  or (_34237_, _34236_, _04678_);
  and (_34239_, _06938_, _05434_);
  or (_34240_, _34239_, _34200_);
  or (_34241_, _34240_, _04679_);
  and (_34242_, _34241_, _34237_);
  or (_34243_, _34242_, _07559_);
  nor (_34244_, _12523_, _11529_);
  or (_34245_, _34200_, _03415_);
  or (_34246_, _34245_, _34244_);
  and (_34247_, _34246_, _04694_);
  and (_34248_, _34247_, _34243_);
  and (_34250_, _05434_, _06457_);
  or (_34251_, _34250_, _34200_);
  and (_34252_, _34251_, _03839_);
  or (_34253_, _34252_, _03483_);
  or (_34254_, _34253_, _34248_);
  nand (_34255_, _13785_, _03483_);
  and (_34256_, _34255_, _34254_);
  or (_34257_, _34256_, _03838_);
  and (_34258_, _12537_, _05434_);
  or (_34259_, _34200_, _04703_);
  or (_34261_, _34259_, _34258_);
  and (_34262_, _34261_, _04701_);
  and (_34263_, _34262_, _34257_);
  and (_34264_, _08707_, _05434_);
  or (_34265_, _34264_, _34200_);
  and (_34266_, _34265_, _03959_);
  or (_34267_, _34266_, _34263_);
  and (_34268_, _34267_, _04708_);
  or (_34269_, _34200_, _05700_);
  and (_34270_, _34251_, _03866_);
  and (_34272_, _34270_, _34269_);
  or (_34273_, _34272_, _34268_);
  and (_34274_, _34273_, _10031_);
  and (_34275_, _34210_, _03967_);
  and (_34276_, _34275_, _34269_);
  and (_34277_, _05326_, _03477_);
  or (_34278_, _34277_, _03835_);
  or (_34279_, _34278_, _34276_);
  or (_34280_, _34279_, _34274_);
  nor (_34281_, _12536_, _11529_);
  or (_34283_, _34200_, _06532_);
  or (_34284_, _34283_, _34281_);
  and (_34285_, _34284_, _34280_);
  or (_34286_, _34285_, _03954_);
  nor (_34287_, _08706_, _11529_);
  or (_34288_, _34287_, _34200_);
  or (_34289_, _34288_, _06537_);
  and (_34290_, _34289_, _11621_);
  and (_34291_, _34290_, _34286_);
  and (_34292_, _13785_, _03974_);
  or (_34294_, _34292_, _03474_);
  or (_34295_, _34294_, _34291_);
  nand (_34296_, _13785_, _03474_);
  and (_34297_, _34296_, _03708_);
  and (_34298_, _34297_, _34295_);
  and (_34299_, _13785_, _03707_);
  or (_34300_, _34299_, _03703_);
  or (_34301_, _34300_, _34298_);
  or (_34302_, _34207_, _03704_);
  and (_34303_, _34302_, _04735_);
  and (_34305_, _34303_, _34301_);
  nor (_34306_, _13785_, _04735_);
  or (_34307_, _34306_, _03701_);
  or (_34308_, _34307_, _34305_);
  and (_34309_, _12596_, _05434_);
  or (_34310_, _34200_, _03702_);
  or (_34311_, _34310_, _34309_);
  and (_34312_, _34311_, _42908_);
  and (_34313_, _34312_, _34308_);
  or (_43324_, _34313_, _34198_);
  nor (_34315_, _42908_, _03754_);
  or (_34316_, _05329_, _04735_);
  nand (_34317_, _13579_, _03474_);
  nand (_34318_, _13579_, _03483_);
  nor (_34319_, _11529_, _05050_);
  nor (_34320_, _05434_, _03754_);
  or (_34321_, _34320_, _04678_);
  or (_34322_, _34321_, _34319_);
  and (_34323_, _34322_, _11528_);
  nor (_34324_, _12610_, _11529_);
  or (_34326_, _34324_, _34320_);
  or (_34327_, _34326_, _04630_);
  and (_34328_, _05434_, \oc8051_golden_model_1.ACC [3]);
  or (_34329_, _34328_, _34320_);
  or (_34330_, _34329_, _04616_);
  or (_34331_, _04615_, \oc8051_golden_model_1.SP [3]);
  and (_34332_, _34331_, _04948_);
  and (_34333_, _34332_, _34330_);
  and (_34334_, _05329_, _04111_);
  or (_34335_, _34334_, _03757_);
  or (_34337_, _34335_, _34333_);
  and (_34338_, _34337_, _03445_);
  and (_34339_, _34338_, _34327_);
  nor (_34340_, _13579_, _03445_);
  or (_34341_, _34340_, _03755_);
  or (_34342_, _34341_, _34339_);
  nand (_34343_, _06157_, _03755_);
  and (_34344_, _34343_, _34342_);
  or (_34345_, _34344_, _03750_);
  or (_34346_, _34329_, _03751_);
  and (_34348_, _34346_, _04759_);
  and (_34349_, _34348_, _34345_);
  or (_34350_, _05099_, _34112_);
  or (_34351_, _34350_, _34349_);
  or (_34352_, _05329_, _04968_);
  and (_34353_, _34352_, _06994_);
  and (_34354_, _34353_, _34351_);
  or (_34355_, _34354_, _34323_);
  and (_34356_, _06937_, _05434_);
  or (_34357_, _34320_, _04679_);
  or (_34359_, _34357_, _34356_);
  and (_34360_, _34359_, _03415_);
  and (_34361_, _34360_, _34355_);
  nor (_34362_, _12724_, _11529_);
  or (_34363_, _34362_, _34320_);
  and (_34364_, _34363_, _07559_);
  or (_34365_, _34364_, _03839_);
  or (_34366_, _34365_, _34361_);
  and (_34367_, _05434_, _06415_);
  or (_34368_, _34367_, _34320_);
  or (_34370_, _34368_, _04694_);
  and (_34371_, _34370_, _34366_);
  or (_34372_, _34371_, _03483_);
  and (_34373_, _34372_, _34318_);
  or (_34374_, _34373_, _03838_);
  and (_34375_, _12738_, _05434_);
  or (_34376_, _34320_, _04703_);
  or (_34377_, _34376_, _34375_);
  and (_34378_, _34377_, _04701_);
  and (_34379_, _34378_, _34374_);
  and (_34381_, _10455_, _05434_);
  or (_34382_, _34381_, _34320_);
  and (_34383_, _34382_, _03959_);
  or (_34384_, _34383_, _34379_);
  and (_34385_, _34384_, _04708_);
  or (_34386_, _34320_, _05554_);
  and (_34387_, _34368_, _03866_);
  and (_34388_, _34387_, _34386_);
  or (_34389_, _34388_, _34385_);
  and (_34390_, _34389_, _10031_);
  and (_34392_, _34329_, _03967_);
  and (_34393_, _34392_, _34386_);
  and (_34394_, _05329_, _03477_);
  or (_34395_, _34394_, _03835_);
  or (_34396_, _34395_, _34393_);
  or (_34397_, _34396_, _34390_);
  nor (_34398_, _12737_, _11529_);
  or (_34399_, _34398_, _34320_);
  or (_34400_, _34399_, _06532_);
  and (_34401_, _34400_, _34397_);
  or (_34403_, _34401_, _03954_);
  nor (_34404_, _08701_, _11529_);
  or (_34405_, _34404_, _34320_);
  or (_34406_, _34405_, _06537_);
  and (_34407_, _34406_, _11621_);
  and (_34408_, _34407_, _34403_);
  nor (_34409_, _06154_, _03754_);
  or (_34410_, _34409_, _06155_);
  and (_34411_, _34410_, _03974_);
  or (_34412_, _34411_, _03474_);
  or (_34414_, _34412_, _34408_);
  and (_34415_, _34414_, _34317_);
  or (_34416_, _34415_, _03707_);
  or (_34417_, _34410_, _03708_);
  and (_34418_, _34417_, _03704_);
  and (_34419_, _34418_, _34416_);
  and (_34420_, _34326_, _03703_);
  or (_34421_, _34420_, _05156_);
  or (_34422_, _34421_, _34419_);
  and (_34423_, _34422_, _34316_);
  or (_34425_, _34423_, _03701_);
  and (_34426_, _12792_, _05434_);
  or (_34427_, _34320_, _03702_);
  or (_34428_, _34427_, _34426_);
  and (_34429_, _34428_, _42908_);
  and (_34430_, _34429_, _34425_);
  or (_34431_, _34430_, _34315_);
  and (_43327_, _34431_, _41654_);
  nor (_34432_, _42908_, _11536_);
  nor (_34433_, _05059_, \oc8051_golden_model_1.SP [4]);
  nor (_34435_, _34433_, _11517_);
  or (_34436_, _34435_, _04735_);
  or (_34437_, _34435_, _06543_);
  and (_34438_, _05060_, \oc8051_golden_model_1.SP [4]);
  nor (_34439_, _05060_, \oc8051_golden_model_1.SP [4]);
  nor (_34440_, _34439_, _34438_);
  and (_34441_, _34440_, _03690_);
  and (_34442_, _11537_, _03674_);
  nor (_34443_, _06156_, _11536_);
  nor (_34444_, _34443_, _34442_);
  nand (_34446_, _34444_, _03755_);
  nor (_34447_, _05434_, _11536_);
  nor (_34448_, _12828_, _11529_);
  or (_34449_, _34448_, _34447_);
  or (_34450_, _34449_, _04630_);
  and (_34451_, _05434_, \oc8051_golden_model_1.ACC [4]);
  or (_34452_, _34451_, _34447_);
  or (_34453_, _34452_, _04616_);
  or (_34454_, _04615_, \oc8051_golden_model_1.SP [4]);
  and (_34455_, _34454_, _04948_);
  and (_34457_, _34455_, _34453_);
  and (_34458_, _34435_, _04111_);
  or (_34459_, _34458_, _03757_);
  or (_34460_, _34459_, _34457_);
  and (_34461_, _34460_, _03445_);
  and (_34462_, _34461_, _34450_);
  and (_34463_, _34435_, _04933_);
  or (_34464_, _34463_, _03755_);
  or (_34465_, _34464_, _34462_);
  and (_34466_, _34465_, _34446_);
  or (_34468_, _34466_, _03750_);
  or (_34469_, _34452_, _03751_);
  and (_34470_, _34469_, _04759_);
  and (_34471_, _34470_, _34468_);
  or (_34472_, _34471_, _34441_);
  and (_34473_, _34472_, _04968_);
  nand (_34474_, _34435_, _34112_);
  nand (_34475_, _34474_, _06994_);
  or (_34476_, _34475_, _34473_);
  nor (_34477_, _05898_, _11529_);
  or (_34479_, _34447_, _06994_);
  or (_34480_, _34479_, _34477_);
  and (_34481_, _34480_, _04679_);
  and (_34482_, _34481_, _34476_);
  and (_34483_, _06942_, _05434_);
  or (_34484_, _34483_, _34447_);
  and (_34485_, _34484_, _04678_);
  or (_34486_, _34485_, _07559_);
  or (_34487_, _34486_, _34482_);
  nor (_34488_, _12919_, _11529_);
  or (_34490_, _34488_, _34447_);
  or (_34491_, _34490_, _03415_);
  and (_34492_, _34491_, _34487_);
  or (_34493_, _34492_, _03839_);
  and (_34494_, _06422_, _05434_);
  or (_34495_, _34494_, _34447_);
  or (_34496_, _34495_, _04694_);
  and (_34497_, _34496_, _11594_);
  and (_34498_, _34497_, _34493_);
  and (_34499_, _34435_, _03483_);
  or (_34501_, _34499_, _03838_);
  or (_34502_, _34501_, _34498_);
  and (_34503_, _12933_, _05434_);
  or (_34504_, _34447_, _04703_);
  or (_34505_, _34504_, _34503_);
  and (_34506_, _34505_, _04701_);
  and (_34507_, _34506_, _34502_);
  and (_34508_, _08700_, _05434_);
  or (_34509_, _34508_, _34447_);
  and (_34510_, _34509_, _03959_);
  or (_34512_, _34510_, _34507_);
  and (_34513_, _34512_, _04708_);
  or (_34514_, _34447_, _08303_);
  and (_34515_, _34495_, _03866_);
  and (_34516_, _34515_, _34514_);
  or (_34517_, _34516_, _34513_);
  and (_34518_, _34517_, _10031_);
  and (_34519_, _34452_, _03967_);
  and (_34520_, _34519_, _34514_);
  and (_34521_, _34435_, _03477_);
  or (_34523_, _34521_, _03835_);
  or (_34524_, _34523_, _34520_);
  or (_34525_, _34524_, _34518_);
  nor (_34526_, _12931_, _11529_);
  or (_34527_, _34447_, _06532_);
  or (_34528_, _34527_, _34526_);
  and (_34529_, _34528_, _34525_);
  or (_34530_, _34529_, _03954_);
  nor (_34531_, _08699_, _11529_);
  or (_34532_, _34531_, _34447_);
  or (_34534_, _34532_, _06537_);
  and (_34535_, _34534_, _11621_);
  and (_34536_, _34535_, _34530_);
  nor (_34537_, _06155_, _11536_);
  or (_34538_, _34537_, _11537_);
  and (_34539_, _34538_, _03974_);
  or (_34540_, _34539_, _03474_);
  or (_34541_, _34540_, _34536_);
  and (_34542_, _34541_, _34437_);
  or (_34543_, _34542_, _03707_);
  or (_34545_, _34538_, _03708_);
  and (_34546_, _34545_, _03704_);
  and (_34547_, _34546_, _34543_);
  and (_34548_, _34449_, _03703_);
  or (_34549_, _34548_, _05156_);
  or (_34550_, _34549_, _34547_);
  and (_34551_, _34550_, _34436_);
  or (_34552_, _34551_, _03701_);
  and (_34553_, _12991_, _05434_);
  or (_34554_, _34447_, _03702_);
  or (_34556_, _34554_, _34553_);
  and (_34557_, _34556_, _42908_);
  and (_34558_, _34557_, _34552_);
  or (_34559_, _34558_, _34432_);
  and (_43328_, _34559_, _41654_);
  nor (_34560_, _42908_, _11535_);
  nor (_34561_, _11517_, \oc8051_golden_model_1.SP [5]);
  nor (_34562_, _34561_, _11518_);
  or (_34563_, _34562_, _04735_);
  or (_34564_, _34562_, _06543_);
  nor (_34566_, _05799_, _11529_);
  nor (_34567_, _05434_, _11535_);
  or (_34568_, _34567_, _06994_);
  or (_34569_, _34568_, _34566_);
  nor (_34570_, _13025_, _11529_);
  or (_34571_, _34570_, _34567_);
  or (_34572_, _34571_, _04630_);
  and (_34573_, _05434_, \oc8051_golden_model_1.ACC [5]);
  or (_34574_, _34573_, _34567_);
  or (_34575_, _34574_, _04616_);
  or (_34577_, _04615_, \oc8051_golden_model_1.SP [5]);
  and (_34578_, _34577_, _04948_);
  and (_34579_, _34578_, _34575_);
  and (_34580_, _34562_, _04111_);
  or (_34581_, _34580_, _03757_);
  or (_34582_, _34581_, _34579_);
  and (_34583_, _34582_, _03445_);
  and (_34584_, _34583_, _34572_);
  and (_34585_, _34562_, _04933_);
  or (_34586_, _34585_, _03755_);
  or (_34588_, _34586_, _34584_);
  and (_34589_, _11538_, _03674_);
  nor (_34590_, _34442_, _11535_);
  nor (_34591_, _34590_, _34589_);
  nand (_34592_, _34591_, _03755_);
  and (_34593_, _34592_, _34588_);
  or (_34594_, _34593_, _03750_);
  or (_34595_, _34574_, _03751_);
  and (_34596_, _34595_, _04759_);
  and (_34597_, _34596_, _34594_);
  nor (_34599_, _34438_, \oc8051_golden_model_1.SP [5]);
  nor (_34600_, _34599_, _11567_);
  and (_34601_, _34600_, _03690_);
  or (_34602_, _34601_, _34597_);
  and (_34603_, _34602_, _04968_);
  nand (_34604_, _34562_, _34112_);
  nand (_34605_, _34604_, _06994_);
  or (_34606_, _34605_, _34603_);
  and (_34607_, _34606_, _34569_);
  or (_34608_, _34607_, _04678_);
  and (_34610_, _06941_, _05434_);
  or (_34611_, _34567_, _04679_);
  or (_34612_, _34611_, _34610_);
  and (_34613_, _34612_, _34608_);
  or (_34614_, _34613_, _07559_);
  nor (_34615_, _13118_, _11529_);
  or (_34616_, _34615_, _34567_);
  or (_34617_, _34616_, _03415_);
  and (_34618_, _34617_, _34614_);
  or (_34619_, _34618_, _03839_);
  and (_34621_, _06371_, _05434_);
  or (_34622_, _34621_, _34567_);
  or (_34623_, _34622_, _04694_);
  and (_34624_, _34623_, _11594_);
  and (_34625_, _34624_, _34619_);
  and (_34626_, _34562_, _03483_);
  or (_34627_, _34626_, _03838_);
  or (_34628_, _34627_, _34625_);
  and (_34629_, _13133_, _05434_);
  or (_34630_, _34567_, _04703_);
  or (_34632_, _34630_, _34629_);
  and (_34633_, _34632_, _04701_);
  and (_34634_, _34633_, _34628_);
  and (_34635_, _10451_, _05434_);
  or (_34636_, _34635_, _34567_);
  and (_34637_, _34636_, _03959_);
  or (_34638_, _34637_, _34634_);
  and (_34639_, _34638_, _04708_);
  or (_34640_, _34567_, _08302_);
  and (_34641_, _34622_, _03866_);
  and (_34643_, _34641_, _34640_);
  or (_34644_, _34643_, _34639_);
  and (_34645_, _34644_, _10031_);
  and (_34646_, _34574_, _03967_);
  and (_34647_, _34646_, _34640_);
  and (_34648_, _34562_, _03477_);
  or (_34649_, _34648_, _03835_);
  or (_34650_, _34649_, _34647_);
  or (_34651_, _34650_, _34645_);
  nor (_34652_, _13131_, _11529_);
  or (_34654_, _34567_, _06532_);
  or (_34655_, _34654_, _34652_);
  and (_34656_, _34655_, _34651_);
  or (_34657_, _34656_, _03954_);
  nor (_34658_, _08697_, _11529_);
  or (_34659_, _34658_, _34567_);
  or (_34660_, _34659_, _06537_);
  and (_34661_, _34660_, _11621_);
  and (_34662_, _34661_, _34657_);
  nor (_34663_, _11537_, _11535_);
  or (_34665_, _34663_, _11538_);
  and (_34666_, _34665_, _03974_);
  or (_34667_, _34666_, _03474_);
  or (_34668_, _34667_, _34662_);
  and (_34669_, _34668_, _34564_);
  or (_34670_, _34669_, _03707_);
  or (_34671_, _34665_, _03708_);
  and (_34672_, _34671_, _03704_);
  and (_34673_, _34672_, _34670_);
  and (_34674_, _34571_, _03703_);
  or (_34675_, _34674_, _05156_);
  or (_34676_, _34675_, _34673_);
  and (_34677_, _34676_, _34563_);
  or (_34678_, _34677_, _03701_);
  and (_34679_, _13193_, _05434_);
  or (_34680_, _34567_, _03702_);
  or (_34681_, _34680_, _34679_);
  and (_34682_, _34681_, _42908_);
  and (_34683_, _34682_, _34678_);
  or (_34684_, _34683_, _34560_);
  and (_43329_, _34684_, _41654_);
  nor (_34687_, _42908_, _11534_);
  nor (_34688_, _06013_, _11529_);
  nor (_34689_, _05434_, _11534_);
  or (_34690_, _34689_, _06994_);
  or (_34691_, _34690_, _34688_);
  nor (_34692_, _34589_, _11534_);
  nor (_34693_, _34692_, _11540_);
  nand (_34694_, _34693_, _03755_);
  nor (_34695_, _13234_, _11529_);
  or (_34697_, _34695_, _34689_);
  or (_34698_, _34697_, _04630_);
  and (_34699_, _05434_, \oc8051_golden_model_1.ACC [6]);
  or (_34700_, _34699_, _34689_);
  or (_34701_, _34700_, _04616_);
  or (_34702_, _04615_, \oc8051_golden_model_1.SP [6]);
  and (_34703_, _34702_, _04948_);
  and (_34704_, _34703_, _34701_);
  nor (_34705_, _11518_, \oc8051_golden_model_1.SP [6]);
  nor (_34706_, _34705_, _11519_);
  and (_34708_, _34706_, _04111_);
  or (_34709_, _34708_, _03757_);
  or (_34710_, _34709_, _34704_);
  and (_34711_, _34710_, _03445_);
  and (_34712_, _34711_, _34698_);
  and (_34713_, _34706_, _04933_);
  or (_34714_, _34713_, _03755_);
  or (_34715_, _34714_, _34712_);
  and (_34716_, _34715_, _34694_);
  or (_34717_, _34716_, _03750_);
  or (_34719_, _34700_, _03751_);
  and (_34720_, _34719_, _04759_);
  and (_34721_, _34720_, _34717_);
  nor (_34722_, _11567_, \oc8051_golden_model_1.SP [6]);
  nor (_34723_, _34722_, _11568_);
  and (_34724_, _34723_, _03690_);
  or (_34725_, _34724_, _34721_);
  and (_34726_, _34725_, _04968_);
  nand (_34727_, _34706_, _34112_);
  nand (_34728_, _34727_, _06994_);
  or (_34730_, _34728_, _34726_);
  and (_34731_, _34730_, _34691_);
  or (_34732_, _34731_, _04678_);
  and (_34733_, _06933_, _05434_);
  or (_34734_, _34689_, _04679_);
  or (_34735_, _34734_, _34733_);
  and (_34736_, _34735_, _03415_);
  and (_34737_, _34736_, _34732_);
  nor (_34738_, _13326_, _11529_);
  or (_34739_, _34738_, _34689_);
  and (_34741_, _34739_, _07559_);
  or (_34742_, _34741_, _03839_);
  or (_34743_, _34742_, _34737_);
  and (_34744_, _13333_, _05434_);
  or (_34745_, _34744_, _34689_);
  or (_34746_, _34745_, _04694_);
  and (_34747_, _34746_, _34743_);
  or (_34748_, _34747_, _03483_);
  or (_34749_, _34706_, _11594_);
  and (_34750_, _34749_, _34748_);
  or (_34752_, _34750_, _03838_);
  and (_34753_, _13341_, _05434_);
  or (_34754_, _34753_, _34689_);
  or (_34755_, _34754_, _04703_);
  and (_34756_, _34755_, _04701_);
  and (_34757_, _34756_, _34752_);
  and (_34758_, _08695_, _05434_);
  or (_34759_, _34758_, _34689_);
  and (_34760_, _34759_, _03959_);
  or (_34761_, _34760_, _34757_);
  and (_34763_, _34761_, _04708_);
  or (_34764_, _34689_, _08289_);
  and (_34765_, _34745_, _03866_);
  and (_34766_, _34765_, _34764_);
  or (_34767_, _34766_, _34763_);
  and (_34768_, _34767_, _10031_);
  and (_34769_, _34700_, _03967_);
  and (_34770_, _34769_, _34764_);
  and (_34771_, _34706_, _03477_);
  or (_34772_, _34771_, _03835_);
  or (_34774_, _34772_, _34770_);
  or (_34775_, _34774_, _34768_);
  nor (_34776_, _13340_, _11529_);
  or (_34777_, _34689_, _06532_);
  or (_34778_, _34777_, _34776_);
  and (_34779_, _34778_, _34775_);
  or (_34780_, _34779_, _03954_);
  nor (_34781_, _08694_, _11529_);
  or (_34782_, _34781_, _34689_);
  or (_34783_, _34782_, _06537_);
  and (_34785_, _34783_, _11621_);
  and (_34786_, _34785_, _34780_);
  nor (_34787_, _11538_, _11534_);
  or (_34788_, _34787_, _11539_);
  and (_34789_, _34788_, _03974_);
  or (_34790_, _34789_, _03474_);
  or (_34791_, _34790_, _34786_);
  or (_34792_, _34706_, _06543_);
  and (_34793_, _34792_, _03708_);
  and (_34794_, _34793_, _34791_);
  and (_34796_, _34788_, _03707_);
  or (_34797_, _34796_, _03703_);
  or (_34798_, _34797_, _34794_);
  or (_34799_, _34697_, _03704_);
  and (_34800_, _34799_, _04735_);
  and (_34801_, _34800_, _34798_);
  and (_34802_, _34706_, _05156_);
  or (_34803_, _34802_, _03701_);
  or (_34804_, _34803_, _34801_);
  nor (_34805_, _13399_, _11529_);
  or (_34807_, _34689_, _03702_);
  or (_34808_, _34807_, _34805_);
  and (_34809_, _34808_, _42908_);
  and (_34810_, _34809_, _34804_);
  or (_34811_, _34810_, _34687_);
  and (_43330_, _34811_, _41654_);
  not (_34812_, \oc8051_golden_model_1.PSW [0]);
  nor (_34813_, _42908_, _34812_);
  nor (_34814_, _07681_, _07680_);
  nor (_34815_, _34814_, _07586_);
  and (_34817_, _34814_, _07586_);
  nor (_34818_, _34817_, _34815_);
  nor (_34819_, _07605_, _07603_);
  nor (_34820_, _34819_, _15422_);
  and (_34821_, _34819_, _15422_);
  nor (_34822_, _34821_, _34820_);
  and (_34823_, _34822_, _34818_);
  nor (_34824_, _34822_, _34818_);
  nor (_34825_, _34824_, _34823_);
  or (_34826_, _34825_, _06142_);
  nand (_34828_, _34825_, _06142_);
  and (_34829_, _34828_, _34826_);
  and (_34830_, _34829_, _12199_);
  or (_34831_, _34829_, _04735_);
  and (_34832_, _12353_, _03473_);
  not (_34833_, _34832_);
  not (_34834_, _15767_);
  nor (_34835_, _15020_, _08554_);
  not (_34836_, _15020_);
  nor (_34837_, _15381_, _34836_);
  nor (_34839_, _34837_, _34835_);
  nor (_34840_, _34839_, _15686_);
  and (_34841_, _34839_, _15686_);
  nor (_34842_, _34841_, _34840_);
  and (_34843_, _34842_, _34834_);
  nor (_34844_, _34842_, _34834_);
  nor (_34845_, _34844_, _34843_);
  and (_34846_, _34845_, _16329_);
  nor (_34847_, _34845_, _16329_);
  nor (_34848_, _34847_, _34846_);
  nor (_34850_, _34848_, _16411_);
  and (_34851_, _34848_, _16411_);
  or (_34852_, _34851_, _34850_);
  nor (_34853_, _34852_, _16986_);
  and (_34854_, _34852_, _16986_);
  or (_34855_, _34854_, _34853_);
  and (_34856_, _34855_, _08571_);
  nor (_34857_, _34855_, _08571_);
  or (_34858_, _34857_, _34856_);
  and (_34859_, _34858_, _15379_);
  nor (_34861_, _14945_, _08665_);
  and (_34862_, _14945_, _08665_);
  nor (_34863_, _34862_, _34861_);
  nor (_34864_, _08659_, _15667_);
  and (_34865_, _08659_, _15667_);
  nor (_34866_, _34865_, _34864_);
  and (_34867_, _34866_, _34863_);
  nor (_34868_, _34866_, _34863_);
  nor (_34869_, _34868_, _34867_);
  not (_34870_, _08652_);
  nor (_34872_, _08656_, _08649_);
  and (_34873_, _08656_, _08649_);
  nor (_34874_, _34873_, _34872_);
  nor (_34875_, _34874_, _34870_);
  and (_34876_, _34874_, _34870_);
  nor (_34877_, _34876_, _34875_);
  and (_34878_, _34877_, _34869_);
  nor (_34879_, _34877_, _34869_);
  or (_34880_, _34879_, _34878_);
  and (_34881_, _34880_, _08082_);
  nor (_34883_, _34880_, _08082_);
  or (_34884_, _34883_, _34881_);
  and (_34885_, _34884_, _10019_);
  and (_34886_, _03850_, _03476_);
  and (_34887_, _34829_, _29313_);
  not (_34888_, _16747_);
  and (_34889_, _34888_, _08490_);
  nor (_34890_, _34888_, _08490_);
  nor (_34891_, _34890_, _34889_);
  and (_34892_, _16420_, _16076_);
  nor (_34894_, _16420_, _16076_);
  or (_34895_, _34894_, _34892_);
  nor (_34896_, _15192_, _14956_);
  and (_34897_, _15192_, _14956_);
  nor (_34898_, _34897_, _34896_);
  nor (_34899_, _15772_, _15640_);
  and (_34900_, _15772_, _15640_);
  nor (_34901_, _34900_, _34899_);
  nor (_34902_, _34901_, _34898_);
  and (_34903_, _34901_, _34898_);
  nor (_34905_, _34903_, _34902_);
  nor (_34906_, _34905_, _34895_);
  and (_34907_, _34905_, _34895_);
  nor (_34908_, _34907_, _34906_);
  nand (_34909_, _34908_, _34891_);
  or (_34910_, _34908_, _34891_);
  and (_34911_, _34910_, _03838_);
  and (_34912_, _34911_, _34909_);
  or (_34913_, _34829_, _28600_);
  and (_34914_, _12353_, _03689_);
  not (_34916_, _34914_);
  or (_34917_, _06939_, _06790_);
  nand (_34918_, _34917_, _12197_);
  or (_34919_, _34917_, _12197_);
  nand (_34920_, _34919_, _34918_);
  nor (_34921_, _06943_, _06882_);
  or (_34922_, _06933_, _06280_);
  or (_34923_, _06607_, _06237_);
  and (_34924_, _34923_, _34922_);
  nand (_34925_, _34924_, _34921_);
  or (_34927_, _34924_, _34921_);
  nand (_34928_, _34927_, _34925_);
  nand (_34929_, _34928_, _34920_);
  or (_34930_, _34928_, _34920_);
  and (_34931_, _34930_, _34929_);
  or (_34932_, _34931_, _34916_);
  nor (_34933_, _06916_, _06132_);
  and (_34934_, _34933_, _12216_);
  nor (_34935_, _34933_, _12216_);
  or (_34936_, _34935_, _34934_);
  nor (_34938_, _06918_, _06130_);
  nor (_34939_, _34938_, _06924_);
  and (_34940_, _34938_, _06924_);
  nor (_34941_, _34940_, _34939_);
  or (_34942_, _34941_, _34936_);
  nand (_34943_, _34941_, _34936_);
  and (_34944_, _34943_, _34942_);
  or (_34945_, _34944_, _10342_);
  and (_34946_, _04944_, _30104_);
  nand (_34947_, _34946_, _34812_);
  or (_34949_, _34946_, _34829_);
  and (_34950_, _34949_, _34947_);
  or (_34951_, _34950_, _08105_);
  and (_34952_, _34951_, _08108_);
  and (_34953_, _34952_, _34945_);
  and (_34954_, _34931_, _08107_);
  or (_34955_, _34954_, _34953_);
  and (_34956_, _06140_, _03450_);
  and (_34957_, _34956_, _34955_);
  and (_34958_, _34829_, _10320_);
  or (_34960_, _34958_, _04624_);
  or (_34961_, _34960_, _34957_);
  nor (_34962_, _34819_, \oc8051_golden_model_1.ACC [6]);
  and (_34963_, _34819_, \oc8051_golden_model_1.ACC [6]);
  nor (_34964_, _34963_, _34962_);
  nor (_34965_, _34964_, \oc8051_golden_model_1.ACC [7]);
  and (_34966_, _34964_, \oc8051_golden_model_1.ACC [7]);
  nor (_34967_, _34966_, _34965_);
  not (_34968_, _34967_);
  nor (_34969_, _34968_, _34920_);
  and (_34971_, _34968_, _34920_);
  or (_34972_, _34971_, _34969_);
  or (_34973_, _34972_, _04625_);
  and (_34974_, _34973_, _04630_);
  and (_34975_, _34974_, _34961_);
  not (_34976_, _14985_);
  nor (_34977_, _15224_, _34976_);
  and (_34978_, _15224_, _34976_);
  nor (_34979_, _34978_, _34977_);
  and (_34980_, _34979_, _15472_);
  nor (_34982_, _34979_, _15472_);
  nor (_34983_, _34982_, _34980_);
  nor (_34984_, _34983_, _16477_);
  and (_34985_, _34983_, _16477_);
  or (_34986_, _34985_, _34984_);
  nor (_34987_, _16097_, _15828_);
  and (_34988_, _16097_, _15828_);
  nor (_34989_, _34988_, _34987_);
  not (_34990_, _34989_);
  not (_34991_, _16782_);
  nand (_34993_, _34991_, _08123_);
  or (_34994_, _34991_, _08123_);
  and (_34995_, _34994_, _34993_);
  nand (_34996_, _34995_, _34990_);
  or (_34997_, _34995_, _34990_);
  and (_34998_, _34997_, _34996_);
  nor (_34999_, _34998_, _34986_);
  and (_35000_, _34998_, _34986_);
  or (_35001_, _35000_, _34999_);
  and (_35002_, _35001_, _03757_);
  or (_35004_, _35002_, _08120_);
  or (_35005_, _35004_, _34975_);
  and (_35006_, _15228_, _07740_);
  or (_35007_, _35006_, _15478_);
  and (_35008_, _35007_, _16104_);
  nor (_35009_, _35007_, _16104_);
  nor (_35010_, _35009_, _35008_);
  nor (_35011_, _15835_, _15423_);
  and (_35012_, _15835_, _15423_);
  nor (_35013_, _35012_, _35011_);
  and (_35015_, _35013_, _35010_);
  nor (_35016_, _35013_, _35010_);
  nor (_35017_, _35016_, _35015_);
  and (_35018_, _35017_, _16484_);
  nor (_35019_, _35017_, _16484_);
  nor (_35020_, _35019_, _35018_);
  nor (_35021_, _16790_, _08146_);
  and (_35022_, _16790_, _08146_);
  nor (_35023_, _35022_, _35021_);
  nand (_35024_, _35023_, _35020_);
  or (_35026_, _35023_, _35020_);
  and (_35027_, _35026_, _35024_);
  or (_35028_, _35027_, _11746_);
  and (_35029_, _35028_, _35005_);
  or (_35030_, _35029_, _10353_);
  or (_35031_, _34829_, _11759_);
  and (_35032_, _35031_, _03697_);
  and (_35033_, _35032_, _35030_);
  not (_35034_, _15839_);
  and (_35035_, _35034_, _15486_);
  nor (_35037_, _35034_, _15486_);
  nor (_35038_, _35037_, _35035_);
  nor (_35039_, _15237_, _14991_);
  and (_35040_, _15237_, _14991_);
  nor (_35041_, _35040_, _35039_);
  not (_35042_, _35041_);
  and (_35043_, _35042_, _35038_);
  nor (_35044_, _35042_, _35038_);
  nor (_35045_, _35044_, _35043_);
  not (_35046_, _16796_);
  nor (_35048_, _16488_, _16111_);
  and (_35049_, _16488_, _16111_);
  nor (_35050_, _35049_, _35048_);
  nor (_35051_, _35050_, _35046_);
  and (_35052_, _35050_, _35046_);
  nor (_35053_, _35052_, _35051_);
  nor (_35054_, _35053_, _35045_);
  and (_35055_, _35053_, _35045_);
  nor (_35056_, _35055_, _35054_);
  and (_35057_, _35056_, _08152_);
  nor (_35059_, _35056_, _08152_);
  or (_35060_, _35059_, _35057_);
  and (_35061_, _35060_, _03696_);
  or (_35062_, _35061_, _04933_);
  or (_35063_, _35062_, _35033_);
  or (_35064_, _34829_, _03445_);
  and (_35065_, _35064_, _35063_);
  or (_35066_, _35065_, _03755_);
  and (_35067_, _15196_, _14963_);
  nor (_35068_, _15196_, _14963_);
  nor (_35070_, _35068_, _35067_);
  and (_35071_, _35070_, _15454_);
  nor (_35072_, _35070_, _15454_);
  or (_35073_, _35072_, _35071_);
  and (_35074_, _35073_, _15781_);
  nor (_35075_, _35073_, _15781_);
  or (_35076_, _35075_, _35074_);
  nor (_35077_, _16424_, _16082_);
  and (_35078_, _16424_, _16082_);
  nor (_35079_, _35078_, _35077_);
  and (_35081_, _35079_, _16752_);
  nor (_35082_, _35079_, _16752_);
  nor (_35083_, _35082_, _35081_);
  nor (_35084_, _35083_, _35076_);
  and (_35085_, _35083_, _35076_);
  nor (_35086_, _35085_, _35084_);
  nand (_35087_, _35086_, _08096_);
  or (_35088_, _35086_, _08096_);
  and (_35089_, _35088_, _35087_);
  or (_35090_, _35089_, _04537_);
  and (_35092_, _35090_, _14968_);
  and (_35093_, _35092_, _35066_);
  and (_35094_, _34944_, _04839_);
  or (_35095_, _35094_, _34914_);
  or (_35096_, _35095_, _35093_);
  and (_35097_, _35096_, _34932_);
  or (_35098_, _35097_, _04247_);
  not (_35099_, _04247_);
  or (_35100_, _34931_, _35099_);
  and (_35101_, _35100_, _03751_);
  and (_35103_, _35101_, _35098_);
  nor (_35104_, _12225_, _05699_);
  and (_35105_, _12595_, _06242_);
  nor (_35106_, _35105_, _35104_);
  nor (_35107_, _06241_, _05901_);
  nor (_35108_, _35107_, _05554_);
  and (_35109_, _35107_, _05554_);
  nor (_35110_, _35109_, _35108_);
  nor (_35111_, _35110_, _06018_);
  and (_35112_, _35110_, _06018_);
  nor (_35114_, _35112_, _35111_);
  not (_35115_, _35114_);
  nand (_35116_, _35115_, _35106_);
  or (_35117_, _35115_, _35106_);
  and (_35118_, _35117_, _03750_);
  and (_35119_, _35118_, _35116_);
  or (_35120_, _35119_, _10377_);
  or (_35121_, _35120_, _35103_);
  or (_35122_, _34829_, _10375_);
  and (_35123_, _35122_, _03692_);
  and (_35125_, _35123_, _35121_);
  nor (_35126_, _15255_, _14954_);
  and (_35127_, _15255_, _14954_);
  nor (_35128_, _35127_, _35126_);
  not (_35129_, _35128_);
  not (_35130_, _15858_);
  and (_35131_, _35130_, _15504_);
  nor (_35132_, _35130_, _15504_);
  nor (_35133_, _35132_, _35131_);
  and (_35134_, _35133_, _35129_);
  nor (_35136_, _35133_, _35129_);
  nor (_35137_, _35136_, _35134_);
  nor (_35138_, _16508_, _16130_);
  and (_35139_, _16508_, _16130_);
  nor (_35140_, _35139_, _35138_);
  not (_35141_, _16816_);
  and (_35142_, _35141_, _08169_);
  nor (_35143_, _35141_, _08169_);
  or (_35144_, _35143_, _35142_);
  or (_35145_, _35144_, _35140_);
  nand (_35147_, _35144_, _35140_);
  and (_35148_, _35147_, _35145_);
  nor (_35149_, _35148_, _35137_);
  and (_35150_, _35148_, _35137_);
  or (_35151_, _35150_, _35149_);
  nand (_35152_, _35151_, _03691_);
  not (_35153_, _03851_);
  and (_35154_, _10380_, _35153_);
  nand (_35155_, _35154_, _35152_);
  or (_35156_, _35155_, _35125_);
  or (_35158_, _35154_, _34829_);
  not (_35159_, _03863_);
  nor (_35160_, _03868_, _03859_);
  and (_35161_, _35160_, _03855_);
  and (_35162_, _35161_, _03871_);
  and (_35163_, _35162_, _35159_);
  and (_35164_, _35163_, _35158_);
  and (_35165_, _35164_, _35156_);
  not (_35166_, _35163_);
  nand (_35167_, _35166_, _34829_);
  nand (_35169_, _35167_, _10433_);
  or (_35170_, _35169_, _35165_);
  or (_35171_, _34829_, _10433_);
  and (_35172_, _35171_, _03685_);
  and (_35173_, _35172_, _35170_);
  not (_35174_, _16462_);
  nor (_35175_, _15509_, _15260_);
  and (_35176_, _15509_, _15260_);
  nor (_35177_, _35176_, _35175_);
  nor (_35178_, _35177_, _35174_);
  and (_35180_, _35177_, _35174_);
  nor (_35181_, _35180_, _35178_);
  not (_35182_, _35181_);
  nor (_35183_, _15810_, _34976_);
  and (_35184_, _15810_, _34976_);
  nor (_35185_, _35184_, _35183_);
  and (_35186_, _35185_, _16136_);
  nor (_35187_, _35185_, _16136_);
  nor (_35188_, _35187_, _35186_);
  nor (_35189_, _16821_, _08174_);
  and (_35191_, _16821_, _08174_);
  nor (_35192_, _35191_, _35189_);
  not (_35193_, _35192_);
  nor (_35194_, _35193_, _35188_);
  and (_35195_, _35193_, _35188_);
  nor (_35196_, _35195_, _35194_);
  nand (_35197_, _35196_, _35182_);
  or (_35198_, _35196_, _35182_);
  and (_35199_, _35198_, _03684_);
  nand (_35200_, _35199_, _35197_);
  and (_35202_, _03850_, _03783_);
  or (_35203_, _35202_, _05105_);
  nor (_35204_, _35203_, _03777_);
  nand (_35205_, _35204_, _35200_);
  or (_35206_, _35205_, _35173_);
  or (_35207_, _35204_, _34829_);
  and (_35208_, _03862_, _03783_);
  not (_35209_, _35208_);
  and (_35210_, _26072_, _35209_);
  and (_35211_, _35210_, _35207_);
  and (_35213_, _35211_, _35206_);
  not (_35214_, _35210_);
  and (_35215_, _35214_, _34829_);
  and (_35216_, _08102_, _03783_);
  or (_35217_, _35216_, _35215_);
  or (_35218_, _35217_, _35213_);
  not (_35219_, _35216_);
  or (_35220_, _35219_, _34829_);
  and (_35221_, _35220_, _07030_);
  and (_35222_, _35221_, _35218_);
  nor (_35224_, _09821_, _25787_);
  nand (_35225_, _35224_, _11667_);
  nor (_35226_, _15266_, _15015_);
  and (_35227_, _15266_, _15015_);
  or (_35228_, _35227_, _35226_);
  nor (_35229_, _35228_, _15514_);
  and (_35230_, _35228_, _15514_);
  nor (_35231_, _35230_, _35229_);
  nor (_35232_, _35231_, _15865_);
  and (_35233_, _35231_, _15865_);
  or (_35235_, _35233_, _35232_);
  nor (_35236_, _35235_, _16141_);
  and (_35237_, _35235_, _16141_);
  or (_35238_, _35237_, _35236_);
  nor (_35239_, _35238_, _16516_);
  and (_35240_, _35238_, _16516_);
  or (_35241_, _35240_, _35239_);
  nor (_35242_, _35241_, _16827_);
  and (_35243_, _35241_, _16827_);
  or (_35244_, _35243_, _35242_);
  or (_35246_, _35244_, _08179_);
  nand (_35247_, _35244_, _08179_);
  and (_35248_, _35247_, _07024_);
  and (_35249_, _35248_, _35246_);
  or (_35250_, _35249_, _35225_);
  or (_35251_, _35250_, _35222_);
  not (_35252_, _35225_);
  or (_35253_, _35252_, _34829_);
  and (_35254_, _35253_, _11666_);
  and (_35255_, _35254_, _35251_);
  and (_35257_, _34829_, _03810_);
  or (_35258_, _35257_, _08182_);
  or (_35259_, _35258_, _35255_);
  or (_35260_, _15274_, _15020_);
  nand (_35261_, _15274_, _15020_);
  and (_35262_, _35261_, _35260_);
  nor (_35263_, _35262_, _15532_);
  and (_35264_, _35262_, _15532_);
  nor (_35265_, _35264_, _35263_);
  nand (_35266_, _35265_, _15805_);
  or (_35268_, _35265_, _15805_);
  and (_35269_, _35268_, _35266_);
  or (_35270_, _35269_, _16160_);
  nand (_35271_, _35269_, _16160_);
  and (_35272_, _35271_, _35270_);
  nor (_35273_, _35272_, _16455_);
  and (_35274_, _35272_, _16455_);
  or (_35275_, _35274_, _35273_);
  nor (_35276_, _35275_, _16843_);
  and (_35277_, _35275_, _16843_);
  nor (_35279_, _35277_, _35276_);
  or (_35280_, _08258_, _08181_);
  or (_35281_, _35280_, _35279_);
  not (_35282_, _35279_);
  or (_35283_, _35282_, _08259_);
  and (_35284_, _35283_, _08261_);
  and (_35285_, _35284_, _35281_);
  and (_35286_, _35285_, _35259_);
  not (_35287_, _08283_);
  or (_35288_, _15205_, _14966_);
  nand (_35290_, _15205_, _14966_);
  and (_35291_, _35290_, _35288_);
  nor (_35292_, _35291_, _15550_);
  and (_35293_, _35291_, _15550_);
  or (_35294_, _35293_, _35292_);
  nor (_35295_, _35294_, _15882_);
  and (_35296_, _35294_, _15882_);
  nor (_35297_, _35296_, _35295_);
  nor (_35298_, _35297_, _16179_);
  and (_35299_, _35297_, _16179_);
  nor (_35301_, _35299_, _35298_);
  nor (_35302_, _35301_, _16535_);
  and (_35303_, _35301_, _16535_);
  or (_35304_, _35303_, _35302_);
  nor (_35305_, _35304_, _16766_);
  and (_35306_, _35304_, _16766_);
  nor (_35307_, _35306_, _35305_);
  nand (_35308_, _35307_, _35287_);
  or (_35309_, _35307_, _35287_);
  and (_35310_, _35309_, _08260_);
  and (_35312_, _35310_, _35308_);
  or (_35313_, _35312_, _03818_);
  or (_35314_, _35313_, _35286_);
  not (_35315_, _08358_);
  nor (_35316_, _15284_, _15027_);
  and (_35317_, _15284_, _15027_);
  or (_35318_, _35317_, _35316_);
  and (_35319_, _35318_, _15565_);
  nor (_35320_, _35318_, _15565_);
  or (_35321_, _35320_, _35319_);
  nor (_35323_, _35321_, _15898_);
  and (_35324_, _35321_, _15898_);
  nor (_35325_, _35324_, _35323_);
  or (_35326_, _35325_, _16195_);
  nand (_35327_, _35325_, _16195_);
  and (_35328_, _35327_, _35326_);
  nor (_35329_, _35328_, _16553_);
  and (_35330_, _35328_, _16553_);
  or (_35331_, _35330_, _35329_);
  and (_35332_, _35331_, _16860_);
  nor (_35334_, _35331_, _16860_);
  nor (_35335_, _35334_, _35332_);
  nand (_35336_, _35335_, _35315_);
  or (_35337_, _35335_, _35315_);
  and (_35338_, _35337_, _08288_);
  and (_35339_, _35338_, _35336_);
  or (_35340_, _35339_, _10492_);
  and (_35341_, _35340_, _35314_);
  nor (_35342_, _15292_, _15032_);
  and (_35343_, _15292_, _15032_);
  or (_35345_, _35343_, _35342_);
  and (_35346_, _35345_, _15582_);
  nor (_35347_, _35345_, _15582_);
  or (_35348_, _35347_, _35346_);
  nor (_35349_, _35348_, _15793_);
  and (_35350_, _35348_, _15793_);
  nor (_35351_, _35350_, _35349_);
  or (_35352_, _35351_, _16212_);
  nand (_35353_, _35351_, _16212_);
  and (_35354_, _35353_, _35352_);
  or (_35356_, _35354_, _16440_);
  nand (_35357_, _35354_, _16440_);
  and (_35358_, _35357_, _35356_);
  nor (_35359_, _35358_, _16874_);
  and (_35360_, _35358_, _16874_);
  nor (_35361_, _35360_, _35359_);
  and (_35362_, _35361_, _08425_);
  nor (_35363_, _35361_, _08425_);
  or (_35364_, _35363_, _35362_);
  and (_35365_, _35364_, _08287_);
  or (_35367_, _35365_, _03547_);
  or (_35368_, _35367_, _35341_);
  nor (_35369_, _05344_, _03741_);
  nor (_35370_, _05363_, _05358_);
  nor (_35371_, _05402_, _05349_);
  or (_35372_, _05388_, _05341_);
  and (_35373_, _35372_, _35371_);
  nor (_35374_, _35372_, _35371_);
  nor (_35375_, _35374_, _35373_);
  nor (_35376_, _35375_, _35370_);
  and (_35378_, _35375_, _35370_);
  nor (_35379_, _35378_, _35376_);
  nor (_35380_, _35379_, _35369_);
  and (_35381_, _35379_, _35369_);
  or (_35382_, _35381_, _35380_);
  or (_35383_, _35382_, _03422_);
  and (_35384_, _35383_, _03680_);
  and (_35385_, _35384_, _35368_);
  and (_35386_, _15300_, _15040_);
  nor (_35387_, _15300_, _15040_);
  or (_35389_, _35387_, _35386_);
  and (_35390_, _35389_, _15590_);
  nor (_35391_, _35389_, _15590_);
  or (_35392_, _35391_, _35390_);
  and (_35393_, _35392_, _15908_);
  nor (_35394_, _35392_, _15908_);
  or (_35395_, _35394_, _35393_);
  not (_35396_, _16883_);
  nor (_35397_, _16564_, _16221_);
  and (_35398_, _16564_, _16221_);
  nor (_35401_, _35398_, _35397_);
  nor (_35402_, _35401_, _35396_);
  and (_35403_, _35401_, _35396_);
  nor (_35404_, _35403_, _35402_);
  nor (_35405_, _35404_, _35395_);
  and (_35406_, _35404_, _35395_);
  or (_35407_, _35406_, _35405_);
  or (_35408_, _35407_, _08434_);
  nand (_35409_, _35407_, _08434_);
  and (_35410_, _35409_, _03679_);
  and (_35412_, _35410_, _35408_);
  or (_35413_, _35412_, _28935_);
  or (_35414_, _35413_, _35385_);
  and (_35415_, _35414_, _34913_);
  or (_35416_, _35415_, _07544_);
  or (_35417_, _35089_, _06994_);
  and (_35418_, _35417_, _04679_);
  and (_35419_, _35418_, _35416_);
  not (_35420_, _16891_);
  and (_35421_, _35420_, _08441_);
  nor (_35424_, _35420_, _08441_);
  nor (_35425_, _35424_, _35421_);
  not (_35426_, _16572_);
  and (_35427_, _35426_, _16228_);
  nor (_35428_, _35426_, _16228_);
  nor (_35429_, _35428_, _35427_);
  and (_35430_, _15307_, _15047_);
  nor (_35431_, _15307_, _15047_);
  nor (_35432_, _35431_, _35430_);
  not (_35433_, _35432_);
  not (_35435_, _15915_);
  and (_35436_, _35435_, _15597_);
  nor (_35437_, _35435_, _15597_);
  nor (_35438_, _35437_, _35436_);
  and (_35439_, _35438_, _35433_);
  nor (_35440_, _35438_, _35433_);
  nor (_35441_, _35440_, _35439_);
  nor (_35442_, _35441_, _35429_);
  and (_35443_, _35441_, _35429_);
  nor (_35444_, _35443_, _35442_);
  or (_35447_, _35444_, _35425_);
  nand (_35448_, _35444_, _35425_);
  and (_35449_, _35448_, _35447_);
  and (_35450_, _35449_, _04678_);
  or (_35451_, _35450_, _07559_);
  or (_35452_, _35451_, _35419_);
  not (_35453_, _16234_);
  and (_35454_, _15312_, _14960_);
  nor (_35455_, _15312_, _14960_);
  nor (_35456_, _35455_, _35454_);
  and (_35458_, _35456_, _15602_);
  nor (_35459_, _35456_, _15602_);
  or (_35460_, _35459_, _35458_);
  nand (_35461_, _35460_, _15920_);
  or (_35462_, _35460_, _15920_);
  and (_35463_, _35462_, _35461_);
  nor (_35464_, _35463_, _35453_);
  and (_35465_, _35463_, _35453_);
  or (_35466_, _35465_, _35464_);
  and (_35467_, _35466_, _16577_);
  nor (_35470_, _35466_, _16577_);
  or (_35471_, _35470_, _35467_);
  and (_35472_, _35471_, _16896_);
  nor (_35473_, _35471_, _16896_);
  or (_35474_, _35473_, _35472_);
  and (_35475_, _35474_, _08446_);
  nor (_35476_, _35474_, _08446_);
  or (_35477_, _35476_, _35475_);
  or (_35478_, _35477_, _03415_);
  and (_35479_, _35478_, _07565_);
  and (_35481_, _35479_, _35452_);
  and (_35482_, _07619_, _16902_);
  nor (_35483_, _07619_, _16902_);
  nor (_35484_, _35483_, _35482_);
  nor (_35485_, _07703_, _07652_);
  and (_35486_, _07703_, _07652_);
  nor (_35487_, _35486_, _35485_);
  not (_35488_, _35487_);
  and (_35489_, _35488_, _07760_);
  nor (_35490_, _35488_, _07760_);
  nor (_35492_, _35490_, _35489_);
  not (_35493_, _35492_);
  nor (_35494_, _35493_, _35484_);
  and (_35495_, _35493_, _35484_);
  or (_35496_, _35495_, _35494_);
  or (_35497_, _35496_, _07577_);
  nand (_35498_, _35496_, _07577_);
  and (_35499_, _35498_, _35497_);
  nor (_35500_, _35499_, _07835_);
  and (_35501_, _35499_, _07835_);
  nor (_35503_, _35501_, _35500_);
  nand (_35504_, _35503_, _14421_);
  or (_35505_, _35503_, _14421_);
  and (_35506_, _35505_, _07558_);
  and (_35507_, _35506_, _35504_);
  or (_35508_, _35507_, _03466_);
  or (_35509_, _35508_, _35481_);
  or (_35510_, _35382_, _03467_);
  and (_35511_, _35510_, _27577_);
  and (_35512_, _35511_, _35509_);
  nand (_35514_, _34829_, _03746_);
  not (_35515_, _03482_);
  not (_35516_, _03797_);
  nor (_35517_, _04110_, _03786_);
  and (_35518_, _35517_, _35516_);
  nor (_35519_, _35518_, _35515_);
  not (_35520_, _35519_);
  nor (_35521_, _04689_, _04685_);
  and (_35522_, _35521_, _06302_);
  and (_35523_, _35522_, _25812_);
  and (_35525_, _35523_, _35520_);
  nand (_35526_, _35525_, _35514_);
  or (_35527_, _35526_, _35512_);
  or (_35528_, _35525_, _34829_);
  and (_35529_, _35528_, _04694_);
  and (_35530_, _35529_, _35527_);
  nor (_35531_, _15930_, _15612_);
  and (_35532_, _15930_, _15612_);
  nor (_35533_, _35532_, _35531_);
  nor (_35534_, _15322_, _15058_);
  and (_35536_, _15322_, _15058_);
  or (_35537_, _35536_, _35534_);
  nor (_35538_, _35537_, _35533_);
  and (_35539_, _35537_, _35533_);
  nor (_35540_, _35539_, _35538_);
  not (_35541_, _16909_);
  nor (_35542_, _16588_, _16245_);
  and (_35543_, _16588_, _16245_);
  nor (_35544_, _35543_, _35542_);
  nor (_35545_, _35544_, _35541_);
  and (_35547_, _35544_, _35541_);
  nor (_35548_, _35547_, _35545_);
  nor (_35549_, _35548_, _35540_);
  and (_35550_, _35548_, _35540_);
  or (_35551_, _35550_, _35549_);
  or (_35552_, _35551_, _08459_);
  nand (_35553_, _35551_, _08459_);
  and (_35554_, _35553_, _03839_);
  and (_35555_, _35554_, _35552_);
  or (_35556_, _35555_, _35530_);
  and (_35558_, _35556_, _08457_);
  nand (_35559_, _35382_, _08456_);
  nor (_35560_, _10540_, _10145_);
  and (_35561_, _35560_, _10543_);
  nand (_35562_, _35561_, _35559_);
  or (_35563_, _35562_, _35558_);
  and (_35564_, _03850_, _03485_);
  nor (_35565_, _35561_, _34829_);
  nor (_35566_, _35565_, _35564_);
  and (_35567_, _35566_, _35563_);
  and (_35569_, _16923_, _08468_);
  nor (_35570_, _16923_, _08468_);
  nor (_35571_, _35570_, _35569_);
  and (_35572_, _15065_, _08666_);
  nor (_35573_, _35572_, _15525_);
  nor (_35574_, _15761_, _08662_);
  and (_35575_, _15761_, _08662_);
  nor (_35576_, _35575_, _35574_);
  nor (_35577_, _35576_, _35573_);
  and (_35578_, _35576_, _35573_);
  nor (_35580_, _35578_, _35577_);
  nor (_35581_, _08653_, _08657_);
  and (_35582_, _08653_, _08657_);
  nor (_35583_, _35582_, _35581_);
  nor (_35584_, _35583_, _35580_);
  and (_35585_, _35583_, _35580_);
  nor (_35586_, _35585_, _35584_);
  nor (_35587_, _35586_, _35571_);
  and (_35588_, _35586_, _35571_);
  or (_35589_, _35588_, _35587_);
  and (_35591_, _35589_, _35564_);
  nor (_35592_, _04970_, _03785_);
  nor (_35593_, _35592_, _15620_);
  or (_35594_, _35593_, _35591_);
  or (_35595_, _35594_, _35567_);
  not (_35596_, _35593_);
  or (_35597_, _35596_, _35589_);
  and (_35598_, _35597_, _16260_);
  and (_35599_, _35598_, _35595_);
  not (_35600_, _07972_);
  and (_35602_, _35600_, _07969_);
  nor (_35603_, _35600_, _07969_);
  nor (_35604_, _35603_, _35602_);
  and (_35605_, _14941_, _07988_);
  nor (_35606_, _35605_, _15543_);
  and (_35607_, _15871_, _07984_);
  nor (_35608_, _15871_, _07984_);
  nor (_35609_, _35608_, _35607_);
  nor (_35610_, _35609_, _35606_);
  and (_35611_, _35609_, _35606_);
  nor (_35613_, _35611_, _35610_);
  and (_35614_, _07979_, _07975_);
  nor (_35615_, _07979_, _07975_);
  nor (_35616_, _35615_, _35614_);
  nor (_35617_, _35616_, _35613_);
  and (_35618_, _35616_, _35613_);
  nor (_35619_, _35618_, _35617_);
  nor (_35620_, _35619_, _35604_);
  and (_35621_, _35619_, _35604_);
  or (_35622_, _35621_, _35620_);
  and (_35624_, _35622_, _16259_);
  or (_35625_, _35624_, _04339_);
  or (_35626_, _35625_, _35599_);
  or (_35627_, _35622_, _16078_);
  and (_35628_, _35627_, _03958_);
  and (_35629_, _35628_, _35626_);
  and (_35630_, _10455_, _08707_);
  nor (_35631_, _35630_, _10456_);
  and (_35632_, _35631_, _08700_);
  nor (_35633_, _35631_, _08700_);
  nor (_35635_, _35633_, _35632_);
  not (_35636_, _10459_);
  and (_35637_, _35636_, _08711_);
  nor (_35638_, _35637_, _10460_);
  nor (_35639_, _10451_, _06523_);
  and (_35640_, _10451_, _06523_);
  nor (_35641_, _35640_, _35639_);
  nor (_35642_, _35641_, _35638_);
  and (_35643_, _35641_, _35638_);
  nor (_35644_, _35643_, _35642_);
  and (_35646_, _35644_, _08695_);
  nor (_35647_, _35644_, _08695_);
  nor (_35648_, _35647_, _35646_);
  not (_35649_, _35648_);
  nor (_35650_, _35649_, _35635_);
  and (_35651_, _35649_, _35635_);
  or (_35652_, _35651_, _08478_);
  or (_35653_, _35652_, _35650_);
  and (_35654_, _35653_, _10590_);
  or (_35655_, _35654_, _35629_);
  and (_35657_, _08736_, _08740_);
  nor (_35658_, _35657_, _10436_);
  not (_35659_, _35658_);
  and (_35660_, _10439_, _08745_);
  nor (_35661_, _35660_, _10440_);
  nor (_35662_, _08751_, _10443_);
  nor (_35663_, _35662_, _10444_);
  and (_35664_, _35663_, _35661_);
  nor (_35665_, _35663_, _35661_);
  nor (_35666_, _35665_, _35664_);
  nor (_35668_, _35666_, _35659_);
  and (_35669_, _35666_, _35659_);
  nor (_35670_, _35669_, _35668_);
  and (_35671_, _08733_, _08485_);
  nor (_35672_, _35671_, _10437_);
  nor (_35673_, _35672_, _35670_);
  and (_35674_, _35672_, _35670_);
  or (_35675_, _35674_, _35673_);
  or (_35676_, _35675_, _08479_);
  and (_35677_, _35676_, _04703_);
  and (_35679_, _35677_, _35655_);
  or (_35680_, _35679_, _34912_);
  and (_35681_, _35680_, _10597_);
  nand (_35682_, _34829_, _03959_);
  nor (_35683_, _35682_, _05365_);
  or (_35684_, _35683_, _35681_);
  and (_35685_, _35684_, _10602_);
  nor (_35686_, _35685_, _34887_);
  nor (_35687_, _35686_, _34886_);
  and (_35688_, _25955_, _03420_);
  or (_35690_, _08667_, _08664_);
  nand (_35691_, _08667_, _08664_);
  and (_35692_, _35691_, _35690_);
  and (_35693_, _15959_, _08660_);
  nor (_35694_, _15959_, _08660_);
  nor (_35695_, _35694_, _35693_);
  not (_35696_, _35695_);
  and (_35697_, _35696_, _35692_);
  nor (_35698_, _35696_, _35692_);
  nor (_35699_, _35698_, _35697_);
  not (_35701_, _08651_);
  nor (_35702_, _08655_, _08648_);
  and (_35703_, _08655_, _08648_);
  nor (_35704_, _35703_, _35702_);
  nor (_35705_, _35704_, _35701_);
  and (_35706_, _35704_, _35701_);
  nor (_35707_, _35706_, _35705_);
  not (_35708_, _35707_);
  nor (_35709_, _35708_, _35699_);
  and (_35710_, _35708_, _35699_);
  nor (_35712_, _35710_, _35709_);
  nand (_35713_, _35712_, _08467_);
  or (_35714_, _35712_, _08467_);
  and (_35715_, _35714_, _35713_);
  and (_35716_, _35715_, _34886_);
  or (_35717_, _35716_, _35688_);
  or (_35718_, _35717_, _35687_);
  not (_35719_, _35688_);
  nor (_35720_, _35715_, _35719_);
  and (_35721_, _14951_, _03382_);
  nor (_35723_, _35721_, _35720_);
  and (_35724_, _35723_, _35718_);
  and (_35725_, _35721_, _35715_);
  or (_35726_, _35725_, _16739_);
  or (_35727_, _35726_, _35724_);
  not (_35728_, _16739_);
  or (_35729_, _35715_, _35728_);
  and (_35730_, _35729_, _08086_);
  and (_35731_, _35730_, _35727_);
  and (_35732_, _35715_, _08085_);
  or (_35734_, _35732_, _08502_);
  or (_35735_, _35734_, _35731_);
  not (_35736_, _07982_);
  or (_35737_, _07989_, _07986_);
  nand (_35738_, _07989_, _07986_);
  and (_35739_, _35738_, _35737_);
  nand (_35740_, _35739_, _35736_);
  or (_35741_, _35739_, _35736_);
  and (_35742_, _35741_, _35740_);
  nor (_35743_, _35742_, _07980_);
  and (_35745_, _35742_, _07980_);
  or (_35746_, _35745_, _35743_);
  nor (_35747_, _07977_, _07973_);
  and (_35748_, _07977_, _07973_);
  nor (_35749_, _35748_, _35747_);
  nor (_35750_, _35749_, _07970_);
  and (_35751_, _35749_, _07970_);
  nor (_35752_, _35751_, _35750_);
  not (_35753_, _35752_);
  and (_35754_, _35753_, _35746_);
  nor (_35756_, _35753_, _35746_);
  nor (_35757_, _35756_, _35754_);
  and (_35758_, _35757_, _07968_);
  nor (_35759_, _35757_, _07968_);
  or (_35760_, _35759_, _08503_);
  or (_35761_, _35760_, _35758_);
  and (_35762_, _35761_, _03966_);
  and (_35763_, _35762_, _35735_);
  not (_35764_, _08698_);
  or (_35765_, _08712_, _08709_);
  nand (_35767_, _08712_, _08709_);
  and (_35768_, _35767_, _35765_);
  and (_35769_, _08704_, _08705_);
  nor (_35770_, _08704_, _08705_);
  nor (_35771_, _35770_, _35769_);
  not (_35772_, _35771_);
  and (_35773_, _35772_, _35768_);
  nor (_35774_, _35772_, _35768_);
  nor (_35775_, _35774_, _35773_);
  nand (_35776_, _35775_, _35764_);
  or (_35778_, _35775_, _35764_);
  and (_35779_, _35778_, _35776_);
  or (_35780_, _35779_, _08696_);
  nand (_35781_, _35779_, _08696_);
  and (_35782_, _35781_, _35780_);
  nor (_35783_, _35782_, _08693_);
  and (_35784_, _35782_, _08693_);
  or (_35785_, _35784_, _35783_);
  and (_35786_, _35785_, _11960_);
  nor (_35787_, _35785_, _11960_);
  or (_35789_, _35787_, _35786_);
  and (_35790_, _35789_, _03965_);
  or (_35791_, _35790_, _08508_);
  or (_35792_, _35791_, _35763_);
  not (_35793_, _08738_);
  or (_35794_, _08747_, _08748_);
  nand (_35795_, _08747_, _08748_);
  and (_35796_, _35795_, _35794_);
  not (_35797_, _08741_);
  and (_35798_, _35797_, _08743_);
  nor (_35800_, _35797_, _08743_);
  nor (_35801_, _35800_, _35798_);
  not (_35802_, _35801_);
  and (_35803_, _35802_, _35796_);
  nor (_35804_, _35802_, _35796_);
  nor (_35805_, _35804_, _35803_);
  nand (_35806_, _35805_, _35793_);
  or (_35807_, _35805_, _35793_);
  and (_35808_, _35807_, _35806_);
  or (_35809_, _35808_, _08734_);
  nand (_35811_, _35808_, _08734_);
  and (_35812_, _35811_, _35809_);
  or (_35813_, _35812_, _08731_);
  nand (_35814_, _35812_, _08731_);
  and (_35815_, _35814_, _35813_);
  nand (_35816_, _35815_, _11966_);
  or (_35817_, _35815_, _11966_);
  and (_35818_, _35817_, _35816_);
  or (_35819_, _35818_, _08509_);
  and (_35820_, _35819_, _04708_);
  and (_35822_, _35820_, _35792_);
  and (_35823_, _10031_, _10030_);
  nor (_35824_, _15659_, _15097_);
  and (_35825_, _15659_, _15097_);
  nor (_35826_, _35825_, _35824_);
  nor (_35827_, _16963_, _16301_);
  and (_35828_, _16963_, _16301_);
  nor (_35829_, _35828_, _35827_);
  and (_35830_, _35829_, _35826_);
  nor (_35831_, _35829_, _35826_);
  nor (_35833_, _35831_, _35830_);
  not (_35834_, _35833_);
  nor (_35835_, _15975_, _15359_);
  and (_35836_, _15975_, _15359_);
  nor (_35837_, _35836_, _35835_);
  nor (_35838_, _16634_, _08516_);
  and (_35839_, _16634_, _08516_);
  nor (_35840_, _35839_, _35838_);
  and (_35841_, _35840_, _35837_);
  nor (_35842_, _35840_, _35837_);
  nor (_35844_, _35842_, _35841_);
  nand (_35845_, _35844_, _35834_);
  or (_35846_, _35844_, _35834_);
  and (_35847_, _35846_, _03866_);
  nand (_35848_, _35847_, _35845_);
  nand (_35849_, _35848_, _35823_);
  or (_35850_, _35849_, _35822_);
  or (_35851_, _34829_, _35823_);
  and (_35852_, _35851_, _10020_);
  and (_35853_, _35852_, _35850_);
  or (_35855_, _35853_, _34885_);
  and (_35856_, _35855_, _10025_);
  nor (_35857_, _34884_, _08521_);
  nor (_35858_, _35857_, _10026_);
  or (_35859_, _35858_, _35856_);
  nor (_35860_, _14940_, _07987_);
  and (_35861_, _14940_, _07987_);
  nor (_35862_, _35861_, _35860_);
  and (_35863_, _35862_, _07983_);
  nor (_35864_, _35862_, _07983_);
  or (_35866_, _35864_, _35863_);
  nand (_35867_, _35866_, _07981_);
  or (_35868_, _35866_, _07981_);
  and (_35869_, _35868_, _35867_);
  nor (_35870_, _07978_, _07971_);
  and (_35871_, _07978_, _07971_);
  nor (_35872_, _35871_, _35870_);
  and (_35873_, _35872_, _07974_);
  nor (_35874_, _35872_, _07974_);
  nor (_35875_, _35874_, _35873_);
  and (_35877_, _35875_, _35869_);
  nor (_35878_, _35875_, _35869_);
  or (_35879_, _35878_, _35877_);
  and (_35880_, _35879_, _11952_);
  nor (_35881_, _35879_, _11952_);
  or (_35882_, _35881_, _10021_);
  or (_35883_, _35882_, _35880_);
  and (_35884_, _35883_, _03953_);
  and (_35885_, _35884_, _35859_);
  nor (_35886_, _10458_, _08710_);
  and (_35888_, _10458_, _08710_);
  nor (_35889_, _35888_, _35886_);
  not (_35890_, _35889_);
  and (_35891_, _08702_, _08706_);
  nor (_35892_, _08702_, _08706_);
  nor (_35893_, _35892_, _35891_);
  nor (_35894_, _35893_, _35890_);
  and (_35895_, _35893_, _35890_);
  nor (_35896_, _35895_, _35894_);
  and (_35897_, _35896_, _08699_);
  nor (_35899_, _35896_, _08699_);
  or (_35900_, _35899_, _35897_);
  and (_35901_, _35900_, _08697_);
  nor (_35902_, _35900_, _08697_);
  or (_35903_, _35902_, _35901_);
  nand (_35904_, _35903_, _08694_);
  or (_35905_, _35903_, _08694_);
  and (_35906_, _35905_, _35904_);
  and (_35907_, _35906_, _11959_);
  nor (_35908_, _35906_, _11959_);
  or (_35910_, _35908_, _35907_);
  and (_35911_, _35910_, _03952_);
  or (_35912_, _35911_, _08526_);
  or (_35913_, _35912_, _35885_);
  nor (_35914_, _08750_, _10441_);
  and (_35915_, _08750_, _10441_);
  nor (_35916_, _35915_, _35914_);
  not (_35917_, _08742_);
  and (_35918_, _35917_, _08744_);
  nor (_35919_, _35917_, _08744_);
  nor (_35921_, _35919_, _35918_);
  and (_35922_, _35921_, _35916_);
  nor (_35923_, _35921_, _35916_);
  nor (_35924_, _35923_, _35922_);
  not (_35925_, _08739_);
  nor (_35926_, _08735_, _08732_);
  and (_35927_, _08735_, _08732_);
  nor (_35928_, _35927_, _35926_);
  nor (_35929_, _35928_, _35925_);
  and (_35930_, _35928_, _35925_);
  nor (_35932_, _35930_, _35929_);
  and (_35933_, _35932_, _35924_);
  nor (_35934_, _35932_, _35924_);
  or (_35935_, _35934_, _35933_);
  and (_35936_, _35935_, _08483_);
  nor (_35937_, _35935_, _08483_);
  or (_35938_, _35937_, _35936_);
  or (_35939_, _35938_, _08529_);
  and (_35940_, _35939_, _06532_);
  and (_35941_, _35940_, _35913_);
  and (_35943_, _10016_, _10015_);
  nor (_35944_, _15375_, _15121_);
  and (_35945_, _15375_, _15121_);
  or (_35946_, _35945_, _35944_);
  nor (_35947_, _15991_, _15681_);
  and (_35948_, _15991_, _15681_);
  nor (_35949_, _35948_, _35947_);
  nor (_35950_, _35949_, _35946_);
  and (_35951_, _35949_, _35946_);
  nor (_35952_, _35951_, _35950_);
  nor (_35954_, _16981_, _16654_);
  and (_35955_, _16981_, _16654_);
  nor (_35956_, _35955_, _35954_);
  not (_35957_, _16323_);
  and (_35958_, _35957_, _08537_);
  nor (_35959_, _35957_, _08537_);
  nor (_35960_, _35959_, _35958_);
  nor (_35961_, _35960_, _35956_);
  and (_35962_, _35960_, _35956_);
  nor (_35963_, _35962_, _35961_);
  not (_35965_, _35963_);
  nand (_35966_, _35965_, _35952_);
  or (_35967_, _35965_, _35952_);
  and (_35968_, _35967_, _03835_);
  nand (_35969_, _35968_, _35966_);
  nand (_35970_, _35969_, _35943_);
  or (_35971_, _35970_, _35941_);
  or (_35972_, _34829_, _35943_);
  and (_35973_, _35972_, _08547_);
  and (_35974_, _35973_, _35971_);
  or (_35976_, _35974_, _34859_);
  and (_35977_, _35976_, _34833_);
  and (_35978_, _08079_, _04083_);
  not (_35979_, _15998_);
  nor (_35980_, _15386_, _14966_);
  and (_35981_, _15386_, _14966_);
  or (_35982_, _35981_, _35980_);
  nor (_35983_, _35982_, _15691_);
  and (_35984_, _35982_, _15691_);
  nor (_35985_, _35984_, _35983_);
  and (_35987_, _35985_, _35979_);
  nor (_35988_, _35985_, _35979_);
  nor (_35989_, _35988_, _35987_);
  and (_35990_, _35989_, _16070_);
  nor (_35991_, _35989_, _16070_);
  nor (_35992_, _35991_, _35990_);
  nor (_35993_, _35992_, _16662_);
  and (_35994_, _35992_, _16662_);
  or (_35995_, _35994_, _35993_);
  nor (_35996_, _35995_, _16992_);
  and (_35998_, _35995_, _16992_);
  or (_35999_, _35998_, _35996_);
  and (_36000_, _35999_, _08078_);
  nor (_36001_, _35999_, _08078_);
  or (_36002_, _36001_, _36000_);
  and (_36003_, _36002_, _35978_);
  or (_36004_, _36003_, _04371_);
  or (_36005_, _36004_, _35977_);
  or (_36006_, _36002_, _04372_);
  and (_36007_, _36006_, _03964_);
  and (_36009_, _36007_, _36005_);
  not (_36010_, _16003_);
  nor (_36011_, _15391_, _15027_);
  and (_36012_, _15391_, _15027_);
  or (_36013_, _36012_, _36011_);
  nor (_36014_, _36013_, _15696_);
  and (_36015_, _36013_, _15696_);
  nor (_36016_, _36015_, _36014_);
  and (_36017_, _36016_, _36010_);
  nor (_36018_, _36016_, _36010_);
  nor (_36020_, _36018_, _36017_);
  nor (_36021_, _36020_, _16336_);
  and (_36022_, _36020_, _16336_);
  or (_36023_, _36022_, _36021_);
  and (_36024_, _36023_, _16667_);
  nor (_36025_, _36023_, _16667_);
  nor (_36026_, _36025_, _36024_);
  and (_36027_, _36026_, _16997_);
  nor (_36028_, _36026_, _16997_);
  or (_36029_, _36028_, _36027_);
  nor (_36031_, _36029_, _08605_);
  and (_36032_, _36029_, _08605_);
  or (_36033_, _36032_, _36031_);
  and (_36034_, _36033_, _03963_);
  or (_36035_, _36034_, _08580_);
  or (_36036_, _36035_, _36009_);
  and (_36037_, _15186_, _15032_);
  nor (_36038_, _15186_, _15032_);
  nor (_36039_, _36038_, _36037_);
  nor (_36040_, _36039_, _15701_);
  and (_36042_, _36039_, _15701_);
  nor (_36043_, _36042_, _36040_);
  and (_36044_, _36043_, _16008_);
  nor (_36045_, _36043_, _16008_);
  nor (_36046_, _36045_, _36044_);
  nor (_36047_, _36046_, _16342_);
  and (_36048_, _36046_, _16342_);
  or (_36049_, _36048_, _36047_);
  nor (_36050_, _36049_, _16673_);
  and (_36051_, _36049_, _16673_);
  or (_36053_, _36051_, _36050_);
  and (_36054_, _36053_, _17003_);
  nor (_36055_, _36053_, _17003_);
  nor (_36056_, _36055_, _36054_);
  nor (_36057_, _36056_, _08632_);
  and (_36058_, _36056_, _08632_);
  or (_36059_, _36058_, _08581_);
  or (_36060_, _36059_, _36057_);
  and (_36061_, _36060_, _08007_);
  and (_36062_, _36061_, _36036_);
  nor (_36064_, _15199_, _15198_);
  nor (_36065_, _15477_, \oc8051_golden_model_1.ACC [3]);
  and (_36066_, _15477_, \oc8051_golden_model_1.ACC [3]);
  nor (_36067_, _36066_, _36065_);
  and (_36068_, _36067_, _34964_);
  nor (_36069_, _36067_, _34964_);
  nor (_36070_, _36069_, _36068_);
  nor (_36071_, _36070_, _36064_);
  and (_36072_, _36070_, _36064_);
  or (_36073_, _36072_, _36071_);
  nand (_36075_, _36073_, _08006_);
  and (_36076_, _29052_, _11621_);
  nand (_36077_, _36076_, _36075_);
  or (_36078_, _36077_, _36062_);
  nor (_36079_, _36076_, _34829_);
  nor (_36080_, _36079_, _08639_);
  and (_36081_, _36080_, _36078_);
  nor (_36082_, _15401_, _15065_);
  nor (_36083_, _36082_, _35572_);
  nor (_36084_, _36083_, _15709_);
  and (_36086_, _36083_, _15709_);
  or (_36087_, _36086_, _36084_);
  nor (_36088_, _36087_, _15764_);
  and (_36089_, _36087_, _15764_);
  nor (_36090_, _36089_, _36088_);
  and (_36091_, _36090_, _16349_);
  nor (_36092_, _36090_, _16349_);
  nor (_36093_, _36092_, _36091_);
  nor (_36094_, _36093_, _16408_);
  and (_36095_, _36093_, _16408_);
  or (_36097_, _36095_, _36094_);
  nor (_36098_, _36097_, _17012_);
  and (_36099_, _36097_, _17012_);
  or (_36100_, _36099_, _36098_);
  or (_36101_, _36100_, _08682_);
  nand (_36102_, _36100_, _08682_);
  and (_36103_, _36102_, _36101_);
  nand (_36104_, _36103_, _08639_);
  nor (_36105_, _08642_, _08637_);
  nand (_36106_, _36105_, _36104_);
  or (_36108_, _36106_, _36081_);
  or (_36109_, _36105_, _36103_);
  and (_36110_, _36109_, _08647_);
  and (_36111_, _36110_, _36108_);
  and (_36112_, _36103_, _04392_);
  or (_36113_, _36112_, _07966_);
  or (_36114_, _36113_, _36111_);
  nor (_36115_, _14940_, _07988_);
  and (_36116_, _14940_, _07988_);
  nor (_36117_, _36116_, _36115_);
  and (_36119_, _36117_, _15714_);
  nor (_36120_, _36117_, _15714_);
  nor (_36121_, _36120_, _36119_);
  and (_36122_, _36121_, _16019_);
  nor (_36123_, _36121_, _16019_);
  nor (_36124_, _36123_, _36122_);
  nor (_36125_, _36124_, _16355_);
  and (_36126_, _36124_, _16355_);
  or (_36127_, _36126_, _36125_);
  nor (_36128_, _36127_, _16684_);
  and (_36130_, _36127_, _16684_);
  or (_36131_, _36130_, _36128_);
  and (_36132_, _36131_, _17017_);
  nor (_36133_, _36131_, _17017_);
  or (_36134_, _36133_, _36132_);
  or (_36135_, _36134_, _08004_);
  nand (_36136_, _36134_, _08004_);
  and (_36137_, _36136_, _36135_);
  or (_36138_, _36137_, _10004_);
  and (_36139_, _36138_, _09989_);
  and (_36141_, _36139_, _36114_);
  nor (_36142_, _15408_, _35636_);
  nor (_36143_, _36142_, _35637_);
  nor (_36144_, _36143_, _15719_);
  and (_36145_, _36143_, _15719_);
  or (_36146_, _36145_, _36144_);
  nor (_36147_, _36146_, _16025_);
  and (_36148_, _36146_, _16025_);
  nor (_36149_, _36148_, _36147_);
  nor (_36150_, _36149_, _16360_);
  and (_36152_, _36149_, _16360_);
  or (_36153_, _36152_, _36150_);
  nor (_36154_, _36153_, _16690_);
  and (_36155_, _36153_, _16690_);
  nor (_36156_, _36155_, _36154_);
  nor (_36157_, _36156_, _17023_);
  and (_36158_, _36156_, _17023_);
  or (_36159_, _36158_, _36157_);
  or (_36160_, _36159_, _08727_);
  nand (_36161_, _36159_, _08727_);
  and (_36163_, _36161_, _03709_);
  and (_36164_, _36163_, _36160_);
  nor (_36165_, _15413_, _10442_);
  nor (_36166_, _36165_, _35662_);
  nor (_36167_, _36166_, _15724_);
  and (_36168_, _36166_, _15724_);
  or (_36169_, _36168_, _36167_);
  nor (_36170_, _36169_, _16031_);
  and (_36171_, _36169_, _16031_);
  or (_36172_, _36171_, _36170_);
  nor (_36174_, _36172_, _16366_);
  and (_36175_, _36172_, _16366_);
  or (_36176_, _36175_, _36174_);
  and (_36177_, _36176_, _16696_);
  nor (_36178_, _36176_, _16696_);
  nor (_36179_, _36178_, _36177_);
  and (_36180_, _36179_, _17028_);
  nor (_36181_, _36179_, _17028_);
  or (_36182_, _36181_, _36180_);
  and (_36183_, _36182_, _08766_);
  nor (_36185_, _36182_, _08766_);
  or (_36186_, _36185_, _36183_);
  nand (_36187_, _36186_, _08691_);
  and (_36188_, _03850_, _03254_);
  not (_36189_, _36188_);
  nor (_36190_, _07964_, _03707_);
  and (_36191_, _36190_, _36189_);
  and (_36192_, _36191_, _29074_);
  nand (_36193_, _36192_, _36187_);
  or (_36194_, _36193_, _36164_);
  or (_36196_, _36194_, _36141_);
  and (_36197_, _03862_, _03254_);
  nor (_36198_, _36192_, _34829_);
  nor (_36199_, _36198_, _36197_);
  and (_36200_, _36199_, _36196_);
  nand (_36201_, _34829_, _36197_);
  and (_36202_, _04927_, _04728_);
  nand (_36203_, _36202_, _36201_);
  or (_36204_, _36203_, _36200_);
  or (_36205_, _36202_, _34829_);
  and (_36207_, _36205_, _03704_);
  and (_36208_, _36207_, _36204_);
  and (_36209_, _35001_, _03703_);
  or (_36210_, _36209_, _08772_);
  or (_36211_, _36210_, _36208_);
  not (_36212_, _08778_);
  and (_36213_, _15477_, _36212_);
  and (_36214_, _36213_, \oc8051_golden_model_1.ACC [3]);
  nor (_36215_, _36213_, \oc8051_golden_model_1.ACC [3]);
  nor (_36216_, _36215_, _36214_);
  and (_36218_, _36216_, _16379_);
  nor (_36219_, _36216_, _16379_);
  nor (_36220_, _36219_, _36218_);
  and (_36221_, _16707_, _07586_);
  nor (_36222_, _16707_, _07586_);
  nor (_36223_, _36222_, _36221_);
  nor (_36224_, _36223_, _36220_);
  and (_36225_, _36223_, _36220_);
  or (_36226_, _36225_, _36224_);
  nor (_36227_, _36226_, _08784_);
  and (_36229_, _36226_, _08784_);
  nor (_36230_, _36229_, _36227_);
  nand (_36231_, _36230_, _08772_);
  and (_36232_, _36231_, _11972_);
  and (_36233_, _36232_, _36211_);
  and (_36234_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_36235_, _36234_, _08142_);
  nand (_36236_, _36235_, _36070_);
  or (_36237_, _36235_, _36070_);
  and (_36238_, _36237_, _36236_);
  nand (_36240_, _36238_, _08777_);
  nand (_36241_, _36240_, _04735_);
  or (_36242_, _36241_, _36233_);
  and (_36243_, _36242_, _34831_);
  or (_36244_, _36243_, _03384_);
  or (_36245_, _35151_, _03385_);
  and (_36246_, _36245_, _12377_);
  and (_36247_, _36246_, _36244_);
  or (_36248_, _36247_, _34830_);
  and (_36249_, _04110_, _03398_);
  not (_36251_, _36249_);
  and (_36252_, _06909_, _04925_);
  and (_36253_, _36252_, _36251_);
  and (_36254_, _36253_, _36248_);
  not (_36255_, _36253_);
  nand (_36256_, _36255_, _34829_);
  nand (_36257_, _36256_, _04947_);
  or (_36258_, _36257_, _36254_);
  or (_36259_, _34829_, _04947_);
  and (_36260_, _36259_, _03702_);
  and (_36262_, _36260_, _36258_);
  not (_36263_, _16053_);
  nor (_36264_, _15433_, _14985_);
  and (_36265_, _15433_, _14985_);
  nor (_36266_, _36265_, _36264_);
  nor (_36267_, _36266_, _15746_);
  and (_36268_, _36266_, _15746_);
  nor (_36269_, _36268_, _36267_);
  nor (_36270_, _36269_, _36263_);
  and (_36271_, _36269_, _36263_);
  or (_36273_, _36271_, _36270_);
  and (_36274_, _36273_, _16391_);
  nor (_36275_, _36273_, _16391_);
  or (_36276_, _36275_, _36274_);
  and (_36277_, _36276_, _16720_);
  nor (_36278_, _36276_, _16720_);
  or (_36279_, _36278_, _36277_);
  and (_36280_, _36279_, _17051_);
  nor (_36281_, _36279_, _17051_);
  or (_36282_, _36281_, _36280_);
  and (_36284_, _36282_, _08797_);
  nor (_36285_, _36282_, _08797_);
  or (_36286_, _36285_, _36284_);
  and (_36287_, _36286_, _03701_);
  or (_36288_, _36287_, _08794_);
  or (_36289_, _36288_, _36262_);
  not (_36290_, _08802_);
  and (_36291_, _15477_, _36290_);
  and (_36292_, _36291_, _07734_);
  nor (_36293_, _36291_, _07734_);
  nor (_36295_, _36293_, _36292_);
  nor (_36296_, _36295_, _16397_);
  and (_36297_, _36295_, _16397_);
  or (_36298_, _36297_, _36296_);
  nor (_36299_, _36298_, _17057_);
  and (_36300_, _36298_, _17057_);
  or (_36301_, _36300_, _36299_);
  nor (_36302_, _16726_, _08809_);
  and (_36303_, _16726_, _08809_);
  nor (_36304_, _36303_, _36302_);
  nand (_36306_, _36304_, _36301_);
  or (_36307_, _36304_, _36301_);
  nand (_36308_, _36307_, _36306_);
  nand (_36309_, _36308_, _08794_);
  and (_36310_, _36309_, _36289_);
  or (_36311_, _36310_, _08801_);
  not (_36312_, _08801_);
  or (_36313_, _34829_, _36312_);
  and (_36314_, _36313_, _10921_);
  and (_36315_, _36314_, _36311_);
  nand (_36317_, _34829_, _03841_);
  nand (_36318_, _36317_, _28781_);
  or (_36319_, _36318_, _36315_);
  or (_36320_, _34829_, _28781_);
  and (_36321_, _36320_, _42908_);
  and (_36322_, _36321_, _36319_);
  or (_36323_, _36322_, _34813_);
  and (_43331_, _36323_, _41654_);
  not (_36324_, \oc8051_golden_model_1.PSW [1]);
  nor (_36325_, _42908_, _36324_);
  nor (_36327_, _05360_, _36324_);
  and (_36328_, _05360_, _04813_);
  or (_36329_, _36328_, _36327_);
  or (_36330_, _36329_, _04537_);
  or (_36331_, _05360_, \oc8051_golden_model_1.PSW [1]);
  and (_36332_, _12225_, _05360_);
  not (_36333_, _36332_);
  and (_36334_, _36333_, _36331_);
  or (_36335_, _36334_, _04630_);
  and (_36336_, _05360_, \oc8051_golden_model_1.ACC [1]);
  or (_36338_, _36336_, _36327_);
  and (_36339_, _36338_, _04615_);
  nor (_36340_, _04615_, _36324_);
  or (_36341_, _36340_, _03757_);
  or (_36342_, _36341_, _36339_);
  and (_36343_, _36342_, _03697_);
  and (_36344_, _36343_, _36335_);
  nor (_36345_, _06092_, _36324_);
  and (_36346_, _12212_, _06092_);
  or (_36347_, _36346_, _36345_);
  and (_36349_, _36347_, _03696_);
  or (_36350_, _36349_, _03755_);
  or (_36351_, _36350_, _36344_);
  and (_36352_, _36351_, _36330_);
  or (_36353_, _36352_, _03750_);
  or (_36354_, _36338_, _03751_);
  and (_36355_, _36354_, _03692_);
  and (_36356_, _36355_, _36353_);
  and (_36357_, _12200_, _06092_);
  or (_36358_, _36357_, _36345_);
  and (_36360_, _36358_, _03691_);
  or (_36361_, _36360_, _03684_);
  or (_36362_, _36361_, _36356_);
  and (_36363_, _36346_, _12211_);
  or (_36364_, _36345_, _03685_);
  or (_36365_, _36364_, _36363_);
  and (_36366_, _36365_, _36362_);
  and (_36367_, _36366_, _03680_);
  not (_36368_, _06092_);
  nor (_36369_, _12256_, _36368_);
  or (_36371_, _36345_, _36369_);
  and (_36372_, _36371_, _03679_);
  or (_36373_, _36372_, _07544_);
  or (_36374_, _36373_, _36367_);
  or (_36375_, _36329_, _06994_);
  and (_36376_, _36375_, _36374_);
  or (_36377_, _36376_, _04678_);
  and (_36378_, _06934_, _05360_);
  or (_36379_, _36378_, _36327_);
  or (_36380_, _36379_, _04679_);
  and (_36382_, _36380_, _03415_);
  and (_36383_, _36382_, _36377_);
  nand (_36384_, _12313_, _05360_);
  and (_36385_, _36331_, _07559_);
  and (_36386_, _36385_, _36384_);
  or (_36387_, _36386_, _36383_);
  and (_36388_, _36387_, _03840_);
  or (_36389_, _12207_, _11659_);
  and (_36390_, _36331_, _03838_);
  and (_36391_, _36390_, _36389_);
  nand (_36393_, _05360_, _04515_);
  and (_36394_, _36393_, _03839_);
  and (_36395_, _36394_, _36331_);
  or (_36396_, _36395_, _03959_);
  or (_36397_, _36396_, _36391_);
  or (_36398_, _36397_, _36388_);
  nor (_36399_, _08710_, _11659_);
  or (_36400_, _36399_, _36327_);
  nand (_36401_, _08709_, _05360_);
  and (_36402_, _36401_, _36400_);
  or (_36404_, _36402_, _04701_);
  and (_36405_, _36404_, _04708_);
  and (_36406_, _36405_, _36398_);
  or (_36407_, _12206_, _11659_);
  and (_36408_, _36331_, _03866_);
  and (_36409_, _36408_, _36407_);
  or (_36410_, _36409_, _03967_);
  or (_36411_, _36410_, _36406_);
  nor (_36412_, _36327_, _04706_);
  nand (_36413_, _36412_, _36401_);
  and (_36415_, _36413_, _06532_);
  and (_36416_, _36415_, _36411_);
  or (_36417_, _36393_, _05603_);
  and (_36418_, _36417_, _03835_);
  and (_36419_, _36418_, _36331_);
  or (_36420_, _36419_, _03954_);
  or (_36421_, _36420_, _36416_);
  or (_36422_, _36400_, _06537_);
  and (_36423_, _36422_, _36421_);
  or (_36424_, _36423_, _03703_);
  or (_36426_, _36334_, _03704_);
  and (_36427_, _36426_, _03385_);
  and (_36428_, _36427_, _36424_);
  and (_36429_, _36358_, _03384_);
  or (_36430_, _36429_, _03701_);
  or (_36431_, _36430_, _36428_);
  or (_36432_, _36327_, _03702_);
  or (_36433_, _36432_, _36332_);
  and (_36434_, _36433_, _42908_);
  and (_36435_, _36434_, _36431_);
  or (_36437_, _36435_, _36325_);
  and (_43332_, _36437_, _41654_);
  and (_36438_, _42912_, \oc8051_golden_model_1.PSW [2]);
  nor (_36439_, _08001_, _11952_);
  and (_36440_, _08001_, _07968_);
  or (_36441_, _36440_, _36439_);
  and (_36442_, _36441_, _07966_);
  and (_36443_, _11659_, \oc8051_golden_model_1.PSW [2]);
  nor (_36444_, _11659_, _05236_);
  or (_36445_, _36444_, _36443_);
  or (_36447_, _36445_, _06994_);
  and (_36448_, _11856_, _08367_);
  nor (_36449_, _11856_, _08367_);
  nor (_36450_, _36449_, _36448_);
  and (_36451_, _36450_, _08422_);
  nor (_36452_, _36450_, _08422_);
  or (_36453_, _36452_, _36451_);
  and (_36454_, _36453_, _08287_);
  and (_36455_, _08188_, \oc8051_golden_model_1.ACC [7]);
  nor (_36456_, _08188_, \oc8051_golden_model_1.ACC [7]);
  or (_36458_, _36456_, _36455_);
  and (_36459_, _36458_, _11821_);
  nor (_36460_, _36458_, _11821_);
  nor (_36461_, _36460_, _36459_);
  and (_36462_, _36461_, _08258_);
  nor (_36463_, _36461_, _08258_);
  or (_36464_, _36463_, _36462_);
  or (_36465_, _36464_, _08181_);
  or (_36466_, _36445_, _04537_);
  nor (_36467_, _12427_, _11659_);
  or (_36469_, _36467_, _36443_);
  or (_36470_, _36469_, _04630_);
  and (_36471_, _05360_, \oc8051_golden_model_1.ACC [2]);
  or (_36472_, _36471_, _36443_);
  and (_36473_, _36472_, _04615_);
  and (_36474_, _04616_, \oc8051_golden_model_1.PSW [2]);
  or (_36475_, _36474_, _03757_);
  or (_36476_, _36475_, _36473_);
  and (_36477_, _36476_, _03697_);
  and (_36478_, _36477_, _36470_);
  and (_36480_, _36368_, \oc8051_golden_model_1.PSW [2]);
  and (_36481_, _12419_, _06092_);
  or (_36482_, _36481_, _36480_);
  and (_36483_, _36482_, _03696_);
  or (_36484_, _36483_, _03755_);
  or (_36485_, _36484_, _36478_);
  and (_36486_, _36485_, _36466_);
  or (_36487_, _36486_, _03750_);
  or (_36488_, _36472_, _03751_);
  and (_36489_, _36488_, _03692_);
  and (_36491_, _36489_, _36487_);
  and (_36492_, _12422_, _06092_);
  or (_36493_, _36492_, _36480_);
  and (_36494_, _36493_, _03691_);
  or (_36495_, _36494_, _03684_);
  or (_36496_, _36495_, _36491_);
  and (_36497_, _36481_, _12418_);
  or (_36498_, _36480_, _03685_);
  or (_36499_, _36498_, _36497_);
  and (_36500_, _36499_, _07030_);
  and (_36502_, _36500_, _36496_);
  or (_36503_, _14286_, _14171_);
  or (_36504_, _36503_, _14394_);
  or (_36505_, _36504_, _14513_);
  or (_36506_, _36505_, _14629_);
  or (_36507_, _36506_, _14746_);
  or (_36508_, _36507_, _07540_);
  or (_36509_, _36508_, _14863_);
  and (_36510_, _36509_, _07024_);
  or (_36511_, _36510_, _08182_);
  or (_36513_, _36511_, _36502_);
  and (_36514_, _36513_, _08261_);
  and (_36515_, _36514_, _36465_);
  or (_36516_, _36515_, _03818_);
  nor (_36517_, _08009_, \oc8051_golden_model_1.ACC [7]);
  and (_36518_, _08009_, \oc8051_golden_model_1.ACC [7]);
  nor (_36519_, _36518_, _36517_);
  not (_36520_, _36519_);
  nor (_36521_, _36520_, _11833_);
  and (_36522_, _36520_, _11833_);
  or (_36524_, _36522_, _36521_);
  nor (_36525_, _36524_, _08283_);
  and (_36526_, _36524_, _08283_);
  or (_36527_, _36526_, _36525_);
  and (_36528_, _36527_, _08260_);
  or (_36529_, _36528_, _36516_);
  not (_36530_, _08355_);
  not (_36531_, _08293_);
  nor (_36532_, _11846_, _36531_);
  and (_36533_, _11846_, _36531_);
  nor (_36535_, _36533_, _36532_);
  nor (_36536_, _36535_, _36530_);
  and (_36537_, _36535_, _36530_);
  or (_36538_, _36537_, _03823_);
  or (_36539_, _36538_, _36536_);
  and (_36540_, _36539_, _08288_);
  and (_36541_, _36540_, _36529_);
  or (_36542_, _36541_, _36454_);
  and (_36543_, _36542_, _03680_);
  nor (_36544_, _12465_, _36368_);
  or (_36546_, _36544_, _36480_);
  and (_36547_, _36546_, _03679_);
  or (_36548_, _36547_, _07544_);
  or (_36549_, _36548_, _36543_);
  and (_36550_, _36549_, _36447_);
  or (_36551_, _36550_, _04678_);
  and (_36552_, _06938_, _05360_);
  or (_36553_, _36552_, _36443_);
  or (_36554_, _36553_, _04679_);
  and (_36555_, _36554_, _36551_);
  or (_36557_, _36555_, _07559_);
  nor (_36558_, _12523_, _11659_);
  or (_36559_, _36443_, _03415_);
  or (_36560_, _36559_, _36558_);
  and (_36561_, _36560_, _07565_);
  and (_36562_, _36561_, _36557_);
  nor (_36563_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and (_36564_, _36563_, _07585_);
  nand (_36565_, _36564_, _07558_);
  nand (_36566_, _36565_, _03840_);
  or (_36568_, _36566_, _36562_);
  and (_36569_, _12537_, _05360_);
  or (_36570_, _36443_, _04703_);
  or (_36571_, _36570_, _36569_);
  and (_36572_, _05360_, _06457_);
  or (_36573_, _36572_, _36443_);
  or (_36574_, _36573_, _04694_);
  and (_36575_, _36574_, _04701_);
  and (_36576_, _36575_, _36571_);
  and (_36577_, _36576_, _36568_);
  and (_36579_, _08707_, _05360_);
  or (_36580_, _36579_, _36443_);
  and (_36581_, _36580_, _03959_);
  or (_36582_, _36581_, _36577_);
  and (_36583_, _36582_, _04708_);
  or (_36584_, _36443_, _05700_);
  and (_36585_, _36573_, _03866_);
  and (_36586_, _36585_, _36584_);
  or (_36587_, _36586_, _36583_);
  and (_36588_, _36587_, _04706_);
  and (_36590_, _36472_, _03967_);
  and (_36591_, _36590_, _36584_);
  or (_36592_, _36591_, _03835_);
  or (_36593_, _36592_, _36588_);
  nor (_36594_, _12536_, _11659_);
  or (_36595_, _36443_, _06532_);
  or (_36596_, _36595_, _36594_);
  and (_36597_, _36596_, _06537_);
  and (_36598_, _36597_, _36593_);
  nor (_36599_, _08706_, _11659_);
  or (_36601_, _36599_, _36443_);
  and (_36602_, _36601_, _03954_);
  or (_36603_, _36602_, _08543_);
  or (_36604_, _36603_, _36598_);
  nor (_36605_, _36458_, _11913_);
  nor (_36606_, _36605_, _36455_);
  and (_36607_, _36606_, _08571_);
  and (_36608_, _36455_, _08568_);
  or (_36609_, _36608_, _36607_);
  or (_36610_, _36609_, _08542_);
  and (_36612_, _36610_, _08546_);
  and (_36613_, _36612_, _36604_);
  and (_36614_, _36609_, _04374_);
  or (_36615_, _36614_, _36613_);
  and (_36616_, _36615_, _34833_);
  and (_36617_, _36518_, _08075_);
  nor (_36618_, _36520_, _11924_);
  nor (_36619_, _36618_, _36518_);
  and (_36620_, _36619_, _08078_);
  or (_36621_, _36620_, _36617_);
  and (_36623_, _36621_, _34832_);
  or (_36624_, _36623_, _36616_);
  and (_36625_, _36624_, _04372_);
  and (_36626_, _36621_, _04371_);
  or (_36627_, _36626_, _03963_);
  or (_36628_, _36627_, _36625_);
  and (_36629_, _08292_, \oc8051_golden_model_1.ACC [7]);
  and (_36630_, _36629_, _08602_);
  nor (_36631_, _08292_, \oc8051_golden_model_1.ACC [7]);
  nor (_36632_, _36631_, _11929_);
  nor (_36634_, _36632_, _36629_);
  and (_36635_, _36634_, _08605_);
  or (_36636_, _36635_, _36630_);
  or (_36637_, _36636_, _03964_);
  and (_36638_, _36637_, _08581_);
  and (_36639_, _36638_, _36628_);
  and (_36640_, _08366_, \oc8051_golden_model_1.ACC [7]);
  nor (_36641_, _08366_, \oc8051_golden_model_1.ACC [7]);
  nor (_36642_, _36641_, _11935_);
  nor (_36643_, _36642_, _36640_);
  and (_36645_, _36643_, _08632_);
  and (_36646_, _36640_, _08629_);
  or (_36647_, _36646_, _36645_);
  and (_36648_, _36647_, _08580_);
  or (_36649_, _36648_, _15145_);
  or (_36650_, _36649_, _36639_);
  and (_36651_, _08679_, _08467_);
  nor (_36652_, _08679_, _11944_);
  or (_36653_, _36652_, _36651_);
  or (_36654_, _36653_, _10007_);
  and (_36656_, _36654_, _10004_);
  and (_36657_, _36656_, _36650_);
  or (_36658_, _36657_, _36442_);
  and (_36659_, _36658_, _09989_);
  or (_36660_, _08724_, _06522_);
  and (_36661_, _11962_, _36660_);
  nand (_36662_, _08763_, _11966_);
  and (_36663_, _36662_, _11968_);
  or (_36664_, _36663_, _03703_);
  or (_36665_, _36664_, _36661_);
  or (_36667_, _36665_, _36659_);
  or (_36668_, _36469_, _03704_);
  and (_36669_, _36668_, _03385_);
  and (_36670_, _36669_, _36667_);
  and (_36671_, _36493_, _03384_);
  or (_36672_, _36671_, _03701_);
  or (_36673_, _36672_, _36670_);
  and (_36674_, _12596_, _05360_);
  or (_36675_, _36443_, _03702_);
  or (_36676_, _36675_, _36674_);
  and (_36678_, _36676_, _42908_);
  and (_36679_, _36678_, _36673_);
  or (_36680_, _36679_, _36438_);
  and (_43333_, _36680_, _41654_);
  nor (_36681_, _42908_, _05064_);
  nor (_36682_, _05360_, _05064_);
  nor (_36683_, _11659_, _05050_);
  or (_36684_, _36683_, _36682_);
  or (_36685_, _36684_, _06994_);
  nor (_36686_, _12610_, _11659_);
  or (_36688_, _36686_, _36682_);
  or (_36689_, _36688_, _04630_);
  and (_36690_, _05360_, \oc8051_golden_model_1.ACC [3]);
  or (_36691_, _36690_, _36682_);
  and (_36692_, _36691_, _04615_);
  nor (_36693_, _04615_, _05064_);
  or (_36694_, _36693_, _03757_);
  or (_36695_, _36694_, _36692_);
  and (_36696_, _36695_, _03697_);
  and (_36697_, _36696_, _36689_);
  nor (_36699_, _06092_, _05064_);
  and (_36700_, _12619_, _06092_);
  or (_36701_, _36700_, _36699_);
  and (_36702_, _36701_, _03696_);
  or (_36703_, _36702_, _03755_);
  or (_36704_, _36703_, _36697_);
  or (_36705_, _36684_, _04537_);
  and (_36706_, _36705_, _36704_);
  or (_36707_, _36706_, _03750_);
  or (_36708_, _36691_, _03751_);
  and (_36710_, _36708_, _03692_);
  and (_36711_, _36710_, _36707_);
  and (_36712_, _12622_, _06092_);
  or (_36713_, _36712_, _36699_);
  and (_36714_, _36713_, _03691_);
  or (_36715_, _36714_, _03684_);
  or (_36716_, _36715_, _36711_);
  or (_36717_, _36699_, _12618_);
  and (_36718_, _36717_, _36701_);
  or (_36719_, _36718_, _03685_);
  and (_36721_, _36719_, _03680_);
  and (_36722_, _36721_, _36716_);
  nor (_36723_, _12665_, _36368_);
  or (_36724_, _36723_, _36699_);
  and (_36725_, _36724_, _03679_);
  or (_36726_, _36725_, _07544_);
  or (_36727_, _36726_, _36722_);
  and (_36728_, _36727_, _36685_);
  or (_36729_, _36728_, _04678_);
  and (_36730_, _06937_, _05360_);
  or (_36732_, _36682_, _04679_);
  or (_36733_, _36732_, _36730_);
  and (_36734_, _36733_, _36729_);
  or (_36735_, _36734_, _07559_);
  nor (_36736_, _12724_, _11659_);
  or (_36737_, _36682_, _03415_);
  or (_36738_, _36737_, _36736_);
  and (_36739_, _36738_, _04694_);
  and (_36740_, _36739_, _36735_);
  and (_36741_, _05360_, _06415_);
  or (_36743_, _36741_, _36682_);
  and (_36744_, _36743_, _03839_);
  or (_36745_, _36744_, _03838_);
  or (_36746_, _36745_, _36740_);
  and (_36747_, _12738_, _05360_);
  or (_36748_, _36682_, _04703_);
  or (_36749_, _36748_, _36747_);
  and (_36750_, _36749_, _04701_);
  and (_36751_, _36750_, _36746_);
  and (_36752_, _10455_, _05360_);
  or (_36754_, _36752_, _36682_);
  and (_36755_, _36754_, _03959_);
  or (_36756_, _36755_, _36751_);
  and (_36757_, _36756_, _04708_);
  or (_36758_, _36682_, _05554_);
  and (_36759_, _36743_, _03866_);
  and (_36760_, _36759_, _36758_);
  or (_36761_, _36760_, _36757_);
  and (_36762_, _36761_, _04706_);
  and (_36763_, _36691_, _03967_);
  and (_36765_, _36763_, _36758_);
  or (_36766_, _36765_, _03835_);
  or (_36767_, _36766_, _36762_);
  nor (_36768_, _12737_, _11659_);
  or (_36769_, _36682_, _06532_);
  or (_36770_, _36769_, _36768_);
  and (_36771_, _36770_, _06537_);
  and (_36772_, _36771_, _36767_);
  nor (_36773_, _08701_, _11659_);
  or (_36774_, _36773_, _36682_);
  and (_36776_, _36774_, _03954_);
  or (_36777_, _36776_, _03703_);
  or (_36778_, _36777_, _36772_);
  or (_36779_, _36688_, _03704_);
  and (_36780_, _36779_, _03385_);
  and (_36781_, _36780_, _36778_);
  and (_36782_, _36713_, _03384_);
  or (_36783_, _36782_, _03701_);
  or (_36784_, _36783_, _36781_);
  and (_36785_, _12792_, _05360_);
  or (_36787_, _36682_, _03702_);
  or (_36788_, _36787_, _36785_);
  and (_36789_, _36788_, _42908_);
  and (_36790_, _36789_, _36784_);
  or (_36791_, _36790_, _36681_);
  and (_43334_, _36791_, _41654_);
  and (_36792_, _42912_, \oc8051_golden_model_1.PSW [4]);
  and (_36793_, _11659_, \oc8051_golden_model_1.PSW [4]);
  nor (_36794_, _05898_, _11659_);
  or (_36795_, _36794_, _36793_);
  or (_36797_, _36795_, _06994_);
  and (_36798_, _36368_, \oc8051_golden_model_1.PSW [4]);
  and (_36799_, _12808_, _06092_);
  or (_36800_, _36799_, _36798_);
  and (_36801_, _36800_, _03691_);
  nor (_36802_, _12828_, _11659_);
  or (_36803_, _36802_, _36793_);
  or (_36804_, _36803_, _04630_);
  and (_36805_, _05360_, \oc8051_golden_model_1.ACC [4]);
  or (_36806_, _36805_, _36793_);
  and (_36808_, _36806_, _04615_);
  and (_36809_, _04616_, \oc8051_golden_model_1.PSW [4]);
  or (_36810_, _36809_, _03757_);
  or (_36811_, _36810_, _36808_);
  and (_36812_, _36811_, _03697_);
  and (_36813_, _36812_, _36804_);
  and (_36814_, _12832_, _06092_);
  or (_36815_, _36814_, _36798_);
  and (_36816_, _36815_, _03696_);
  or (_36817_, _36816_, _03755_);
  or (_36819_, _36817_, _36813_);
  or (_36820_, _36795_, _04537_);
  and (_36821_, _36820_, _36819_);
  or (_36822_, _36821_, _03750_);
  or (_36823_, _36806_, _03751_);
  and (_36824_, _36823_, _03692_);
  and (_36825_, _36824_, _36822_);
  or (_36826_, _36825_, _36801_);
  and (_36827_, _36826_, _03685_);
  and (_36828_, _12848_, _06092_);
  or (_36830_, _36828_, _36798_);
  and (_36831_, _36830_, _03684_);
  or (_36832_, _36831_, _36827_);
  and (_36833_, _36832_, _03680_);
  nor (_36834_, _12810_, _36368_);
  or (_36835_, _36834_, _36798_);
  and (_36836_, _36835_, _03679_);
  or (_36837_, _36836_, _07544_);
  or (_36838_, _36837_, _36833_);
  and (_36839_, _36838_, _36797_);
  or (_36841_, _36839_, _04678_);
  and (_36842_, _06942_, _05360_);
  or (_36843_, _36842_, _36793_);
  or (_36844_, _36843_, _04679_);
  and (_36845_, _36844_, _36841_);
  or (_36846_, _36845_, _07559_);
  nor (_36847_, _12919_, _11659_);
  or (_36848_, _36793_, _03415_);
  or (_36849_, _36848_, _36847_);
  and (_36850_, _36849_, _04694_);
  and (_36852_, _36850_, _36846_);
  and (_36853_, _06422_, _05360_);
  or (_36854_, _36853_, _36793_);
  and (_36855_, _36854_, _03839_);
  or (_36856_, _36855_, _03838_);
  or (_36857_, _36856_, _36852_);
  and (_36858_, _12933_, _05360_);
  or (_36859_, _36793_, _04703_);
  or (_36860_, _36859_, _36858_);
  and (_36861_, _36860_, _04701_);
  and (_36863_, _36861_, _36857_);
  and (_36864_, _08700_, _05360_);
  or (_36865_, _36864_, _36793_);
  and (_36866_, _36865_, _03959_);
  or (_36867_, _36866_, _36863_);
  and (_36868_, _36867_, _04708_);
  or (_36869_, _36793_, _08303_);
  and (_36870_, _36854_, _03866_);
  and (_36871_, _36870_, _36869_);
  or (_36872_, _36871_, _36868_);
  and (_36874_, _36872_, _04706_);
  and (_36875_, _36806_, _03967_);
  and (_36876_, _36875_, _36869_);
  or (_36877_, _36876_, _03835_);
  or (_36878_, _36877_, _36874_);
  nor (_36879_, _12931_, _11659_);
  or (_36880_, _36793_, _06532_);
  or (_36881_, _36880_, _36879_);
  and (_36882_, _36881_, _06537_);
  and (_36883_, _36882_, _36878_);
  nor (_36885_, _08699_, _11659_);
  or (_36886_, _36885_, _36793_);
  and (_36887_, _36886_, _03954_);
  or (_36888_, _36887_, _03703_);
  or (_36889_, _36888_, _36883_);
  or (_36890_, _36803_, _03704_);
  and (_36891_, _36890_, _03385_);
  and (_36892_, _36891_, _36889_);
  and (_36893_, _36800_, _03384_);
  or (_36894_, _36893_, _03701_);
  or (_36896_, _36894_, _36892_);
  and (_36897_, _12991_, _05360_);
  or (_36898_, _36793_, _03702_);
  or (_36899_, _36898_, _36897_);
  and (_36900_, _36899_, _42908_);
  and (_36901_, _36900_, _36896_);
  or (_36902_, _36901_, _36792_);
  and (_43335_, _36902_, _41654_);
  and (_36903_, _42912_, \oc8051_golden_model_1.PSW [5]);
  and (_36904_, _11659_, \oc8051_golden_model_1.PSW [5]);
  nor (_36906_, _05799_, _11659_);
  or (_36907_, _36906_, _36904_);
  or (_36908_, _36907_, _06994_);
  nor (_36909_, _13025_, _11659_);
  or (_36910_, _36909_, _36904_);
  or (_36911_, _36910_, _04630_);
  and (_36912_, _05360_, \oc8051_golden_model_1.ACC [5]);
  or (_36913_, _36912_, _36904_);
  and (_36914_, _36913_, _04615_);
  and (_36915_, _04616_, \oc8051_golden_model_1.PSW [5]);
  or (_36917_, _36915_, _03757_);
  or (_36918_, _36917_, _36914_);
  and (_36919_, _36918_, _03697_);
  and (_36920_, _36919_, _36911_);
  and (_36921_, _36368_, \oc8051_golden_model_1.PSW [5]);
  and (_36922_, _13029_, _06092_);
  or (_36923_, _36922_, _36921_);
  and (_36924_, _36923_, _03696_);
  or (_36925_, _36924_, _03755_);
  or (_36926_, _36925_, _36920_);
  or (_36928_, _36907_, _04537_);
  and (_36929_, _36928_, _36926_);
  or (_36930_, _36929_, _03750_);
  or (_36931_, _36913_, _03751_);
  and (_36932_, _36931_, _03692_);
  and (_36933_, _36932_, _36930_);
  and (_36934_, _13007_, _06092_);
  or (_36935_, _36934_, _36921_);
  and (_36936_, _36935_, _03691_);
  or (_36937_, _36936_, _03684_);
  or (_36939_, _36937_, _36933_);
  or (_36940_, _36921_, _13044_);
  and (_36941_, _36940_, _36923_);
  or (_36942_, _36941_, _03685_);
  and (_36943_, _36942_, _03680_);
  and (_36944_, _36943_, _36939_);
  nor (_36945_, _13009_, _36368_);
  or (_36946_, _36945_, _36921_);
  and (_36947_, _36946_, _03679_);
  or (_36948_, _36947_, _07544_);
  or (_36950_, _36948_, _36944_);
  and (_36951_, _36950_, _36908_);
  or (_36952_, _36951_, _04678_);
  and (_36953_, _06941_, _05360_);
  or (_36954_, _36953_, _36904_);
  or (_36955_, _36954_, _04679_);
  and (_36956_, _36955_, _36952_);
  or (_36957_, _36956_, _07559_);
  nor (_36958_, _13118_, _11659_);
  or (_36959_, _36904_, _03415_);
  or (_36961_, _36959_, _36958_);
  and (_36962_, _36961_, _04694_);
  and (_36963_, _36962_, _36957_);
  and (_36964_, _06371_, _05360_);
  or (_36965_, _36964_, _36904_);
  and (_36966_, _36965_, _03839_);
  or (_36967_, _36966_, _03838_);
  or (_36968_, _36967_, _36963_);
  and (_36969_, _13133_, _05360_);
  or (_36970_, _36904_, _04703_);
  or (_36972_, _36970_, _36969_);
  and (_36973_, _36972_, _04701_);
  and (_36974_, _36973_, _36968_);
  and (_36975_, _10451_, _05360_);
  or (_36976_, _36975_, _36904_);
  and (_36977_, _36976_, _03959_);
  or (_36978_, _36977_, _36974_);
  and (_36979_, _36978_, _04708_);
  or (_36980_, _36904_, _08302_);
  and (_36981_, _36965_, _03866_);
  and (_36983_, _36981_, _36980_);
  or (_36984_, _36983_, _36979_);
  and (_36985_, _36984_, _04706_);
  and (_36986_, _36913_, _03967_);
  and (_36987_, _36986_, _36980_);
  or (_36988_, _36987_, _03835_);
  or (_36989_, _36988_, _36985_);
  nor (_36990_, _13131_, _11659_);
  or (_36991_, _36904_, _06532_);
  or (_36992_, _36991_, _36990_);
  and (_36994_, _36992_, _06537_);
  and (_36995_, _36994_, _36989_);
  nor (_36996_, _08697_, _11659_);
  or (_36997_, _36996_, _36904_);
  and (_36998_, _36997_, _03954_);
  or (_36999_, _36998_, _03703_);
  or (_37000_, _36999_, _36995_);
  or (_37001_, _36910_, _03704_);
  and (_37002_, _37001_, _03385_);
  and (_37003_, _37002_, _37000_);
  and (_37005_, _36935_, _03384_);
  or (_37006_, _37005_, _03701_);
  or (_37007_, _37006_, _37003_);
  and (_37008_, _13193_, _05360_);
  or (_37009_, _36904_, _03702_);
  or (_37010_, _37009_, _37008_);
  and (_37011_, _37010_, _42908_);
  and (_37012_, _37011_, _37007_);
  or (_37013_, _37012_, _36903_);
  and (_43336_, _37013_, _41654_);
  nor (_37015_, _42908_, _15832_);
  or (_37016_, _10007_, _08673_);
  or (_37017_, _08080_, _08031_);
  or (_37018_, _37017_, _08069_);
  or (_37019_, _08562_, _08209_);
  and (_37020_, _04671_, _03473_);
  and (_37021_, _37020_, _37019_);
  nor (_37022_, _13340_, _11659_);
  nor (_37023_, _05360_, _15832_);
  or (_37024_, _37023_, _06532_);
  or (_37026_, _37024_, _37022_);
  nor (_37027_, _06013_, _11659_);
  or (_37028_, _37027_, _37023_);
  or (_37029_, _37028_, _06994_);
  or (_37030_, _08276_, _08031_);
  and (_37031_, _37030_, _08260_);
  nor (_37032_, _06092_, _15832_);
  and (_37033_, _13218_, _06092_);
  or (_37034_, _37033_, _37032_);
  and (_37035_, _37034_, _03691_);
  nor (_37037_, _13234_, _11659_);
  or (_37038_, _37037_, _37023_);
  or (_37039_, _37038_, _04630_);
  and (_37040_, _05360_, \oc8051_golden_model_1.ACC [6]);
  or (_37041_, _37040_, _37023_);
  and (_37042_, _37041_, _04615_);
  nor (_37043_, _04615_, _15832_);
  or (_37044_, _37043_, _03757_);
  or (_37045_, _37044_, _37042_);
  and (_37046_, _37045_, _03697_);
  and (_37048_, _37046_, _37039_);
  and (_37049_, _13238_, _06092_);
  or (_37050_, _37049_, _37032_);
  and (_37051_, _37050_, _03696_);
  or (_37052_, _37051_, _03755_);
  or (_37053_, _37052_, _37048_);
  or (_37054_, _37028_, _04537_);
  and (_37055_, _37054_, _37053_);
  or (_37056_, _37055_, _03750_);
  or (_37057_, _37041_, _03751_);
  and (_37059_, _37057_, _03692_);
  and (_37060_, _37059_, _37056_);
  or (_37061_, _37060_, _37035_);
  and (_37062_, _37061_, _03685_);
  or (_37063_, _37032_, _13253_);
  and (_37064_, _37050_, _03684_);
  and (_37065_, _37064_, _37063_);
  or (_37066_, _37065_, _08182_);
  or (_37067_, _37066_, _37062_);
  or (_37068_, _08209_, _08181_);
  or (_37070_, _37068_, _08245_);
  and (_37071_, _37070_, _08261_);
  and (_37072_, _37071_, _37067_);
  or (_37073_, _37072_, _03818_);
  or (_37074_, _37073_, _37031_);
  or (_37075_, _08345_, _08307_);
  or (_37076_, _37075_, _03823_);
  and (_37077_, _37076_, _37074_);
  or (_37078_, _37077_, _08287_);
  or (_37079_, _08363_, _08288_);
  or (_37081_, _37079_, _08412_);
  and (_37082_, _37081_, _03680_);
  and (_37083_, _37082_, _37078_);
  nor (_37084_, _13220_, _36368_);
  or (_37085_, _37084_, _37032_);
  and (_37086_, _37085_, _03679_);
  or (_37087_, _37086_, _07544_);
  or (_37088_, _37087_, _37083_);
  and (_37089_, _37088_, _37029_);
  or (_37090_, _37089_, _04678_);
  and (_37092_, _06933_, _05360_);
  or (_37093_, _37023_, _04679_);
  or (_37094_, _37093_, _37092_);
  and (_37095_, _37094_, _03415_);
  and (_37096_, _37095_, _37090_);
  nor (_37097_, _13326_, _11659_);
  or (_37098_, _37097_, _37023_);
  and (_37099_, _37098_, _07559_);
  or (_37100_, _37099_, _08854_);
  or (_37101_, _37100_, _37096_);
  and (_37103_, _13341_, _05360_);
  or (_37104_, _37023_, _04703_);
  or (_37105_, _37104_, _37103_);
  and (_37106_, _13333_, _05360_);
  or (_37107_, _37106_, _37023_);
  or (_37108_, _37107_, _04694_);
  and (_37109_, _37108_, _04701_);
  and (_37110_, _37109_, _37105_);
  and (_37111_, _37110_, _37101_);
  and (_37112_, _08695_, _05360_);
  or (_37114_, _37112_, _37023_);
  and (_37115_, _37114_, _03959_);
  or (_37116_, _37115_, _37111_);
  and (_37117_, _37116_, _04708_);
  or (_37118_, _37023_, _08289_);
  and (_37119_, _37107_, _03866_);
  and (_37120_, _37119_, _37118_);
  or (_37121_, _37120_, _37117_);
  and (_37122_, _37121_, _04706_);
  and (_37123_, _37041_, _03967_);
  and (_37125_, _37123_, _37118_);
  or (_37126_, _37125_, _03835_);
  or (_37127_, _37126_, _37122_);
  and (_37128_, _37127_, _37026_);
  or (_37129_, _37128_, _03954_);
  nor (_37130_, _08694_, _11659_);
  or (_37131_, _37130_, _37023_);
  nor (_37132_, _37131_, _06537_);
  nor (_37133_, _37132_, _37020_);
  and (_37134_, _37133_, _37129_);
  nor (_37136_, _37134_, _37021_);
  nor (_37137_, _37136_, _04373_);
  and (_37138_, _03797_, _03473_);
  and (_37139_, _37019_, _04373_);
  or (_37140_, _37139_, _37138_);
  or (_37141_, _37140_, _37137_);
  not (_37142_, _37138_);
  or (_37143_, _37019_, _37142_);
  and (_37144_, _37143_, _37141_);
  or (_37145_, _37144_, _04366_);
  nor (_37147_, _37019_, _04367_);
  nor (_37148_, _37147_, _15126_);
  and (_37149_, _37148_, _37145_);
  and (_37150_, _37019_, _15126_);
  or (_37151_, _37150_, _08079_);
  or (_37152_, _37151_, _37149_);
  and (_37153_, _37152_, _37018_);
  or (_37154_, _37153_, _03963_);
  or (_37155_, _08307_, _03964_);
  or (_37156_, _37155_, _08596_);
  and (_37158_, _37156_, _08581_);
  and (_37159_, _37158_, _37154_);
  or (_37160_, _08623_, _08363_);
  and (_37161_, _37160_, _08580_);
  or (_37162_, _37161_, _15145_);
  or (_37163_, _37162_, _37159_);
  and (_37164_, _37163_, _37016_);
  or (_37165_, _37164_, _07966_);
  or (_37166_, _07995_, _10004_);
  and (_37167_, _37166_, _04166_);
  and (_37169_, _37167_, _37165_);
  and (_37170_, _08718_, _03709_);
  or (_37171_, _37170_, _08691_);
  or (_37172_, _37171_, _37169_);
  or (_37173_, _08757_, _08692_);
  and (_37174_, _37173_, _37172_);
  or (_37175_, _37174_, _03703_);
  or (_37176_, _37038_, _03704_);
  and (_37177_, _37176_, _03385_);
  and (_37178_, _37177_, _37175_);
  and (_37180_, _37034_, _03384_);
  or (_37181_, _37180_, _03701_);
  or (_37182_, _37181_, _37178_);
  nor (_37183_, _13399_, _11659_);
  or (_37184_, _37023_, _03702_);
  or (_37185_, _37184_, _37183_);
  and (_37186_, _37185_, _42908_);
  and (_37187_, _37186_, _37182_);
  or (_37188_, _37187_, _37015_);
  and (_43337_, _37188_, _41654_);
  and (_37190_, _42912_, \oc8051_golden_model_1.P0INREG [0]);
  or (_37191_, _37190_, _01248_);
  and (_43340_, _37191_, _41654_);
  and (_37192_, _42912_, \oc8051_golden_model_1.P0INREG [1]);
  or (_37193_, _37192_, _01270_);
  and (_43341_, _37193_, _41654_);
  and (_37194_, _42912_, \oc8051_golden_model_1.P0INREG [2]);
  or (_37195_, _37194_, _01263_);
  and (_43342_, _37195_, _41654_);
  and (_37196_, _42912_, \oc8051_golden_model_1.P0INREG [3]);
  or (_37198_, _37196_, _01256_);
  and (_43343_, _37198_, _41654_);
  and (_37199_, _42912_, \oc8051_golden_model_1.P0INREG [4]);
  or (_37200_, _37199_, _01281_);
  and (_43344_, _37200_, _41654_);
  and (_37201_, _42912_, \oc8051_golden_model_1.P0INREG [5]);
  or (_37202_, _37201_, _01303_);
  and (_43347_, _37202_, _41654_);
  and (_37203_, _42912_, \oc8051_golden_model_1.P0INREG [6]);
  or (_37204_, _37203_, _01296_);
  and (_43348_, _37204_, _41654_);
  and (_37206_, _42912_, \oc8051_golden_model_1.P1INREG [0]);
  or (_37207_, _37206_, _01355_);
  and (_43349_, _37207_, _41654_);
  and (_37208_, _42912_, \oc8051_golden_model_1.P1INREG [1]);
  or (_37209_, _37208_, _01348_);
  and (_43351_, _37209_, _41654_);
  and (_37210_, _42912_, \oc8051_golden_model_1.P1INREG [2]);
  or (_37211_, _37210_, _01333_);
  and (_43352_, _37211_, _41654_);
  and (_37213_, _42912_, \oc8051_golden_model_1.P1INREG [3]);
  or (_37214_, _37213_, _01341_);
  and (_43353_, _37214_, _41654_);
  and (_37215_, _42912_, \oc8051_golden_model_1.P1INREG [4]);
  or (_37216_, _37215_, _01400_);
  and (_43354_, _37216_, _41654_);
  and (_37217_, _42912_, \oc8051_golden_model_1.P1INREG [5]);
  or (_37218_, _37217_, _01390_);
  and (_43355_, _37218_, _41654_);
  and (_37219_, _42912_, \oc8051_golden_model_1.P1INREG [6]);
  or (_37221_, _37219_, _01369_);
  and (_43356_, _37221_, _41654_);
  and (_37222_, _42912_, \oc8051_golden_model_1.P2INREG [0]);
  or (_37223_, _37222_, _01167_);
  and (_43359_, _37223_, _41654_);
  and (_37224_, _42912_, \oc8051_golden_model_1.P2INREG [1]);
  or (_37225_, _37224_, _01152_);
  and (_43360_, _37225_, _41654_);
  and (_37226_, _42912_, \oc8051_golden_model_1.P2INREG [2]);
  or (_37227_, _37226_, _01174_);
  and (_43361_, _37227_, _41654_);
  and (_37229_, _42912_, \oc8051_golden_model_1.P2INREG [3]);
  or (_37230_, _37229_, _01160_);
  and (_43362_, _37230_, _41654_);
  and (_37231_, _42912_, \oc8051_golden_model_1.P2INREG [4]);
  or (_37232_, _37231_, _01132_);
  and (_43363_, _37232_, _41654_);
  and (_37233_, _42912_, \oc8051_golden_model_1.P2INREG [5]);
  or (_37234_, _37233_, _01117_);
  and (_43364_, _37234_, _41654_);
  and (_37236_, _42912_, \oc8051_golden_model_1.P2INREG [6]);
  or (_37237_, _37236_, _01139_);
  and (_43365_, _37237_, _41654_);
  and (_37238_, _42912_, \oc8051_golden_model_1.P3INREG [0]);
  or (_37239_, _37238_, _01105_);
  and (_43367_, _37239_, _41654_);
  and (_37240_, _42912_, \oc8051_golden_model_1.P3INREG [1]);
  or (_37241_, _37240_, _01098_);
  and (_43368_, _37241_, _41654_);
  and (_37242_, _42912_, \oc8051_golden_model_1.P3INREG [2]);
  or (_37244_, _37242_, _01083_);
  and (_43369_, _37244_, _41654_);
  and (_37245_, _42912_, \oc8051_golden_model_1.P3INREG [3]);
  or (_37246_, _37245_, _01091_);
  and (_43370_, _37246_, _41654_);
  and (_37247_, _42912_, \oc8051_golden_model_1.P3INREG [4]);
  or (_37248_, _37247_, _01069_);
  and (_43371_, _37248_, _41654_);
  and (_37249_, _42912_, \oc8051_golden_model_1.P3INREG [5]);
  or (_37250_, _37249_, _01062_);
  and (_43372_, _37250_, _41654_);
  and (_37252_, _42912_, \oc8051_golden_model_1.P3INREG [6]);
  or (_37253_, _37252_, _01046_);
  and (_43373_, _37253_, _41654_);
  and (_00005_[6], _01047_, _41654_);
  and (_00005_[5], _01063_, _41654_);
  and (_00005_[4], _01070_, _41654_);
  and (_00005_[3], _01092_, _41654_);
  and (_00005_[2], _01084_, _41654_);
  and (_00005_[1], _01099_, _41654_);
  and (_00005_[0], _01106_, _41654_);
  and (_00004_[6], _01140_, _41654_);
  and (_00004_[5], _01118_, _41654_);
  and (_00004_[4], _01133_, _41654_);
  and (_00004_[3], _01161_, _41654_);
  and (_00004_[2], _01175_, _41654_);
  and (_00004_[1], _01153_, _41654_);
  and (_00004_[0], _01168_, _41654_);
  and (_00003_[6], _01371_, _41654_);
  and (_00003_[5], _01392_, _41654_);
  and (_00003_[4], _01401_, _41654_);
  and (_00003_[3], _01342_, _41654_);
  and (_00003_[2], _01334_, _41654_);
  and (_00003_[1], _01349_, _41654_);
  and (_00003_[0], _01356_, _41654_);
  and (_00002_[6], _01297_, _41654_);
  and (_00002_[5], _01304_, _41654_);
  and (_00002_[4], _01282_, _41654_);
  and (_00002_[3], _01257_, _41654_);
  and (_00002_[2], _01264_, _41654_);
  and (_00002_[1], _01271_, _41654_);
  and (_00002_[0], _01249_, _41654_);
  not (_37257_, _20509_);
  and (_37258_, _20596_, _37257_);
  not (_37259_, _21102_);
  and (_37260_, _21186_, _37259_);
  and (_37261_, _37260_, _37258_);
  not (_37262_, _18525_);
  and (_37263_, _18612_, _37262_);
  not (_37264_, _19904_);
  and (_37266_, _19991_, _37264_);
  and (_37267_, _37266_, _37263_);
  and (_37268_, _37267_, _37261_);
  not (_37269_, _21702_);
  and (_37270_, _21789_, _37269_);
  not (_37271_, _22305_);
  and (_37272_, _22393_, _37271_);
  nand (_37273_, _37272_, _37270_);
  nor (_37274_, _37273_, _17405_);
  and (_37275_, _37274_, _37268_);
  nor (_37277_, _20682_, _20081_);
  nor (_37278_, _22481_, _21272_);
  and (_37279_, _37278_, _37277_);
  or (_37280_, _03440_, _03383_);
  nor (_37281_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_37282_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and (_37283_, _37282_, _37281_);
  nor (_37284_, \oc8051_golden_model_1.IP [5], \oc8051_golden_model_1.IP [4]);
  nor (_37285_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [3]);
  and (_37286_, _37285_, _37284_);
  and (_37288_, _37286_, _37283_);
  nor (_37289_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor (_37290_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and (_37291_, _37290_, _37289_);
  nor (_37292_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor (_37293_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and (_37294_, _37293_, _37292_);
  and (_37295_, _37294_, _37291_);
  and (_37296_, _37295_, _37288_);
  nor (_37297_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor (_37299_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor (_37300_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and (_37301_, _37300_, _37299_);
  and (_37302_, _37301_, _37297_);
  nor (_37303_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_37304_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and (_37305_, _37304_, _37303_);
  nor (_37306_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor (_37307_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and (_37308_, _37307_, _37306_);
  and (_37310_, _37308_, _37305_);
  and (_37311_, _37310_, _37302_);
  and (_37312_, _37311_, _37296_);
  nor (_37313_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor (_37314_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and (_37315_, _37314_, _37313_);
  nor (_37316_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_37317_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and (_37318_, _37317_, _37316_);
  and (_37319_, _37318_, _37315_);
  nor (_37321_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  nor (_37322_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  and (_37323_, _37322_, _37321_);
  nor (_37324_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor (_37325_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and (_37326_, _37325_, _37324_);
  and (_37327_, _37326_, _37323_);
  and (_37328_, _37327_, _37319_);
  nor (_37329_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_37330_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and (_37332_, _37330_, _37329_);
  nor (_37333_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  nor (_37334_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  and (_37335_, _37334_, _37333_);
  and (_37336_, _37335_, _37332_);
  nor (_37337_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor (_37338_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and (_37339_, _37338_, _37337_);
  nor (_37340_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor (_37341_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and (_37343_, _37341_, _37340_);
  and (_37344_, _37343_, _37339_);
  and (_37345_, _37344_, _37336_);
  and (_37346_, _37345_, _37328_);
  nor (_37347_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and (_37348_, _37347_, op0_cnst);
  nor (_37349_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor (_37350_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and (_37351_, _37350_, _37349_);
  nor (_37352_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor (_37354_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and (_37355_, _37354_, _37352_);
  and (_37356_, _37355_, _37351_);
  and (_37357_, _37356_, _37348_);
  nor (_37358_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_37359_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and (_37360_, _37359_, _37358_);
  nor (_37361_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor (_37362_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and (_37363_, _37362_, _37361_);
  and (_37365_, _37363_, _37360_);
  and (_37366_, \oc8051_golden_model_1.TCON [1], _19051_);
  nor (_37367_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and (_37368_, _37367_, _37366_);
  nor (_37369_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor (_37370_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and (_37371_, _37370_, _37369_);
  and (_37372_, _37371_, _37368_);
  and (_37373_, _37372_, _37365_);
  and (_37374_, _37373_, _37357_);
  and (_37376_, _37374_, _37346_);
  and (_37377_, _37376_, _37312_);
  and (_37378_, _37377_, _03188_);
  nand (_37379_, _37378_, _37280_);
  nor (_37380_, _37379_, _17145_);
  nor (_37381_, _18700_, _17318_);
  and (_37382_, _37381_, _37380_);
  and (_37383_, _37382_, _37279_);
  and (_37384_, _37383_, _37275_);
  or (_37385_, _22134_, _21531_);
  or (_37387_, _37385_, _22740_);
  nor (_37388_, _37387_, _17885_);
  and (_37389_, _37388_, _37384_);
  not (_37390_, _18873_);
  and (_37391_, _37390_, _17774_);
  not (_37392_, _19047_);
  and (_37393_, _19155_, _37392_);
  and (_37394_, _37393_, _37391_);
  and (_37395_, _09509_, _09428_);
  and (_37396_, _37395_, _09590_);
  and (_37398_, _09086_, _08895_);
  and (_37399_, _09348_, _09268_);
  and (_37400_, _37399_, _37398_);
  and (_37401_, _37400_, _37396_);
  nor (_37402_, _17665_, _17493_);
  and (_37403_, _37402_, _37401_);
  and (_37404_, _37403_, _37394_);
  and (_37405_, _37404_, _37389_);
  not (_37406_, _23048_);
  nand (_37407_, _37406_, _19266_);
  or (_37409_, _37407_, _23822_);
  nor (_37410_, _37409_, _09006_);
  and (_37411_, _37410_, _37405_);
  or (_37412_, _23164_, _19381_);
  nor (_37413_, _37412_, _23934_);
  nor (_37414_, _21617_, _21444_);
  nor (_37415_, _22224_, _22047_);
  and (_37416_, _37415_, _37414_);
  nor (_37417_, _20426_, _20253_);
  nor (_37418_, _21023_, _20854_);
  and (_37420_, _37418_, _37417_);
  and (_37421_, _37420_, _37416_);
  nor (_37422_, _22828_, _22653_);
  and (_37423_, _23712_, _22936_);
  nand (_37424_, _37423_, _37422_);
  nor (_37425_, _37424_, _18001_);
  and (_37426_, _37425_, _37421_);
  and (_37427_, _37426_, _37413_);
  and (_37428_, _37427_, _37411_);
  or (_00001_, _37428_, rst);
  and (_00005_[7], _01056_, _41654_);
  and (_00004_[7], _01126_, _41654_);
  and (_00003_[7], _01382_, _41654_);
  and (_00002_[7], _01290_, _41654_);
  and (_37430_, _37428_, inst_finished_r);
  not (_37431_, word_in[1]);
  and (_37432_, _37431_, word_in[0]);
  and (_37433_, _37432_, \oc8051_golden_model_1.IRAM[5] [0]);
  nor (_37434_, _37431_, word_in[0]);
  and (_37435_, _37434_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_37437_, _37435_, _37433_);
  nor (_37438_, word_in[1], word_in[0]);
  and (_37439_, _37438_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_37440_, word_in[1], word_in[0]);
  and (_37441_, _37440_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_37442_, _37441_, _37439_);
  and (_37443_, _37442_, _37437_);
  not (_37444_, word_in[3]);
  and (_37445_, _37444_, word_in[2]);
  not (_37446_, _37445_);
  nor (_37448_, _37446_, _37443_);
  and (_37449_, _37432_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_37450_, _37434_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor (_37451_, _37450_, _37449_);
  and (_37452_, _37438_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_37453_, _37440_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor (_37454_, _37453_, _37452_);
  and (_37455_, _37454_, _37451_);
  nor (_37456_, _37444_, word_in[2]);
  not (_37457_, _37456_);
  nor (_37459_, _37457_, _37455_);
  nor (_37460_, _37459_, _37448_);
  and (_37461_, _37432_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_37462_, _37434_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor (_37463_, _37462_, _37461_);
  and (_37464_, _37438_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_37465_, _37440_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor (_37466_, _37465_, _37464_);
  and (_37467_, _37466_, _37463_);
  nor (_37468_, word_in[3], word_in[2]);
  not (_37470_, _37468_);
  nor (_37471_, _37470_, _37467_);
  and (_37472_, _37432_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_37473_, _37434_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor (_37474_, _37473_, _37472_);
  and (_37475_, _37438_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_37476_, _37440_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor (_37477_, _37476_, _37475_);
  and (_37478_, _37477_, _37474_);
  and (_37479_, word_in[3], word_in[2]);
  not (_37481_, _37479_);
  nor (_37482_, _37481_, _37478_);
  nor (_37483_, _37482_, _37471_);
  and (_37484_, _37483_, _37460_);
  and (_37485_, _37456_, _37432_);
  and (_37486_, _37485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_37487_, _37468_, _37434_);
  and (_37488_, _37487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_37489_, _37488_, _37486_);
  and (_37490_, _37479_, _37434_);
  and (_37492_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_37493_, _37445_, _37432_);
  and (_37494_, _37493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_37495_, _37494_, _37492_);
  and (_37496_, _37495_, _37489_);
  and (_37497_, _37456_, _37440_);
  and (_37498_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_37499_, _37456_, _37438_);
  and (_37500_, _37499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_37501_, _37500_, _37498_);
  and (_37503_, _37479_, _37438_);
  and (_37504_, _37503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_37505_, _37468_, _37440_);
  and (_37506_, _37505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_37507_, _37506_, _37504_);
  and (_37508_, _37507_, _37501_);
  and (_37509_, _37508_, _37496_);
  and (_37510_, _37445_, _37440_);
  and (_37511_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_37512_, _37445_, _37434_);
  and (_37514_, _37512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_37515_, _37514_, _37511_);
  and (_37516_, _37445_, _37438_);
  and (_37517_, _37516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_37518_, _37468_, _37438_);
  and (_37519_, _37518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_37520_, _37519_, _37517_);
  and (_37521_, _37520_, _37515_);
  and (_37522_, _37456_, _37434_);
  and (_37523_, _37522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_37525_, _37468_, _37432_);
  and (_37526_, _37525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_37527_, _37526_, _37523_);
  and (_37528_, _37479_, _37440_);
  and (_37529_, _37528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_37530_, _37479_, _37432_);
  and (_37531_, _37530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_37532_, _37531_, _37529_);
  and (_37533_, _37532_, _37527_);
  and (_37534_, _37533_, _37521_);
  and (_37536_, _37534_, _37509_);
  nand (_37537_, _37536_, _37484_);
  or (_37538_, _37536_, _37484_);
  and (_37539_, _37538_, _37537_);
  and (_37540_, _37432_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_37541_, _37434_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor (_37542_, _37541_, _37540_);
  and (_37543_, _37438_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_37544_, _37440_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_37545_, _37544_, _37543_);
  and (_37547_, _37545_, _37542_);
  nor (_37548_, _37547_, _37446_);
  and (_37549_, _37432_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_37550_, _37434_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor (_37551_, _37550_, _37549_);
  and (_37552_, _37438_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_37553_, _37440_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor (_37554_, _37553_, _37552_);
  and (_37555_, _37554_, _37551_);
  nor (_37556_, _37555_, _37481_);
  nor (_37558_, _37556_, _37548_);
  and (_37559_, _37432_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_37560_, _37434_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor (_37561_, _37560_, _37559_);
  and (_37562_, _37438_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_37563_, _37440_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor (_37564_, _37563_, _37562_);
  and (_37565_, _37564_, _37561_);
  nor (_37566_, _37565_, _37470_);
  and (_37567_, _37432_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_37569_, _37434_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor (_37570_, _37569_, _37567_);
  and (_37571_, _37438_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_37572_, _37440_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor (_37573_, _37572_, _37571_);
  and (_37574_, _37573_, _37570_);
  nor (_37575_, _37574_, _37457_);
  nor (_37576_, _37575_, _37566_);
  and (_37577_, _37576_, _37558_);
  and (_37578_, _37528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_37580_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_37581_, _37580_, _37578_);
  and (_37582_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37583_, _37518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_37584_, _37583_, _37582_);
  and (_37585_, _37584_, _37581_);
  and (_37586_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_37587_, _37530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_37588_, _37587_, _37586_);
  and (_37589_, _37522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_37591_, _37485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_37592_, _37591_, _37589_);
  and (_37593_, _37592_, _37588_);
  and (_37594_, _37593_, _37585_);
  and (_37595_, _37516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_37596_, _37505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_37597_, _37596_, _37595_);
  and (_37598_, _37512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_37599_, _37493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_37600_, _37599_, _37598_);
  and (_37602_, _37600_, _37597_);
  and (_37603_, _37487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_37604_, _37525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_37605_, _37604_, _37603_);
  and (_37606_, _37503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_37607_, _37499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_37608_, _37607_, _37606_);
  and (_37609_, _37608_, _37605_);
  and (_37610_, _37609_, _37602_);
  and (_37611_, _37610_, _37594_);
  nand (_37613_, _37611_, _37577_);
  or (_37614_, _37611_, _37577_);
  and (_37615_, _37614_, _37613_);
  or (_37616_, _37615_, _37539_);
  and (_37617_, _37432_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_37618_, _37434_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor (_37619_, _37618_, _37617_);
  and (_37620_, _37438_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_37621_, _37440_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor (_37622_, _37621_, _37620_);
  and (_37624_, _37622_, _37619_);
  nor (_37625_, _37624_, _37470_);
  and (_37626_, _37432_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_37627_, _37434_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor (_37628_, _37627_, _37626_);
  and (_37629_, _37438_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_37630_, _37440_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor (_37631_, _37630_, _37629_);
  and (_37632_, _37631_, _37628_);
  nor (_37633_, _37632_, _37481_);
  nor (_37635_, _37633_, _37625_);
  and (_37636_, _37432_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_37637_, _37434_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_37638_, _37637_, _37636_);
  and (_37639_, _37438_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_37640_, _37440_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor (_37641_, _37640_, _37639_);
  and (_37642_, _37641_, _37638_);
  nor (_37643_, _37642_, _37446_);
  and (_37644_, _37432_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_37646_, _37434_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor (_37647_, _37646_, _37644_);
  and (_37648_, _37438_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_37649_, _37440_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor (_37650_, _37649_, _37648_);
  and (_37651_, _37650_, _37647_);
  nor (_37652_, _37651_, _37457_);
  nor (_37653_, _37652_, _37643_);
  and (_37654_, _37653_, _37635_);
  and (_37655_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_37657_, _37505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_37658_, _37657_, _37655_);
  and (_37659_, _37530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_37660_, _37503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_37661_, _37660_, _37659_);
  and (_37662_, _37661_, _37658_);
  and (_37663_, _37512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_37664_, _37493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_37665_, _37664_, _37663_);
  and (_37666_, _37516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_37668_, _37518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_37669_, _37668_, _37666_);
  and (_37670_, _37669_, _37665_);
  and (_37671_, _37670_, _37662_);
  and (_37672_, _37528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_37673_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_37674_, _37673_, _37672_);
  and (_37675_, _37522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_37676_, _37499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_37677_, _37676_, _37675_);
  and (_37679_, _37677_, _37674_);
  and (_37680_, _37487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_37681_, _37525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_37682_, _37681_, _37680_);
  and (_37683_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_37684_, _37485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_37685_, _37684_, _37683_);
  and (_37686_, _37685_, _37682_);
  and (_37687_, _37686_, _37679_);
  and (_37688_, _37687_, _37671_);
  nand (_37690_, _37688_, _37654_);
  or (_37691_, _37688_, _37654_);
  and (_37692_, _37691_, _37690_);
  and (_37693_, _37432_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_37694_, _37434_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor (_37695_, _37694_, _37693_);
  and (_37696_, _37438_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_37697_, _37440_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor (_37698_, _37697_, _37696_);
  and (_37699_, _37698_, _37695_);
  nor (_37701_, _37699_, _37446_);
  and (_37702_, _37432_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_37703_, _37434_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor (_37704_, _37703_, _37702_);
  and (_37705_, _37438_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_37706_, _37440_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor (_37707_, _37706_, _37705_);
  and (_37708_, _37707_, _37704_);
  nor (_37709_, _37708_, _37457_);
  nor (_37710_, _37709_, _37701_);
  and (_37712_, _37432_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_37713_, _37434_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor (_37714_, _37713_, _37712_);
  and (_37715_, _37438_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_37716_, _37440_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor (_37717_, _37716_, _37715_);
  and (_37718_, _37717_, _37714_);
  nor (_37719_, _37718_, _37470_);
  and (_37720_, _37432_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_37721_, _37434_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor (_37723_, _37721_, _37720_);
  and (_37724_, _37438_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_37725_, _37440_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor (_37726_, _37725_, _37724_);
  and (_37727_, _37726_, _37723_);
  nor (_37728_, _37727_, _37481_);
  nor (_37729_, _37728_, _37719_);
  and (_37730_, _37729_, _37710_);
  not (_37731_, _37730_);
  and (_37732_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_37734_, _37522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_37735_, _37734_, _37732_);
  and (_37736_, _37530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_37737_, _37485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_37738_, _37737_, _37736_);
  and (_37739_, _37738_, _37735_);
  and (_37740_, _37516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_37741_, _37487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_37742_, _37741_, _37740_);
  and (_37743_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_37745_, _37493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_37746_, _37745_, _37743_);
  and (_37747_, _37746_, _37742_);
  and (_37748_, _37747_, _37739_);
  and (_37749_, _37503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_37750_, _37525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_37751_, _37750_, _37749_);
  and (_37752_, _37499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_37753_, _37505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_37754_, _37753_, _37752_);
  and (_37756_, _37754_, _37751_);
  and (_37757_, _37528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_37758_, _37518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_37759_, _37758_, _37757_);
  and (_37760_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_37761_, _37512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_37762_, _37761_, _37760_);
  and (_37763_, _37762_, _37759_);
  and (_37764_, _37763_, _37756_);
  and (_37765_, _37764_, _37748_);
  nor (_37767_, _37765_, _37731_);
  and (_37768_, _37765_, _37731_);
  or (_37769_, _37768_, _37767_);
  or (_37770_, _37769_, _37692_);
  or (_37771_, _37770_, _37616_);
  and (_37772_, _37432_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_37773_, _37434_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor (_37774_, _37773_, _37772_);
  and (_37775_, _37438_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_37776_, _37440_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor (_37778_, _37776_, _37775_);
  and (_37779_, _37778_, _37774_);
  nor (_37780_, _37779_, _37446_);
  and (_37781_, _37432_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_37782_, _37434_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor (_37783_, _37782_, _37781_);
  and (_37784_, _37438_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_37785_, _37440_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor (_37786_, _37785_, _37784_);
  and (_37787_, _37786_, _37783_);
  nor (_37789_, _37787_, _37481_);
  nor (_37790_, _37789_, _37780_);
  and (_37791_, _37432_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_37792_, _37434_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor (_37793_, _37792_, _37791_);
  and (_37794_, _37438_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_37795_, _37440_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor (_37796_, _37795_, _37794_);
  and (_37797_, _37796_, _37793_);
  nor (_37798_, _37797_, _37470_);
  and (_37800_, _37432_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_37801_, _37434_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor (_37802_, _37801_, _37800_);
  and (_37803_, _37438_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_37804_, _37440_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor (_37805_, _37804_, _37803_);
  and (_37806_, _37805_, _37802_);
  nor (_37807_, _37806_, _37457_);
  nor (_37808_, _37807_, _37798_);
  and (_37809_, _37808_, _37790_);
  and (_37811_, _37503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_37812_, _37525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_37813_, _37812_, _37811_);
  and (_37814_, _37530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_37815_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_37816_, _37815_, _37814_);
  and (_37817_, _37816_, _37813_);
  and (_37818_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_37819_, _37522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_37820_, _37819_, _37818_);
  and (_37822_, _37505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_37823_, _37518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_37824_, _37823_, _37822_);
  and (_37825_, _37824_, _37820_);
  and (_37826_, _37825_, _37817_);
  and (_37827_, _37499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_37828_, _37493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_37829_, _37828_, _37827_);
  and (_37830_, _37528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_37831_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_37833_, _37831_, _37830_);
  and (_37834_, _37833_, _37829_);
  and (_37835_, _37485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_37836_, _37512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_37837_, _37836_, _37835_);
  and (_37838_, _37516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_37839_, _37487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_37840_, _37839_, _37838_);
  and (_37841_, _37840_, _37837_);
  and (_37842_, _37841_, _37834_);
  and (_37844_, _37842_, _37826_);
  or (_37845_, _37844_, _37809_);
  nand (_37846_, _37844_, _37809_);
  and (_37847_, _37846_, _37845_);
  and (_37848_, _37432_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_37849_, _37434_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor (_37850_, _37849_, _37848_);
  and (_37851_, _37438_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_37852_, _37440_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor (_37853_, _37852_, _37851_);
  and (_37855_, _37853_, _37850_);
  nor (_37856_, _37855_, _37446_);
  and (_37857_, _37432_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_37858_, _37434_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor (_37859_, _37858_, _37857_);
  and (_37860_, _37438_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_37861_, _37440_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor (_37862_, _37861_, _37860_);
  and (_37863_, _37862_, _37859_);
  nor (_37864_, _37863_, _37481_);
  nor (_37866_, _37864_, _37856_);
  and (_37867_, _37432_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_37868_, _37434_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor (_37869_, _37868_, _37867_);
  and (_37870_, _37438_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_37871_, _37440_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor (_37872_, _37871_, _37870_);
  and (_37873_, _37872_, _37869_);
  nor (_37874_, _37873_, _37470_);
  and (_37875_, _37432_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_37877_, _37434_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor (_37878_, _37877_, _37875_);
  and (_37879_, _37438_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_37880_, _37440_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor (_37881_, _37880_, _37879_);
  and (_37882_, _37881_, _37878_);
  nor (_37883_, _37882_, _37457_);
  nor (_37884_, _37883_, _37874_);
  and (_37885_, _37884_, _37866_);
  and (_37886_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_37888_, _37522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_37889_, _37888_, _37886_);
  and (_37890_, _37530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_37891_, _37485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_37892_, _37891_, _37890_);
  and (_37893_, _37892_, _37889_);
  and (_37894_, _37493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_37895_, _37487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_37896_, _37895_, _37894_);
  and (_37897_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_37899_, _37516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_37900_, _37899_, _37897_);
  and (_37901_, _37900_, _37896_);
  and (_37902_, _37901_, _37893_);
  and (_37903_, _37503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_37904_, _37525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_37905_, _37904_, _37903_);
  and (_37906_, _37499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_37907_, _37505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_37908_, _37907_, _37906_);
  and (_37910_, _37908_, _37905_);
  and (_37911_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_37912_, _37518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_37913_, _37912_, _37911_);
  and (_37914_, _37528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_37915_, _37512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_37916_, _37915_, _37914_);
  and (_37917_, _37916_, _37913_);
  and (_37918_, _37917_, _37910_);
  and (_37919_, _37918_, _37902_);
  or (_37921_, _37919_, _37885_);
  nand (_37922_, _37919_, _37885_);
  and (_37923_, _37922_, _37921_);
  or (_37924_, _37923_, _37847_);
  and (_37925_, _37432_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_37926_, _37434_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor (_37927_, _37926_, _37925_);
  and (_37928_, _37438_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_37929_, _37440_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor (_37930_, _37929_, _37928_);
  and (_37932_, _37930_, _37927_);
  nor (_37933_, _37932_, _37446_);
  and (_37934_, _37432_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_37935_, _37434_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_37936_, _37935_, _37934_);
  and (_37937_, _37438_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_37938_, _37440_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor (_37939_, _37938_, _37937_);
  and (_37940_, _37939_, _37936_);
  nor (_37941_, _37940_, _37481_);
  nor (_37943_, _37941_, _37933_);
  and (_37944_, _37432_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_37945_, _37434_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor (_37946_, _37945_, _37944_);
  and (_37947_, _37438_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_37948_, _37440_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor (_37949_, _37948_, _37947_);
  and (_37950_, _37949_, _37946_);
  nor (_37951_, _37950_, _37470_);
  and (_37952_, _37432_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_37954_, _37434_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor (_37955_, _37954_, _37952_);
  and (_37956_, _37438_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_37957_, _37440_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_37958_, _37957_, _37956_);
  and (_37959_, _37958_, _37955_);
  nor (_37960_, _37959_, _37457_);
  nor (_37961_, _37960_, _37951_);
  and (_37962_, _37961_, _37943_);
  and (_37963_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_37965_, _37522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor (_37966_, _37965_, _37963_);
  and (_37967_, _37530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_37968_, _37485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_37969_, _37968_, _37967_);
  and (_37970_, _37969_, _37966_);
  and (_37971_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_37972_, _37512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_37973_, _37972_, _37971_);
  and (_37974_, _37493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_37976_, _37487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_37977_, _37976_, _37974_);
  and (_37978_, _37977_, _37973_);
  and (_37979_, _37978_, _37970_);
  and (_37980_, _37503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_37981_, _37518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_37982_, _37981_, _37980_);
  and (_37983_, _37499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_37984_, _37505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_37985_, _37984_, _37983_);
  and (_37987_, _37985_, _37982_);
  and (_37988_, _37528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_37989_, _37525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_37990_, _37989_, _37988_);
  and (_37991_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_37992_, _37516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_37993_, _37992_, _37991_);
  and (_37994_, _37993_, _37990_);
  and (_37995_, _37994_, _37987_);
  and (_37996_, _37995_, _37979_);
  nand (_37998_, _37996_, _37962_);
  or (_37999_, _37996_, _37962_);
  and (_38000_, _37999_, _37998_);
  and (_38001_, _37432_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_38002_, _37434_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor (_38003_, _38002_, _38001_);
  and (_38004_, _37438_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_38005_, _37440_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor (_38006_, _38005_, _38004_);
  and (_38007_, _38006_, _38003_);
  nor (_38009_, _38007_, _37470_);
  and (_38010_, _37432_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_38011_, _37434_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor (_38012_, _38011_, _38010_);
  and (_38013_, _37438_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_38014_, _37440_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor (_38015_, _38014_, _38013_);
  and (_38016_, _38015_, _38012_);
  nor (_38017_, _38016_, _37457_);
  nor (_38018_, _38017_, _38009_);
  and (_38020_, _37432_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_38021_, _37434_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor (_38022_, _38021_, _38020_);
  and (_38023_, _37438_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_38024_, _37440_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor (_38025_, _38024_, _38023_);
  and (_38026_, _38025_, _38022_);
  nor (_38027_, _38026_, _37446_);
  and (_38028_, _37432_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_38029_, _37434_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_38031_, _38029_, _38028_);
  and (_38032_, _37438_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_38033_, _37440_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_38034_, _38033_, _38032_);
  and (_38035_, _38034_, _38031_);
  nor (_38036_, _38035_, _37481_);
  nor (_38037_, _38036_, _38027_);
  and (_38038_, _38037_, _38018_);
  and (_38039_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_38040_, _37525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_38042_, _38040_, _38039_);
  and (_38043_, _37485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_38044_, _37487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_38045_, _38044_, _38043_);
  and (_38046_, _38045_, _38042_);
  and (_38047_, _37530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_38048_, _37503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_38049_, _38048_, _38047_);
  and (_38050_, _37493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_38051_, _37516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_38053_, _38051_, _38050_);
  and (_38054_, _38053_, _38049_);
  and (_38055_, _38054_, _38046_);
  and (_38056_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_38057_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_38058_, _38057_, _38056_);
  and (_38059_, _37505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_38060_, _37518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_38061_, _38060_, _38059_);
  and (_38062_, _38061_, _38058_);
  and (_38064_, _37528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_38065_, _37512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_38066_, _38065_, _38064_);
  and (_38067_, _37522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_38068_, _37499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_38069_, _38068_, _38067_);
  and (_38070_, _38069_, _38066_);
  and (_38071_, _38070_, _38062_);
  and (_38072_, _38071_, _38055_);
  not (_38073_, _38072_);
  nor (_38075_, _38073_, _38038_);
  and (_38076_, _38073_, _38038_);
  or (_38077_, _38076_, _38075_);
  or (_38078_, _38077_, _38000_);
  or (_38079_, _38078_, _37924_);
  or (_38080_, _38079_, _37771_);
  and (property_invalid_iram, _38080_, _37430_);
  nand (_38081_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38082_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38083_, _38082_, _38081_);
  and (_38085_, _07740_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_38086_, _07740_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_38087_, _38086_, _38085_);
  or (_38088_, _38087_, _38083_);
  nor (_38089_, _03491_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38090_, _03491_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_38091_, _38090_, _38089_);
  and (_38092_, _03558_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38093_, _03558_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_38094_, _38093_, _38092_);
  or (_38096_, _38094_, _38091_);
  or (_38097_, _38096_, _38088_);
  or (_38098_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38099_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38100_, _38099_, _38098_);
  or (_38101_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_38102_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38103_, _38102_, _38101_);
  or (_38104_, _38103_, _38100_);
  and (_38105_, _07586_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_38107_, _07586_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_38108_, _38107_, _38105_);
  nand (_38109_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38110_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_38111_, _38110_, _38109_);
  or (_38112_, _38111_, _38108_);
  or (_38113_, _38112_, _38104_);
  or (_38114_, _38113_, _38097_);
  and (property_invalid_acc, _38114_, _37430_);
  nor (_38115_, _26334_, _43823_);
  and (_38117_, _26334_, _43823_);
  and (_38118_, _28111_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_38119_, _28111_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_38120_, _27403_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_38121_, _27403_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_38122_, _38121_, _38120_);
  nor (_38123_, _27761_, _43838_);
  and (_38124_, _27761_, _43838_);
  nor (_38125_, _27053_, _43831_);
  and (_38126_, _27053_, _43831_);
  nor (_38128_, _29114_, _38413_);
  and (_38129_, _29114_, _38413_);
  or (_38130_, _30049_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_38131_, _30049_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38132_, _38131_, _38130_);
  nand (_38133_, _29430_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_38134_, _29430_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38135_, _38134_, _38133_);
  or (_38136_, _30669_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_38137_, _30669_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38139_, _38137_, _38136_);
  nor (_38140_, _10935_, _38435_);
  and (_38141_, _10935_, _38435_);
  or (_38142_, _38141_, _38140_);
  nor (_38143_, _29735_, _38403_);
  and (_38144_, _29735_, _38403_);
  or (_38145_, _38144_, _38143_);
  or (_38146_, _25933_, _43819_);
  nand (_38147_, _25933_, _43819_);
  and (_38148_, _38147_, _38146_);
  or (_38150_, _38148_, _38145_);
  or (_38151_, _38150_, _38142_);
  or (_38152_, _38151_, _38139_);
  and (_38153_, _30354_, _38399_);
  nor (_38154_, _30354_, _38399_);
  or (_38155_, _38154_, _38153_);
  or (_38156_, _38155_, _38152_);
  and (_38157_, _28785_, _38407_);
  nor (_38158_, _28785_, _38407_);
  or (_38159_, _38158_, _38157_);
  or (_38161_, _38159_, _38156_);
  or (_38162_, _38161_, _38135_);
  or (_38163_, _38162_, _38132_);
  or (_38164_, _38163_, _38129_);
  or (_38165_, _38164_, _38128_);
  or (_38166_, _38165_, _38126_);
  or (_38167_, _38166_, _38125_);
  or (_38168_, _38167_, _38124_);
  or (_38169_, _38168_, _38123_);
  or (_38170_, _38169_, _38122_);
  or (_38172_, _38170_, _38119_);
  or (_38173_, _38172_, _38118_);
  nor (_38174_, _28464_, _43845_);
  and (_38175_, _28464_, _43845_);
  or (_38176_, _38175_, _38174_);
  or (_38177_, _38176_, _38173_);
  and (_38178_, _26703_, _43827_);
  nor (_38179_, _26703_, _43827_);
  or (_38180_, _38179_, _38178_);
  or (_38181_, _38180_, _38177_);
  or (_38183_, _38181_, _38117_);
  or (_38184_, _38183_, _38115_);
  and (_38185_, _37428_, _42908_);
  and (property_invalid_pc, _38185_, _38184_);
  buf (_01387_, _41654_);
  buf (_01440_, _41654_);
  buf (_01493_, _41654_);
  buf (_01545_, _41654_);
  buf (_01597_, _41654_);
  buf (_01649_, _41654_);
  buf (_01701_, _41654_);
  buf (_01752_, _41654_);
  buf (_01804_, _41654_);
  buf (_01855_, _41654_);
  buf (_01894_, _41654_);
  buf (_01947_, _41654_);
  buf (_02000_, _41654_);
  buf (_02051_, _41654_);
  buf (_02103_, _41654_);
  buf (_02155_, _41654_);
  buf (_38725_, _38627_);
  buf (_38726_, _38628_);
  buf (_38738_, _38627_);
  buf (_38739_, _38628_);
  buf (_39052_, _38646_);
  buf (_39053_, _38648_);
  buf (_39054_, _38649_);
  buf (_39055_, _38650_);
  buf (_39056_, _38651_);
  buf (_39057_, _38652_);
  buf (_39058_, _38654_);
  buf (_39060_, _38655_);
  buf (_39061_, _38656_);
  buf (_39062_, _38657_);
  buf (_39063_, _38658_);
  buf (_39064_, _38660_);
  buf (_39065_, _38661_);
  buf (_39066_, _38662_);
  buf (_39118_, _38646_);
  buf (_39119_, _38648_);
  buf (_39120_, _38649_);
  buf (_39121_, _38650_);
  buf (_39122_, _38651_);
  buf (_39123_, _38652_);
  buf (_39124_, _38654_);
  buf (_39126_, _38655_);
  buf (_39127_, _38656_);
  buf (_39128_, _38657_);
  buf (_39129_, _38658_);
  buf (_39130_, _38660_);
  buf (_39131_, _38661_);
  buf (_39132_, _38662_);
  buf (_39524_, _39429_);
  buf (_39639_, _39429_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _01391_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _01395_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _01399_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _01403_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _01407_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _01411_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _01415_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _01384_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _01387_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _01444_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _01448_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _01452_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _01456_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _01460_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _01464_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _01468_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _01437_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _01440_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _01898_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _01902_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _01906_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _01910_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _01914_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _01918_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _01922_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _01892_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _01894_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _01951_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _01955_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _01959_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _01963_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _01967_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _01971_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _01975_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _01944_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _01947_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _02004_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _02007_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _02011_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _02015_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _02019_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _02023_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _02027_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _01997_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _02000_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _02055_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _02059_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _02063_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _02067_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _02071_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _02075_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _02079_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _02048_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _02051_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _02107_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _02111_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _02115_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _02118_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _02122_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _02126_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _02130_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _02100_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _02103_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _02159_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _02163_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _02167_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _02171_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _02174_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _02178_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _02182_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _02152_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _02155_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _01497_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _01501_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _01505_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _01509_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _01513_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _01517_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _01521_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _01490_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _01493_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _01549_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _01552_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _01556_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _01560_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _01564_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _01568_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _01572_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _01542_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _01545_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _01601_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _01605_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _01609_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _01613_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _01617_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _01621_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _01624_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _01594_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _01597_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _01653_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _01657_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _01661_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _01665_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _01668_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _01672_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _01676_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _01646_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _01649_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _01704_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _01708_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _01712_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _01716_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _01720_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _01724_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _01728_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _01698_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _01701_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _01756_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _01760_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _01764_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _01768_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _01772_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _01776_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _01780_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _01749_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _01752_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _01808_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _01812_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _01816_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _01819_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _01823_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _01827_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _01831_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _01801_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _01804_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _01859_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _01863_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _01867_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _01871_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _01875_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _01879_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _01883_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _01852_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _01855_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _40671_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _40672_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _40674_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _40675_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _40676_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _40677_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _40678_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40439_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _40659_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _40660_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _40662_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _40663_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _40664_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _40665_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _40666_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _40668_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _40647_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _40648_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _40650_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _40651_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _40652_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _40653_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _40654_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _40656_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40635_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40636_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40637_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40639_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40640_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40641_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40642_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40643_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40623_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40624_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40625_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40626_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40628_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40629_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40630_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40631_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40611_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40612_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40613_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40614_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40615_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40617_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40618_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40619_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40599_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40600_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40601_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40602_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40603_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40605_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40606_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40607_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40586_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40588_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40589_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40590_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40591_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40592_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40594_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40595_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40574_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40575_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40576_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40577_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40579_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40580_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40581_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40582_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40562_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40563_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40564_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40565_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40566_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40568_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40569_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40570_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40550_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40551_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40552_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40553_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40554_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40556_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40557_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40558_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40537_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40539_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40540_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40541_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40542_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40543_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40545_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40546_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40525_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40526_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40527_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40528_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40530_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40531_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40532_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40533_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40512_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40514_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40515_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40516_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40517_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40518_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40520_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40521_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40500_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40501_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40502_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40503_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40505_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40506_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40507_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40508_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40486_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40487_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40489_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40490_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40491_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40493_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40494_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40495_);
  dff (\oc8051_golden_model_1.B [0], _43136_);
  dff (\oc8051_golden_model_1.B [1], _43137_);
  dff (\oc8051_golden_model_1.B [2], _43138_);
  dff (\oc8051_golden_model_1.B [3], _43139_);
  dff (\oc8051_golden_model_1.B [4], _43140_);
  dff (\oc8051_golden_model_1.B [5], _43141_);
  dff (\oc8051_golden_model_1.B [6], _43142_);
  dff (\oc8051_golden_model_1.B [7], _40440_);
  dff (\oc8051_golden_model_1.ACC [0], _43143_);
  dff (\oc8051_golden_model_1.ACC [1], _43144_);
  dff (\oc8051_golden_model_1.ACC [2], _43145_);
  dff (\oc8051_golden_model_1.ACC [3], _43146_);
  dff (\oc8051_golden_model_1.ACC [4], _43147_);
  dff (\oc8051_golden_model_1.ACC [5], _43150_);
  dff (\oc8051_golden_model_1.ACC [6], _43151_);
  dff (\oc8051_golden_model_1.ACC [7], _40441_);
  dff (\oc8051_golden_model_1.SBUF [0], _43152_);
  dff (\oc8051_golden_model_1.SBUF [1], _43155_);
  dff (\oc8051_golden_model_1.SBUF [2], _43156_);
  dff (\oc8051_golden_model_1.SBUF [3], _43157_);
  dff (\oc8051_golden_model_1.SBUF [4], _43158_);
  dff (\oc8051_golden_model_1.SBUF [5], _43159_);
  dff (\oc8051_golden_model_1.SBUF [6], _43160_);
  dff (\oc8051_golden_model_1.SBUF [7], _40443_);
  dff (\oc8051_golden_model_1.SCON [0], _43161_);
  dff (\oc8051_golden_model_1.SCON [1], _43162_);
  dff (\oc8051_golden_model_1.SCON [2], _43163_);
  dff (\oc8051_golden_model_1.SCON [3], _43164_);
  dff (\oc8051_golden_model_1.SCON [4], _43165_);
  dff (\oc8051_golden_model_1.SCON [5], _43166_);
  dff (\oc8051_golden_model_1.SCON [6], _43167_);
  dff (\oc8051_golden_model_1.SCON [7], _40444_);
  dff (\oc8051_golden_model_1.PCON [0], _43170_);
  dff (\oc8051_golden_model_1.PCON [1], _43171_);
  dff (\oc8051_golden_model_1.PCON [2], _43172_);
  dff (\oc8051_golden_model_1.PCON [3], _43175_);
  dff (\oc8051_golden_model_1.PCON [4], _43176_);
  dff (\oc8051_golden_model_1.PCON [5], _43177_);
  dff (\oc8051_golden_model_1.PCON [6], _43178_);
  dff (\oc8051_golden_model_1.PCON [7], _40445_);
  dff (\oc8051_golden_model_1.TCON [0], _43179_);
  dff (\oc8051_golden_model_1.TCON [1], _43180_);
  dff (\oc8051_golden_model_1.TCON [2], _43181_);
  dff (\oc8051_golden_model_1.TCON [3], _43182_);
  dff (\oc8051_golden_model_1.TCON [4], _43183_);
  dff (\oc8051_golden_model_1.TCON [5], _43184_);
  dff (\oc8051_golden_model_1.TCON [6], _43185_);
  dff (\oc8051_golden_model_1.TCON [7], _40446_);
  dff (\oc8051_golden_model_1.TL0 [0], _43188_);
  dff (\oc8051_golden_model_1.TL0 [1], _43189_);
  dff (\oc8051_golden_model_1.TL0 [2], _43190_);
  dff (\oc8051_golden_model_1.TL0 [3], _43191_);
  dff (\oc8051_golden_model_1.TL0 [4], _43192_);
  dff (\oc8051_golden_model_1.TL0 [5], _43195_);
  dff (\oc8051_golden_model_1.TL0 [6], _43196_);
  dff (\oc8051_golden_model_1.TL0 [7], _40447_);
  dff (\oc8051_golden_model_1.TL1 [0], _43197_);
  dff (\oc8051_golden_model_1.TL1 [1], _43199_);
  dff (\oc8051_golden_model_1.TL1 [2], _43200_);
  dff (\oc8051_golden_model_1.TL1 [3], _43201_);
  dff (\oc8051_golden_model_1.TL1 [4], _43202_);
  dff (\oc8051_golden_model_1.TL1 [5], _43203_);
  dff (\oc8051_golden_model_1.TL1 [6], _43204_);
  dff (\oc8051_golden_model_1.TL1 [7], _40449_);
  dff (\oc8051_golden_model_1.TH0 [0], _43207_);
  dff (\oc8051_golden_model_1.TH0 [1], _43208_);
  dff (\oc8051_golden_model_1.TH0 [2], _43209_);
  dff (\oc8051_golden_model_1.TH0 [3], _43210_);
  dff (\oc8051_golden_model_1.TH0 [4], _43211_);
  dff (\oc8051_golden_model_1.TH0 [5], _43212_);
  dff (\oc8051_golden_model_1.TH0 [6], _43213_);
  dff (\oc8051_golden_model_1.TH0 [7], _40450_);
  dff (\oc8051_golden_model_1.TH1 [0], _43215_);
  dff (\oc8051_golden_model_1.TH1 [1], _43216_);
  dff (\oc8051_golden_model_1.TH1 [2], _43217_);
  dff (\oc8051_golden_model_1.TH1 [3], _43218_);
  dff (\oc8051_golden_model_1.TH1 [4], _43219_);
  dff (\oc8051_golden_model_1.TH1 [5], _43220_);
  dff (\oc8051_golden_model_1.TH1 [6], _43221_);
  dff (\oc8051_golden_model_1.TH1 [7], _40451_);
  dff (\oc8051_golden_model_1.TMOD [0], _43224_);
  dff (\oc8051_golden_model_1.TMOD [1], _43225_);
  dff (\oc8051_golden_model_1.TMOD [2], _43226_);
  dff (\oc8051_golden_model_1.TMOD [3], _43227_);
  dff (\oc8051_golden_model_1.TMOD [4], _43228_);
  dff (\oc8051_golden_model_1.TMOD [5], _43229_);
  dff (\oc8051_golden_model_1.TMOD [6], _43230_);
  dff (\oc8051_golden_model_1.TMOD [7], _40452_);
  dff (\oc8051_golden_model_1.IE [0], _43233_);
  dff (\oc8051_golden_model_1.IE [1], _43234_);
  dff (\oc8051_golden_model_1.IE [2], _43235_);
  dff (\oc8051_golden_model_1.IE [3], _43236_);
  dff (\oc8051_golden_model_1.IE [4], _43237_);
  dff (\oc8051_golden_model_1.IE [5], _43238_);
  dff (\oc8051_golden_model_1.IE [6], _43239_);
  dff (\oc8051_golden_model_1.IE [7], _40453_);
  dff (\oc8051_golden_model_1.IP [0], _43240_);
  dff (\oc8051_golden_model_1.IP [1], _43243_);
  dff (\oc8051_golden_model_1.IP [2], _43244_);
  dff (\oc8051_golden_model_1.IP [3], _43245_);
  dff (\oc8051_golden_model_1.IP [4], _43246_);
  dff (\oc8051_golden_model_1.IP [5], _43247_);
  dff (\oc8051_golden_model_1.IP [6], _43248_);
  dff (\oc8051_golden_model_1.IP [7], _40455_);
  dff (\oc8051_golden_model_1.DPL [0], _43251_);
  dff (\oc8051_golden_model_1.DPL [1], _43252_);
  dff (\oc8051_golden_model_1.DPL [2], _43253_);
  dff (\oc8051_golden_model_1.DPL [3], _43254_);
  dff (\oc8051_golden_model_1.DPL [4], _43255_);
  dff (\oc8051_golden_model_1.DPL [5], _43256_);
  dff (\oc8051_golden_model_1.DPL [6], _43257_);
  dff (\oc8051_golden_model_1.DPL [7], _40456_);
  dff (\oc8051_golden_model_1.DPH [0], _43258_);
  dff (\oc8051_golden_model_1.DPH [1], _43259_);
  dff (\oc8051_golden_model_1.DPH [2], _43260_);
  dff (\oc8051_golden_model_1.DPH [3], _43263_);
  dff (\oc8051_golden_model_1.DPH [4], _43264_);
  dff (\oc8051_golden_model_1.DPH [5], _43265_);
  dff (\oc8051_golden_model_1.DPH [6], _43266_);
  dff (\oc8051_golden_model_1.DPH [7], _40457_);
  dff (\oc8051_golden_model_1.PC [0], _43269_);
  dff (\oc8051_golden_model_1.PC [1], _43270_);
  dff (\oc8051_golden_model_1.PC [2], _43271_);
  dff (\oc8051_golden_model_1.PC [3], _43272_);
  dff (\oc8051_golden_model_1.PC [4], _43273_);
  dff (\oc8051_golden_model_1.PC [5], _43274_);
  dff (\oc8051_golden_model_1.PC [6], _43275_);
  dff (\oc8051_golden_model_1.PC [7], _43276_);
  dff (\oc8051_golden_model_1.PC [8], _43277_);
  dff (\oc8051_golden_model_1.PC [9], _43278_);
  dff (\oc8051_golden_model_1.PC [10], _43279_);
  dff (\oc8051_golden_model_1.PC [11], _43282_);
  dff (\oc8051_golden_model_1.PC [12], _43283_);
  dff (\oc8051_golden_model_1.PC [13], _43284_);
  dff (\oc8051_golden_model_1.PC [14], _43285_);
  dff (\oc8051_golden_model_1.PC [15], _40458_);
  dff (\oc8051_golden_model_1.P2 [0], _43288_);
  dff (\oc8051_golden_model_1.P2 [1], _43289_);
  dff (\oc8051_golden_model_1.P2 [2], _43290_);
  dff (\oc8051_golden_model_1.P2 [3], _43291_);
  dff (\oc8051_golden_model_1.P2 [4], _43292_);
  dff (\oc8051_golden_model_1.P2 [5], _43293_);
  dff (\oc8051_golden_model_1.P2 [6], _43294_);
  dff (\oc8051_golden_model_1.P2 [7], _40459_);
  dff (\oc8051_golden_model_1.P3 [0], _43295_);
  dff (\oc8051_golden_model_1.P3 [1], _43296_);
  dff (\oc8051_golden_model_1.P3 [2], _43297_);
  dff (\oc8051_golden_model_1.P3 [3], _43298_);
  dff (\oc8051_golden_model_1.P3 [4], _43299_);
  dff (\oc8051_golden_model_1.P3 [5], _43302_);
  dff (\oc8051_golden_model_1.P3 [6], _43303_);
  dff (\oc8051_golden_model_1.P3 [7], _40461_);
  dff (\oc8051_golden_model_1.P0 [0], _43304_);
  dff (\oc8051_golden_model_1.P0 [1], _43307_);
  dff (\oc8051_golden_model_1.P0 [2], _43308_);
  dff (\oc8051_golden_model_1.P0 [3], _43309_);
  dff (\oc8051_golden_model_1.P0 [4], _43310_);
  dff (\oc8051_golden_model_1.P0 [5], _43311_);
  dff (\oc8051_golden_model_1.P0 [6], _43312_);
  dff (\oc8051_golden_model_1.P0 [7], _40462_);
  dff (\oc8051_golden_model_1.P1 [0], _43313_);
  dff (\oc8051_golden_model_1.P1 [1], _43314_);
  dff (\oc8051_golden_model_1.P1 [2], _43315_);
  dff (\oc8051_golden_model_1.P1 [3], _43316_);
  dff (\oc8051_golden_model_1.P1 [4], _43317_);
  dff (\oc8051_golden_model_1.P1 [5], _43318_);
  dff (\oc8051_golden_model_1.P1 [6], _43319_);
  dff (\oc8051_golden_model_1.P1 [7], _40463_);
  dff (\oc8051_golden_model_1.SP [0], _43322_);
  dff (\oc8051_golden_model_1.SP [1], _43323_);
  dff (\oc8051_golden_model_1.SP [2], _43324_);
  dff (\oc8051_golden_model_1.SP [3], _43327_);
  dff (\oc8051_golden_model_1.SP [4], _43328_);
  dff (\oc8051_golden_model_1.SP [5], _43329_);
  dff (\oc8051_golden_model_1.SP [6], _43330_);
  dff (\oc8051_golden_model_1.SP [7], _40464_);
  dff (\oc8051_golden_model_1.PSW [0], _43331_);
  dff (\oc8051_golden_model_1.PSW [1], _43332_);
  dff (\oc8051_golden_model_1.PSW [2], _43333_);
  dff (\oc8051_golden_model_1.PSW [3], _43334_);
  dff (\oc8051_golden_model_1.PSW [4], _43335_);
  dff (\oc8051_golden_model_1.PSW [5], _43336_);
  dff (\oc8051_golden_model_1.PSW [6], _43337_);
  dff (\oc8051_golden_model_1.PSW [7], _40465_);
  dff (\oc8051_golden_model_1.P0INREG [0], _43340_);
  dff (\oc8051_golden_model_1.P0INREG [1], _43341_);
  dff (\oc8051_golden_model_1.P0INREG [2], _43342_);
  dff (\oc8051_golden_model_1.P0INREG [3], _43343_);
  dff (\oc8051_golden_model_1.P0INREG [4], _43344_);
  dff (\oc8051_golden_model_1.P0INREG [5], _43347_);
  dff (\oc8051_golden_model_1.P0INREG [6], _43348_);
  dff (\oc8051_golden_model_1.P0INREG [7], _40467_);
  dff (\oc8051_golden_model_1.P1INREG [0], _43349_);
  dff (\oc8051_golden_model_1.P1INREG [1], _43351_);
  dff (\oc8051_golden_model_1.P1INREG [2], _43352_);
  dff (\oc8051_golden_model_1.P1INREG [3], _43353_);
  dff (\oc8051_golden_model_1.P1INREG [4], _43354_);
  dff (\oc8051_golden_model_1.P1INREG [5], _43355_);
  dff (\oc8051_golden_model_1.P1INREG [6], _43356_);
  dff (\oc8051_golden_model_1.P1INREG [7], _40468_);
  dff (\oc8051_golden_model_1.P2INREG [0], _43359_);
  dff (\oc8051_golden_model_1.P2INREG [1], _43360_);
  dff (\oc8051_golden_model_1.P2INREG [2], _43361_);
  dff (\oc8051_golden_model_1.P2INREG [3], _43362_);
  dff (\oc8051_golden_model_1.P2INREG [4], _43363_);
  dff (\oc8051_golden_model_1.P2INREG [5], _43364_);
  dff (\oc8051_golden_model_1.P2INREG [6], _43365_);
  dff (\oc8051_golden_model_1.P2INREG [7], _40469_);
  dff (\oc8051_golden_model_1.P3INREG [0], _43367_);
  dff (\oc8051_golden_model_1.P3INREG [1], _43368_);
  dff (\oc8051_golden_model_1.P3INREG [2], _43369_);
  dff (\oc8051_golden_model_1.P3INREG [3], _43370_);
  dff (\oc8051_golden_model_1.P3INREG [4], _43371_);
  dff (\oc8051_golden_model_1.P3INREG [5], _43372_);
  dff (\oc8051_golden_model_1.P3INREG [6], _43373_);
  dff (\oc8051_golden_model_1.P3INREG [7], _40470_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02972_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02983_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03003_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03025_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03045_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00866_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03056_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00840_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03066_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03077_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03088_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03098_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03109_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03120_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03131_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00884_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02427_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22329_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02622_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02816_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03014_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03222_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03423_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03624_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03825_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04026_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04127_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04228_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04329_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04430_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04531_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04632_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04733_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24502_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38639_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38640_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38641_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38642_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38643_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38644_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38645_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38625_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38646_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38648_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38649_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38650_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38651_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38652_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38654_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38627_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38655_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38656_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38657_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38658_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38660_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38661_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38662_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38628_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _30380_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05965_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _30383_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05968_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _30385_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _30387_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05971_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _30389_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _30391_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05974_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _30393_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05977_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _30395_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _30397_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _30399_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _05980_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _30401_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05983_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _05986_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _06045_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _06047_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _05950_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _06050_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _06053_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _05953_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _06056_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _05956_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _06059_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _06062_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _06065_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _06068_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _06071_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _06074_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _06077_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _05959_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _05962_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39429_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _39462_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _39463_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _39464_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _39465_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _39466_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _39467_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _39468_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39430_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _39469_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _39470_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _39471_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _39472_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _39473_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _39474_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _39475_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39431_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _39476_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _39478_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _39479_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _39480_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _39481_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _39482_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _39483_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39433_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _39484_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _39485_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _39486_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _39487_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _39489_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _39490_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _39491_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39434_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39005_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39006_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39007_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39008_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38722_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38796_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38800_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38802_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38804_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38806_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38808_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _38810_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _38811_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38685_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _38815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _38816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _38817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _38818_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _38819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _38820_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _38821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _38822_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _38824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _38825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _38826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _38827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _38828_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _38829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _38830_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38687_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39009_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39010_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39012_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39013_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39014_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39015_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39016_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39017_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39018_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39019_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39020_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39021_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39023_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39024_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39025_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39026_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39027_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39028_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39029_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39030_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39031_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39032_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39034_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39035_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39036_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39037_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39038_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39039_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39040_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39041_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39042_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38746_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39044_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39045_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39046_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39047_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39048_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39050_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39051_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39052_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39053_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39054_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39057_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39060_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39061_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39062_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39063_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39064_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39065_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39066_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38726_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38727_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38728_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39068_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39069_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39071_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39072_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39073_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39074_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38729_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39075_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39076_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39077_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39078_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39079_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39080_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39082_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39083_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39084_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39085_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39086_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39087_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39088_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39090_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38731_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39091_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39093_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39094_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39095_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39096_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39097_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39098_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39099_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39100_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39101_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39102_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39104_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39105_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39106_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39107_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38732_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38735_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38734_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39108_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39109_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39110_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39111_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39112_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39113_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39115_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38736_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39116_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39117_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38737_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39118_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39119_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39120_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39122_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39123_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39124_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38738_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39126_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39127_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39128_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39129_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39132_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38739_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _38740_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39133_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39134_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39137_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39138_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39139_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39140_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38742_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _38743_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38744_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39141_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39143_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38745_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39144_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39145_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39149_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39151_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39152_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39153_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39155_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39156_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39159_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39160_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39163_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39165_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39167_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39169_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39171_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39173_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39176_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39178_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39181_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39182_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39183_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39184_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39187_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39189_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39191_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39192_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39195_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38753_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38754_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39203_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39209_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39213_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39214_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39216_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39217_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38756_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38757_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39636_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39655_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39656_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39657_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39659_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39660_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39661_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39662_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39638_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39639_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39663_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39664_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _43666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _43670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _43674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _43678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _43682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _43686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _43690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _42719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _43634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _43638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _43642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _43646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _43650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _43654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _43658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _43661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _43602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _43606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _43610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _43614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _43618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _43622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _43626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _43629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _42974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _42980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _42986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _42992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _42998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _43004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _43010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _43013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _43021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _43025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _43029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _43033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _43034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _43038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _43042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _43045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _43053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _43057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _43061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _43065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _43069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _43073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _43077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _43080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _43121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _43125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _43129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _43133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _43149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _43169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _43187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _43198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _43086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _43090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _43094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _43098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _43102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _43106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _43110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _43113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _43473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _43477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _43481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _43485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _43489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _43493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _43497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _43500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _43441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _43445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _43449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _43453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _43457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _43461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _43465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _43468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _43407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _43411_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _43415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _43419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _43423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _43427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _43431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _43434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _43375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _43379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _43383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _43387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _43391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _43395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _43399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _43402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _43223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _43242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _43262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _43281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _43301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _43321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _43339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _43350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _43505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _43509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _43513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _43517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _43521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _43525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _43529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _43532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _43570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _43574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _43578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _43582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _43586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _43590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _43594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _43597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _43537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _43541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _43545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _43549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _43553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _43557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _43561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _43564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _01364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _01366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _01368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _01370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _01372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _01374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _01376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _42707_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39521_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39522_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39586_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39587_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39589_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39590_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39591_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39592_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39593_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39523_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39524_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24099_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24123_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08887_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08898_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08908_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08941_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08952_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13619_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13628_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12656_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13667_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13676_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13686_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _41654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _42571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _42573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42574_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _42576_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _42578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _42580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42582_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _42584_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _41651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _41649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _42586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _42587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _41647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _42589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _42591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _41645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _42593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _42595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _41610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _41608_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _41606_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _41604_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _42597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _42599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _42601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _41601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _42603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _42604_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _42606_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _42608_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _42610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _42612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _42614_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _41599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _42616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _42618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _42620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _42622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _42624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _42626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _42628_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _41597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41059_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41061_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41062_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41068_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41069_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35388_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41071_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41073_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41076_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41080_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35411_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41089_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41092_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35434_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41095_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41097_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41099_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41101_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41103_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41106_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35457_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21381_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21392_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21404_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21416_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21428_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21439_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16448_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09497_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10676_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10687_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09517_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [0], \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [1], \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [2], \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [3], \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [4], \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [5], \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [6], \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [7], \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [0], \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [1], \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [2], \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [3], \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [4], \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [5], \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [6], \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [7], \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [0], \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [1], \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [2], \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [3], \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [4], \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [5], \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [6], \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [7], \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [0], \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [1], \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [2], \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [3], \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [4], \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [5], \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [6], \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [7], \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1283 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1300 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1439 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1439 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1489 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1475 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1489 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1489 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1569 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1605 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1605 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1638 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1638 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1671 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1671 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1732 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1732 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1732 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1732 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1732 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1732 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1732 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1789 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1806 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1823 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1823 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1866 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1866 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1866 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1866 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1866 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1866 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1866 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1923 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1940 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1957 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1957 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2074 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2091 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2108 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2108 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2132 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2148 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2190 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2148 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2216 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2216 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2148 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2457 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2457 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2457 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2457 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2487 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2487 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2487 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2487 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2517 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2517 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2552 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2555 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2583 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2583 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2589 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2629 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2682 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2735 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2735 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2823 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2823 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2845 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2845 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2864 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2735 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2881 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.n2882 [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.n2882 [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.n2882 [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.n2882 [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.n2882 [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.n2882 [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.n2882 [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0988 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n0988 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n0988 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0988 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0988 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n0988 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n0988 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0989 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0990 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0991 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0992 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0993 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0995 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0996 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1003 , \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1011 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1011 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1011 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1011 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1011 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1011 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1011 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1017 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1018 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1019 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1026 , \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.n1027 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1027 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1027 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1027 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1027 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1043 , \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.n1044 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1044 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1044 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1044 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1044 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1044 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1044 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1156 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1156 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1156 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1156 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1158 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1158 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1158 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1158 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1160 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1160 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1160 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1160 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1161 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1161 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1162 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1163 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1164 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1165 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1165 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1166 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1213 , \oc8051_golden_model_1.n2555 [7]);
  buf(\oc8051_golden_model_1.n1258 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1259 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1259 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1259 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1259 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1259 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1259 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1259 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1259 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1259 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1260 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1261 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1261 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1261 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1261 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1261 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1262 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1263 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1263 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1263 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1264 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1265 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1265 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1266 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1266 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1266 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1266 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1266 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1266 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1266 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1267 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1267 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1267 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1267 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1267 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1267 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1268 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1269 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1270 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1271 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1272 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1273 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1274 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1282 , \oc8051_golden_model_1.n1283 [0]);
  buf(\oc8051_golden_model_1.n1283 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1283 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1283 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1283 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1283 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1283 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1283 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1299 , \oc8051_golden_model_1.n1300 [0]);
  buf(\oc8051_golden_model_1.n1300 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1300 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1300 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1300 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1300 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1300 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1300 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1343 [9], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1343 [10], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1343 [11], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1343 [12], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.n1343 [13], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.n1343 [14], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.n1343 [15], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n1345 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1345 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1345 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1345 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1345 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1345 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1345 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1345 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1346 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1352 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1360 , \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.n1361 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1361 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1361 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1361 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1361 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1361 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1361 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1363 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1363 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1363 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1363 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1363 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1363 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1363 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1363 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1363 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1367 [8], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1368 , \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1369 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1369 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1370 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1370 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1370 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1374 [4], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1375 , \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1376 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1376 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1376 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1376 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1376 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1384 , \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1385 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1385 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1385 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1385 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1385 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1385 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1386 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1386 [1], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1386 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1386 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1386 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1386 [5], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1386 [6], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1401 , \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.n1402 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1402 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1402 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1402 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1406 [8], \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.n1407 , \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.n1412 [4], \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.n1413 , \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.n1421 , \oc8051_golden_model_1.n1439 [2]);
  buf(\oc8051_golden_model_1.n1422 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1422 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1422 [2], \oc8051_golden_model_1.n1439 [2]);
  buf(\oc8051_golden_model_1.n1422 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1422 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1422 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1422 [6], \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.n1422 [7], \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.n1423 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1423 [1], \oc8051_golden_model_1.n1439 [2]);
  buf(\oc8051_golden_model_1.n1423 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1423 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1423 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1423 [5], \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.n1423 [6], \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.n1438 , \oc8051_golden_model_1.n1439 [0]);
  buf(\oc8051_golden_model_1.n1439 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1439 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1439 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1439 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1441 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1441 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1441 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1441 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1441 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n1441 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n1441 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n1441 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n1441 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1443 [8], \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.n1444 , \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.n1445 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1445 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1445 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1445 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1446 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1446 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1446 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1446 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1446 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1448 [4], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1449 , \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1450 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1450 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1450 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1450 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1450 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n1450 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n1450 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n1450 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n1450 [8], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n1457 , \oc8051_golden_model_1.n1475 [2]);
  buf(\oc8051_golden_model_1.n1458 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1458 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1458 [2], \oc8051_golden_model_1.n1475 [2]);
  buf(\oc8051_golden_model_1.n1458 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1458 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1458 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1458 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1458 [7], \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.n1459 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1459 [1], \oc8051_golden_model_1.n1475 [2]);
  buf(\oc8051_golden_model_1.n1459 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1459 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1459 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1459 [5], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1459 [6], \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.n1474 , \oc8051_golden_model_1.n1489 [0]);
  buf(\oc8051_golden_model_1.n1475 [0], \oc8051_golden_model_1.n1489 [0]);
  buf(\oc8051_golden_model_1.n1475 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1475 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1475 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1475 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1475 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1478 [8], \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.n1479 , \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.n1486 , \oc8051_golden_model_1.n1489 [2]);
  buf(\oc8051_golden_model_1.n1487 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1487 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1487 [2], \oc8051_golden_model_1.n1489 [2]);
  buf(\oc8051_golden_model_1.n1487 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1487 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1487 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1487 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1487 [7], \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.n1488 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1488 [1], \oc8051_golden_model_1.n1489 [2]);
  buf(\oc8051_golden_model_1.n1488 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1488 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1488 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1488 [5], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1488 [6], \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.n1489 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1489 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1489 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1489 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1491 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1491 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1491 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1491 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1491 [4], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.n1491 [5], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.n1491 [6], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.n1491 [7], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n1491 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1493 [8], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1494 , \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1495 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1495 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1495 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1495 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1495 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1497 [4], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1498 , \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1499 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1499 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1499 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1499 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1499 [4], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.n1499 [5], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.n1499 [6], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.n1499 [7], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n1499 [8], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n1506 , \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1507 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1507 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1507 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1507 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1508 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1508 [1], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1508 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1508 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1508 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1508 [5], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1508 [6], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1523 , \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.n1524 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.n1524 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1524 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1524 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1524 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1524 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1524 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1524 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1527 , \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1528 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1528 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1528 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1528 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1528 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1528 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1528 [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1528 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1529 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1529 [1], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1529 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1529 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1529 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1529 [5], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1529 [6], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1530 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.n1530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1530 [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1532 [8], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1533 , \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1540 , \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1541 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1541 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1541 [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1541 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1541 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1541 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1541 [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1541 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1543 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.n1543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1543 [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1543 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1544 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1544 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1544 [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1544 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1544 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1544 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1544 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1545 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1545 [1], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1545 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1545 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1545 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1545 [5], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1545 [6], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1549 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1549 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1549 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1549 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1549 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1549 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1549 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1549 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1549 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1550 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1550 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1550 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1550 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1550 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1550 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1550 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1550 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1550 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1551 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1551 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1551 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1551 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1551 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1551 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1551 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1551 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1552 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1552 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1552 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1552 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1552 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1552 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1552 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1552 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1553 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1553 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1553 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1553 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1553 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1553 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1553 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1555 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1557 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1559 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1560 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1561 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 , \oc8051_golden_model_1.n1569 [0]);
  buf(\oc8051_golden_model_1.n1569 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1569 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1569 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1569 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1569 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1569 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1569 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1570 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1573 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [8], \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.n1576 , \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.n1577 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1577 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1579 [4], \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.n1580 , \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.n1587 , \oc8051_golden_model_1.n1605 [2]);
  buf(\oc8051_golden_model_1.n1588 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1588 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1588 [2], \oc8051_golden_model_1.n1605 [2]);
  buf(\oc8051_golden_model_1.n1588 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1588 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1588 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1588 [6], \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.n1588 [7], \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.n1589 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1589 [1], \oc8051_golden_model_1.n1605 [2]);
  buf(\oc8051_golden_model_1.n1589 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1589 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1589 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1589 [5], \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.n1589 [6], \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.n1604 , \oc8051_golden_model_1.n1605 [0]);
  buf(\oc8051_golden_model_1.n1605 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1605 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1605 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1605 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1609 [8], \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.n1610 , \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.n1612 [4], \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.n1613 , \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.n1620 , \oc8051_golden_model_1.n1638 [2]);
  buf(\oc8051_golden_model_1.n1621 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1621 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1621 [2], \oc8051_golden_model_1.n1638 [2]);
  buf(\oc8051_golden_model_1.n1621 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1621 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1621 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1621 [6], \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.n1621 [7], \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.n1622 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1622 [1], \oc8051_golden_model_1.n1638 [2]);
  buf(\oc8051_golden_model_1.n1622 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1622 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1622 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1622 [5], \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.n1622 [6], \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.n1637 , \oc8051_golden_model_1.n1638 [0]);
  buf(\oc8051_golden_model_1.n1638 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1638 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1638 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1638 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1642 [8], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.n1643 , \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.n1645 [4], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.n1646 , \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.n1653 , \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.n1654 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1654 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1654 [2], \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.n1654 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1654 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1654 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1654 [6], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.n1654 [7], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.n1655 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1655 [1], \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.n1655 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1655 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1655 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1655 [5], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.n1655 [6], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.n1670 , \oc8051_golden_model_1.n1671 [0]);
  buf(\oc8051_golden_model_1.n1671 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1671 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1671 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1671 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1675 [8], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.n1676 , \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.n1678 [4], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.n1679 , \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.n1686 , \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.n1687 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1687 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1687 [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.n1687 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1687 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1687 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1687 [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.n1687 [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.n1688 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1688 [1], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.n1688 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1688 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1688 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1688 [5], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.n1688 [6], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.n1703 , \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.n1704 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1704 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1704 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1704 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1730 [1], \oc8051_golden_model_1.n1732 [1]);
  buf(\oc8051_golden_model_1.n1730 [2], \oc8051_golden_model_1.n1732 [2]);
  buf(\oc8051_golden_model_1.n1730 [3], \oc8051_golden_model_1.n1732 [3]);
  buf(\oc8051_golden_model_1.n1730 [4], \oc8051_golden_model_1.n1732 [4]);
  buf(\oc8051_golden_model_1.n1730 [5], \oc8051_golden_model_1.n1732 [5]);
  buf(\oc8051_golden_model_1.n1730 [6], \oc8051_golden_model_1.n1732 [6]);
  buf(\oc8051_golden_model_1.n1730 [7], \oc8051_golden_model_1.n1732 [7]);
  buf(\oc8051_golden_model_1.n1731 [0], \oc8051_golden_model_1.n1732 [1]);
  buf(\oc8051_golden_model_1.n1731 [1], \oc8051_golden_model_1.n1732 [2]);
  buf(\oc8051_golden_model_1.n1731 [2], \oc8051_golden_model_1.n1732 [3]);
  buf(\oc8051_golden_model_1.n1731 [3], \oc8051_golden_model_1.n1732 [4]);
  buf(\oc8051_golden_model_1.n1731 [4], \oc8051_golden_model_1.n1732 [5]);
  buf(\oc8051_golden_model_1.n1731 [5], \oc8051_golden_model_1.n1732 [6]);
  buf(\oc8051_golden_model_1.n1731 [6], \oc8051_golden_model_1.n1732 [7]);
  buf(\oc8051_golden_model_1.n1732 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n1788 , \oc8051_golden_model_1.n1789 [0]);
  buf(\oc8051_golden_model_1.n1789 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1789 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1789 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1789 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1789 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1789 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1789 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1805 , \oc8051_golden_model_1.n1806 [0]);
  buf(\oc8051_golden_model_1.n1806 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1806 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1806 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1806 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1806 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1806 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1806 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1822 , \oc8051_golden_model_1.n1823 [0]);
  buf(\oc8051_golden_model_1.n1823 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1823 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1823 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1823 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1823 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1823 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1823 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1839 , \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.n1840 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1840 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1840 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1840 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1840 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1840 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1840 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1864 [1], \oc8051_golden_model_1.n1866 [1]);
  buf(\oc8051_golden_model_1.n1864 [2], \oc8051_golden_model_1.n1866 [2]);
  buf(\oc8051_golden_model_1.n1864 [3], \oc8051_golden_model_1.n1866 [3]);
  buf(\oc8051_golden_model_1.n1864 [4], \oc8051_golden_model_1.n1866 [4]);
  buf(\oc8051_golden_model_1.n1864 [5], \oc8051_golden_model_1.n1866 [5]);
  buf(\oc8051_golden_model_1.n1864 [6], \oc8051_golden_model_1.n1866 [6]);
  buf(\oc8051_golden_model_1.n1864 [7], \oc8051_golden_model_1.n1866 [7]);
  buf(\oc8051_golden_model_1.n1865 [0], \oc8051_golden_model_1.n1866 [1]);
  buf(\oc8051_golden_model_1.n1865 [1], \oc8051_golden_model_1.n1866 [2]);
  buf(\oc8051_golden_model_1.n1865 [2], \oc8051_golden_model_1.n1866 [3]);
  buf(\oc8051_golden_model_1.n1865 [3], \oc8051_golden_model_1.n1866 [4]);
  buf(\oc8051_golden_model_1.n1865 [4], \oc8051_golden_model_1.n1866 [5]);
  buf(\oc8051_golden_model_1.n1865 [5], \oc8051_golden_model_1.n1866 [6]);
  buf(\oc8051_golden_model_1.n1865 [6], \oc8051_golden_model_1.n1866 [7]);
  buf(\oc8051_golden_model_1.n1866 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n1922 , \oc8051_golden_model_1.n1923 [0]);
  buf(\oc8051_golden_model_1.n1923 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1923 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1923 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1923 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1923 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1923 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1923 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1939 , \oc8051_golden_model_1.n1940 [0]);
  buf(\oc8051_golden_model_1.n1940 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1940 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1940 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1940 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1940 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1940 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1940 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1956 , \oc8051_golden_model_1.n1957 [0]);
  buf(\oc8051_golden_model_1.n1957 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1957 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1957 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1957 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1957 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1957 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1957 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1973 , \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.n1974 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1974 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1974 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1974 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1974 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1974 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1974 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2073 , \oc8051_golden_model_1.n2074 [0]);
  buf(\oc8051_golden_model_1.n2074 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2074 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2074 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2074 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2074 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2074 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2074 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2090 , \oc8051_golden_model_1.n2091 [0]);
  buf(\oc8051_golden_model_1.n2091 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2091 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2091 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2091 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2091 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2091 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2091 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2107 , \oc8051_golden_model_1.n2108 [0]);
  buf(\oc8051_golden_model_1.n2108 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2108 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2108 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2108 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2108 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2108 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2108 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2124 , \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.n2125 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2125 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2125 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2125 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2125 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2125 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2125 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2128 , \oc8051_golden_model_1.n2132 [7]);
  buf(\oc8051_golden_model_1.n2129 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2129 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2129 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2129 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2129 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2129 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2129 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2130 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2130 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2130 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2130 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2130 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2130 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2130 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2130 [7], \oc8051_golden_model_1.n2132 [7]);
  buf(\oc8051_golden_model_1.n2131 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2131 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2131 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2131 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2131 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2131 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2131 [6], \oc8051_golden_model_1.n2132 [7]);
  buf(\oc8051_golden_model_1.n2132 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2132 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2132 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2132 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2132 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2132 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2132 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2147 , \oc8051_golden_model_1.n2148 [0]);
  buf(\oc8051_golden_model_1.n2148 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2148 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2148 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2148 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2148 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2148 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2148 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2187 , \oc8051_golden_model_1.n2190 [7]);
  buf(\oc8051_golden_model_1.n2188 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2188 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2188 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2188 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2188 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2188 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2188 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2188 [7], \oc8051_golden_model_1.n2190 [7]);
  buf(\oc8051_golden_model_1.n2189 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2189 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2189 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2189 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2189 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2189 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2189 [6], \oc8051_golden_model_1.n2190 [7]);
  buf(\oc8051_golden_model_1.n2190 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2190 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2190 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2190 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2190 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2190 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2190 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2197 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2197 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2197 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2197 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2198 , \oc8051_golden_model_1.n2216 [2]);
  buf(\oc8051_golden_model_1.n2199 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2199 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2199 [2], \oc8051_golden_model_1.n2216 [2]);
  buf(\oc8051_golden_model_1.n2199 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2199 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2199 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2199 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2199 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2200 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2200 [1], \oc8051_golden_model_1.n2216 [2]);
  buf(\oc8051_golden_model_1.n2200 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2200 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2200 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2200 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2200 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2215 , \oc8051_golden_model_1.n2216 [0]);
  buf(\oc8051_golden_model_1.n2216 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2216 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2216 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2216 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2216 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2216 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2428 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2431 , \oc8051_golden_model_1.n2457 [7]);
  buf(\oc8051_golden_model_1.n2433 , \oc8051_golden_model_1.n2457 [6]);
  buf(\oc8051_golden_model_1.n2439 , \oc8051_golden_model_1.n2457 [2]);
  buf(\oc8051_golden_model_1.n2440 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2440 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2440 [2], \oc8051_golden_model_1.n2457 [2]);
  buf(\oc8051_golden_model_1.n2440 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2440 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2440 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2440 [6], \oc8051_golden_model_1.n2457 [6]);
  buf(\oc8051_golden_model_1.n2440 [7], \oc8051_golden_model_1.n2457 [7]);
  buf(\oc8051_golden_model_1.n2441 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2441 [1], \oc8051_golden_model_1.n2457 [2]);
  buf(\oc8051_golden_model_1.n2441 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2441 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2441 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2441 [5], \oc8051_golden_model_1.n2457 [6]);
  buf(\oc8051_golden_model_1.n2441 [6], \oc8051_golden_model_1.n2457 [7]);
  buf(\oc8051_golden_model_1.n2456 , \oc8051_golden_model_1.n2457 [0]);
  buf(\oc8051_golden_model_1.n2457 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2457 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2457 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2457 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2461 , \oc8051_golden_model_1.n2487 [7]);
  buf(\oc8051_golden_model_1.n2463 , \oc8051_golden_model_1.n2487 [6]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2487 [2]);
  buf(\oc8051_golden_model_1.n2470 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [2], \oc8051_golden_model_1.n2487 [2]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2470 [6], \oc8051_golden_model_1.n2487 [6]);
  buf(\oc8051_golden_model_1.n2470 [7], \oc8051_golden_model_1.n2487 [7]);
  buf(\oc8051_golden_model_1.n2471 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2471 [1], \oc8051_golden_model_1.n2487 [2]);
  buf(\oc8051_golden_model_1.n2471 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2471 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2471 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2471 [5], \oc8051_golden_model_1.n2487 [6]);
  buf(\oc8051_golden_model_1.n2471 [6], \oc8051_golden_model_1.n2487 [7]);
  buf(\oc8051_golden_model_1.n2486 , \oc8051_golden_model_1.n2487 [0]);
  buf(\oc8051_golden_model_1.n2487 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2487 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2487 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2487 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2491 , \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2493 , \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.n2499 , \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.n2500 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [2], \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2500 [6], \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.n2500 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2501 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2501 [1], \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.n2501 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2501 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2501 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2501 [5], \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.n2501 [6], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2516 , \oc8051_golden_model_1.n2517 [0]);
  buf(\oc8051_golden_model_1.n2517 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2517 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2517 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2517 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2521 , \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.n2523 , \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.n2530 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2530 [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.n2530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2530 [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.n2530 [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.n2531 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2531 [1], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.n2531 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2531 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2531 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2531 [5], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.n2531 [6], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.n2546 , \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2549 , \oc8051_golden_model_1.n2552 [7]);
  buf(\oc8051_golden_model_1.n2550 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2550 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2550 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2550 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2550 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2550 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2550 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2550 [7], \oc8051_golden_model_1.n2552 [7]);
  buf(\oc8051_golden_model_1.n2551 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2551 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2551 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2551 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2551 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2551 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2551 [6], \oc8051_golden_model_1.n2552 [7]);
  buf(\oc8051_golden_model_1.n2552 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2552 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2552 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2552 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2552 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2552 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2552 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2553 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2553 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2553 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2553 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2553 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2553 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2553 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2553 [7], \oc8051_golden_model_1.n2555 [7]);
  buf(\oc8051_golden_model_1.n2554 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2554 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2554 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2554 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2554 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2554 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2554 [6], \oc8051_golden_model_1.n2555 [7]);
  buf(\oc8051_golden_model_1.n2555 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2555 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2555 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2555 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2555 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2555 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2555 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2559 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2559 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2559 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2559 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2559 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2559 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2559 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2559 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2559 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2565 , \oc8051_golden_model_1.n2583 [2]);
  buf(\oc8051_golden_model_1.n2566 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.n2583 [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2567 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2567 [1], \oc8051_golden_model_1.n2583 [2]);
  buf(\oc8051_golden_model_1.n2567 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2567 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2567 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2567 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2567 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2582 , \oc8051_golden_model_1.n2583 [0]);
  buf(\oc8051_golden_model_1.n2583 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2583 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2583 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2583 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2583 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2583 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2586 , \oc8051_golden_model_1.n2589 [7]);
  buf(\oc8051_golden_model_1.n2587 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2587 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2587 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2587 [7], \oc8051_golden_model_1.n2589 [7]);
  buf(\oc8051_golden_model_1.n2588 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2588 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2588 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2588 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2588 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2588 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2588 [6], \oc8051_golden_model_1.n2589 [7]);
  buf(\oc8051_golden_model_1.n2589 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2589 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2589 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2589 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2589 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2589 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2589 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2626 , \oc8051_golden_model_1.n2629 [7]);
  buf(\oc8051_golden_model_1.n2627 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2627 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2627 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2627 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2627 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2627 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2627 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2627 [7], \oc8051_golden_model_1.n2629 [7]);
  buf(\oc8051_golden_model_1.n2628 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2628 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2628 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2628 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2628 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2628 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2628 [6], \oc8051_golden_model_1.n2629 [7]);
  buf(\oc8051_golden_model_1.n2629 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2629 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2629 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2629 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2629 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2629 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2629 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2634 , \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2635 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2635 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2635 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2635 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2635 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2635 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2635 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2635 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2636 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2636 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2636 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2636 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2636 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2636 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2636 [6], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2637 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2637 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2637 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2637 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2637 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2637 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2637 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2642 , \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2643 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2643 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2643 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2643 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2643 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2643 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2643 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2644 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2644 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2644 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2644 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2644 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2644 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2644 [6], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2645 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2645 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2645 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2645 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2645 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2645 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2645 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2650 , \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2651 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2651 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2651 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2651 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2651 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2651 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2651 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2651 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2658 , \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2659 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2659 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2659 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2659 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2659 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2659 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2659 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2659 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2660 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2660 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2660 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2660 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2660 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2660 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2660 [6], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2661 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2661 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2661 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2661 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2661 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2661 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2661 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2662 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2662 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2662 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2662 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2662 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2662 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2662 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2662 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2663 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2663 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2663 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2663 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2663 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2663 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2663 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2664 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2664 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2664 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2664 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2664 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2664 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2664 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2664 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2665 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2665 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2665 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2665 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2666 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2666 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2666 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2666 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2666 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2666 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2666 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2666 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2667 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2668 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2669 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2670 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2671 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2672 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2673 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2674 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2681 , \oc8051_golden_model_1.n2682 [0]);
  buf(\oc8051_golden_model_1.n2682 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2682 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2682 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2682 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2682 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2682 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2682 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2702 [1], \oc8051_golden_model_1.n2882 [1]);
  buf(\oc8051_golden_model_1.n2702 [2], \oc8051_golden_model_1.n2882 [2]);
  buf(\oc8051_golden_model_1.n2702 [3], \oc8051_golden_model_1.n2882 [3]);
  buf(\oc8051_golden_model_1.n2702 [4], \oc8051_golden_model_1.n2882 [4]);
  buf(\oc8051_golden_model_1.n2702 [5], \oc8051_golden_model_1.n2882 [5]);
  buf(\oc8051_golden_model_1.n2702 [6], \oc8051_golden_model_1.n2882 [6]);
  buf(\oc8051_golden_model_1.n2702 [7], \oc8051_golden_model_1.n2882 [7]);
  buf(\oc8051_golden_model_1.n2703 [0], \oc8051_golden_model_1.n2882 [1]);
  buf(\oc8051_golden_model_1.n2703 [1], \oc8051_golden_model_1.n2882 [2]);
  buf(\oc8051_golden_model_1.n2703 [2], \oc8051_golden_model_1.n2882 [3]);
  buf(\oc8051_golden_model_1.n2703 [3], \oc8051_golden_model_1.n2882 [4]);
  buf(\oc8051_golden_model_1.n2703 [4], \oc8051_golden_model_1.n2882 [5]);
  buf(\oc8051_golden_model_1.n2703 [5], \oc8051_golden_model_1.n2882 [6]);
  buf(\oc8051_golden_model_1.n2703 [6], \oc8051_golden_model_1.n2882 [7]);
  buf(\oc8051_golden_model_1.n2719 [1], \oc8051_golden_model_1.n2882 [1]);
  buf(\oc8051_golden_model_1.n2719 [2], \oc8051_golden_model_1.n2882 [2]);
  buf(\oc8051_golden_model_1.n2719 [3], \oc8051_golden_model_1.n2882 [3]);
  buf(\oc8051_golden_model_1.n2719 [4], \oc8051_golden_model_1.n2882 [4]);
  buf(\oc8051_golden_model_1.n2719 [5], \oc8051_golden_model_1.n2882 [5]);
  buf(\oc8051_golden_model_1.n2719 [6], \oc8051_golden_model_1.n2882 [6]);
  buf(\oc8051_golden_model_1.n2719 [7], \oc8051_golden_model_1.n2882 [7]);
  buf(\oc8051_golden_model_1.n2720 , \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n2721 , \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n2722 , \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n2723 , \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n2724 , \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n2725 , \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n2726 , \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n2727 , \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n2734 , \oc8051_golden_model_1.n2735 [0]);
  buf(\oc8051_golden_model_1.n2735 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2735 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2735 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2735 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2735 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2735 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2735 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2750 , \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2751 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2751 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2751 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2751 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2751 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2751 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2751 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2784 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2784 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2784 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2784 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2784 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2784 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2784 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2784 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2785 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2785 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2785 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2785 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2785 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2785 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2785 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2786 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2786 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2786 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2786 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2786 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2786 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2786 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2786 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2805 , \oc8051_golden_model_1.n2823 [7]);
  buf(\oc8051_golden_model_1.n2806 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2806 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2806 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2806 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2806 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2806 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2806 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2806 [7], \oc8051_golden_model_1.n2823 [7]);
  buf(\oc8051_golden_model_1.n2807 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2807 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2807 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2807 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2807 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2807 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2807 [6], \oc8051_golden_model_1.n2823 [7]);
  buf(\oc8051_golden_model_1.n2822 , \oc8051_golden_model_1.n2823 [0]);
  buf(\oc8051_golden_model_1.n2823 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2823 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2823 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2823 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2823 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2823 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2827 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n2827 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n2827 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n2827 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n2827 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2827 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2827 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2827 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2828 [0], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n2828 [1], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n2828 [2], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n2828 [3], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n2829 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2829 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2829 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2829 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2830 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2831 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2832 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2833 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2844 , \oc8051_golden_model_1.n2845 [0]);
  buf(\oc8051_golden_model_1.n2845 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2845 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2845 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2845 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2845 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2845 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2845 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2863 , \oc8051_golden_model_1.n2864 [0]);
  buf(\oc8051_golden_model_1.n2864 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2864 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2864 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2864 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2864 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2864 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2864 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2880 , \oc8051_golden_model_1.n2881 [0]);
  buf(\oc8051_golden_model_1.n2881 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2881 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2881 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2881 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2881 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2881 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2881 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(ie_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(ie_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(ie_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(ie_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(ie_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(ie_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(ie_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(ie_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
