
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire _44029_;
  wire _44030_;
  wire _44031_;
  wire _44032_;
  wire _44033_;
  wire _44034_;
  wire _44035_;
  wire _44036_;
  wire _44037_;
  wire _44038_;
  wire _44039_;
  wire _44040_;
  wire _44041_;
  wire _44042_;
  wire _44043_;
  wire _44044_;
  wire _44045_;
  wire _44046_;
  wire _44047_;
  wire _44048_;
  wire _44049_;
  wire _44050_;
  wire _44051_;
  wire _44052_;
  wire _44053_;
  wire _44054_;
  wire _44055_;
  wire _44056_;
  wire _44057_;
  wire _44058_;
  wire _44059_;
  wire _44060_;
  wire _44061_;
  wire _44062_;
  wire _44063_;
  wire _44064_;
  wire _44065_;
  wire _44066_;
  wire _44067_;
  wire _44068_;
  wire _44069_;
  wire _44070_;
  wire _44071_;
  wire _44072_;
  wire _44073_;
  wire _44074_;
  wire _44075_;
  wire _44076_;
  wire _44077_;
  wire _44078_;
  wire _44079_;
  wire _44080_;
  wire _44081_;
  wire _44082_;
  wire _44083_;
  wire _44084_;
  wire _44085_;
  wire _44086_;
  wire _44087_;
  wire _44088_;
  wire _44089_;
  wire _44090_;
  wire _44091_;
  wire _44092_;
  wire _44093_;
  wire _44094_;
  wire _44095_;
  wire _44096_;
  wire _44097_;
  wire _44098_;
  wire _44099_;
  wire _44100_;
  wire _44101_;
  wire _44102_;
  wire _44103_;
  wire _44104_;
  wire _44105_;
  wire _44106_;
  wire _44107_;
  wire _44108_;
  wire _44109_;
  wire _44110_;
  wire _44111_;
  wire _44112_;
  wire _44113_;
  wire _44114_;
  wire _44115_;
  wire _44116_;
  wire _44117_;
  wire _44118_;
  wire _44119_;
  wire _44120_;
  wire _44121_;
  wire _44122_;
  wire _44123_;
  wire _44124_;
  wire _44125_;
  wire _44126_;
  wire _44127_;
  wire _44128_;
  wire _44129_;
  wire _44130_;
  wire _44131_;
  wire _44132_;
  wire _44133_;
  wire _44134_;
  wire _44135_;
  wire _44136_;
  wire _44137_;
  wire _44138_;
  wire _44139_;
  wire _44140_;
  wire _44141_;
  wire _44142_;
  wire _44143_;
  wire _44144_;
  wire _44145_;
  wire _44146_;
  wire _44147_;
  wire _44148_;
  wire _44149_;
  wire _44150_;
  wire _44151_;
  wire _44152_;
  wire [7:0] ACC_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] PCON_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [7:0] ie_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [6:0] \oc8051_golden_model_1.n0988 ;
  wire \oc8051_golden_model_1.n0989 ;
  wire \oc8051_golden_model_1.n0990 ;
  wire \oc8051_golden_model_1.n0991 ;
  wire \oc8051_golden_model_1.n0992 ;
  wire \oc8051_golden_model_1.n0993 ;
  wire \oc8051_golden_model_1.n0994 ;
  wire \oc8051_golden_model_1.n0995 ;
  wire \oc8051_golden_model_1.n0996 ;
  wire \oc8051_golden_model_1.n1003 ;
  wire [7:0] \oc8051_golden_model_1.n1004 ;
  wire [7:0] \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1017 ;
  wire \oc8051_golden_model_1.n1018 ;
  wire \oc8051_golden_model_1.n1019 ;
  wire \oc8051_golden_model_1.n1026 ;
  wire [7:0] \oc8051_golden_model_1.n1027 ;
  wire \oc8051_golden_model_1.n1043 ;
  wire [7:0] \oc8051_golden_model_1.n1044 ;
  wire [3:0] \oc8051_golden_model_1.n1156 ;
  wire [3:0] \oc8051_golden_model_1.n1158 ;
  wire [3:0] \oc8051_golden_model_1.n1160 ;
  wire [3:0] \oc8051_golden_model_1.n1161 ;
  wire [3:0] \oc8051_golden_model_1.n1162 ;
  wire [3:0] \oc8051_golden_model_1.n1163 ;
  wire [3:0] \oc8051_golden_model_1.n1164 ;
  wire [3:0] \oc8051_golden_model_1.n1165 ;
  wire [3:0] \oc8051_golden_model_1.n1166 ;
  wire \oc8051_golden_model_1.n1213 ;
  wire \oc8051_golden_model_1.n1258 ;
  wire [8:0] \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [7:0] \oc8051_golden_model_1.n1261 ;
  wire \oc8051_golden_model_1.n1262 ;
  wire [2:0] \oc8051_golden_model_1.n1263 ;
  wire \oc8051_golden_model_1.n1264 ;
  wire [1:0] \oc8051_golden_model_1.n1265 ;
  wire [7:0] \oc8051_golden_model_1.n1266 ;
  wire [6:0] \oc8051_golden_model_1.n1267 ;
  wire \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1270 ;
  wire \oc8051_golden_model_1.n1271 ;
  wire \oc8051_golden_model_1.n1272 ;
  wire \oc8051_golden_model_1.n1273 ;
  wire \oc8051_golden_model_1.n1274 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire \oc8051_golden_model_1.n1282 ;
  wire [7:0] \oc8051_golden_model_1.n1283 ;
  wire \oc8051_golden_model_1.n1299 ;
  wire [7:0] \oc8051_golden_model_1.n1300 ;
  wire [15:0] \oc8051_golden_model_1.n1343 ;
  wire [7:0] \oc8051_golden_model_1.n1345 ;
  wire \oc8051_golden_model_1.n1346 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1360 ;
  wire [7:0] \oc8051_golden_model_1.n1361 ;
  wire [8:0] \oc8051_golden_model_1.n1363 ;
  wire [8:0] \oc8051_golden_model_1.n1367 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [3:0] \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1370 ;
  wire [4:0] \oc8051_golden_model_1.n1374 ;
  wire \oc8051_golden_model_1.n1375 ;
  wire [8:0] \oc8051_golden_model_1.n1376 ;
  wire \oc8051_golden_model_1.n1384 ;
  wire [7:0] \oc8051_golden_model_1.n1385 ;
  wire [6:0] \oc8051_golden_model_1.n1386 ;
  wire \oc8051_golden_model_1.n1401 ;
  wire [7:0] \oc8051_golden_model_1.n1402 ;
  wire [8:0] \oc8051_golden_model_1.n1406 ;
  wire \oc8051_golden_model_1.n1407 ;
  wire [4:0] \oc8051_golden_model_1.n1412 ;
  wire \oc8051_golden_model_1.n1413 ;
  wire \oc8051_golden_model_1.n1421 ;
  wire [7:0] \oc8051_golden_model_1.n1422 ;
  wire [6:0] \oc8051_golden_model_1.n1423 ;
  wire \oc8051_golden_model_1.n1438 ;
  wire [7:0] \oc8051_golden_model_1.n1439 ;
  wire [8:0] \oc8051_golden_model_1.n1441 ;
  wire [8:0] \oc8051_golden_model_1.n1443 ;
  wire \oc8051_golden_model_1.n1444 ;
  wire [3:0] \oc8051_golden_model_1.n1445 ;
  wire [4:0] \oc8051_golden_model_1.n1446 ;
  wire [4:0] \oc8051_golden_model_1.n1448 ;
  wire \oc8051_golden_model_1.n1449 ;
  wire [8:0] \oc8051_golden_model_1.n1450 ;
  wire \oc8051_golden_model_1.n1457 ;
  wire [7:0] \oc8051_golden_model_1.n1458 ;
  wire [6:0] \oc8051_golden_model_1.n1459 ;
  wire \oc8051_golden_model_1.n1474 ;
  wire [7:0] \oc8051_golden_model_1.n1475 ;
  wire [8:0] \oc8051_golden_model_1.n1478 ;
  wire \oc8051_golden_model_1.n1479 ;
  wire \oc8051_golden_model_1.n1486 ;
  wire [7:0] \oc8051_golden_model_1.n1487 ;
  wire [6:0] \oc8051_golden_model_1.n1488 ;
  wire [7:0] \oc8051_golden_model_1.n1489 ;
  wire [8:0] \oc8051_golden_model_1.n1491 ;
  wire [8:0] \oc8051_golden_model_1.n1493 ;
  wire \oc8051_golden_model_1.n1494 ;
  wire [4:0] \oc8051_golden_model_1.n1495 ;
  wire [4:0] \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1498 ;
  wire [8:0] \oc8051_golden_model_1.n1499 ;
  wire \oc8051_golden_model_1.n1506 ;
  wire [7:0] \oc8051_golden_model_1.n1507 ;
  wire [6:0] \oc8051_golden_model_1.n1508 ;
  wire \oc8051_golden_model_1.n1523 ;
  wire [7:0] \oc8051_golden_model_1.n1524 ;
  wire [4:0] \oc8051_golden_model_1.n1526 ;
  wire \oc8051_golden_model_1.n1527 ;
  wire [7:0] \oc8051_golden_model_1.n1528 ;
  wire [6:0] \oc8051_golden_model_1.n1529 ;
  wire [7:0] \oc8051_golden_model_1.n1530 ;
  wire [8:0] \oc8051_golden_model_1.n1532 ;
  wire \oc8051_golden_model_1.n1533 ;
  wire \oc8051_golden_model_1.n1540 ;
  wire [7:0] \oc8051_golden_model_1.n1541 ;
  wire [6:0] \oc8051_golden_model_1.n1542 ;
  wire [7:0] \oc8051_golden_model_1.n1543 ;
  wire [7:0] \oc8051_golden_model_1.n1544 ;
  wire [6:0] \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [8:0] \oc8051_golden_model_1.n1549 ;
  wire [8:0] \oc8051_golden_model_1.n1550 ;
  wire [7:0] \oc8051_golden_model_1.n1551 ;
  wire [7:0] \oc8051_golden_model_1.n1552 ;
  wire [6:0] \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire \oc8051_golden_model_1.n1555 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire \oc8051_golden_model_1.n1557 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1559 ;
  wire \oc8051_golden_model_1.n1560 ;
  wire \oc8051_golden_model_1.n1561 ;
  wire \oc8051_golden_model_1.n1568 ;
  wire [7:0] \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [8:0] \oc8051_golden_model_1.n1573 ;
  wire [8:0] \oc8051_golden_model_1.n1575 ;
  wire \oc8051_golden_model_1.n1576 ;
  wire [4:0] \oc8051_golden_model_1.n1577 ;
  wire [4:0] \oc8051_golden_model_1.n1579 ;
  wire \oc8051_golden_model_1.n1580 ;
  wire \oc8051_golden_model_1.n1587 ;
  wire [7:0] \oc8051_golden_model_1.n1588 ;
  wire [6:0] \oc8051_golden_model_1.n1589 ;
  wire \oc8051_golden_model_1.n1604 ;
  wire [7:0] \oc8051_golden_model_1.n1605 ;
  wire [8:0] \oc8051_golden_model_1.n1609 ;
  wire \oc8051_golden_model_1.n1610 ;
  wire [4:0] \oc8051_golden_model_1.n1612 ;
  wire \oc8051_golden_model_1.n1613 ;
  wire \oc8051_golden_model_1.n1620 ;
  wire [7:0] \oc8051_golden_model_1.n1621 ;
  wire [6:0] \oc8051_golden_model_1.n1622 ;
  wire \oc8051_golden_model_1.n1637 ;
  wire [7:0] \oc8051_golden_model_1.n1638 ;
  wire [8:0] \oc8051_golden_model_1.n1642 ;
  wire \oc8051_golden_model_1.n1643 ;
  wire [4:0] \oc8051_golden_model_1.n1645 ;
  wire \oc8051_golden_model_1.n1646 ;
  wire \oc8051_golden_model_1.n1653 ;
  wire [7:0] \oc8051_golden_model_1.n1654 ;
  wire [6:0] \oc8051_golden_model_1.n1655 ;
  wire \oc8051_golden_model_1.n1670 ;
  wire [7:0] \oc8051_golden_model_1.n1671 ;
  wire [8:0] \oc8051_golden_model_1.n1675 ;
  wire \oc8051_golden_model_1.n1676 ;
  wire [4:0] \oc8051_golden_model_1.n1678 ;
  wire \oc8051_golden_model_1.n1679 ;
  wire \oc8051_golden_model_1.n1686 ;
  wire [7:0] \oc8051_golden_model_1.n1687 ;
  wire [6:0] \oc8051_golden_model_1.n1688 ;
  wire \oc8051_golden_model_1.n1703 ;
  wire [7:0] \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1730 ;
  wire [6:0] \oc8051_golden_model_1.n1731 ;
  wire [7:0] \oc8051_golden_model_1.n1732 ;
  wire \oc8051_golden_model_1.n1788 ;
  wire [7:0] \oc8051_golden_model_1.n1789 ;
  wire \oc8051_golden_model_1.n1805 ;
  wire [7:0] \oc8051_golden_model_1.n1806 ;
  wire \oc8051_golden_model_1.n1822 ;
  wire [7:0] \oc8051_golden_model_1.n1823 ;
  wire \oc8051_golden_model_1.n1839 ;
  wire [7:0] \oc8051_golden_model_1.n1840 ;
  wire [7:0] \oc8051_golden_model_1.n1864 ;
  wire [6:0] \oc8051_golden_model_1.n1865 ;
  wire [7:0] \oc8051_golden_model_1.n1866 ;
  wire \oc8051_golden_model_1.n1922 ;
  wire [7:0] \oc8051_golden_model_1.n1923 ;
  wire \oc8051_golden_model_1.n1939 ;
  wire [7:0] \oc8051_golden_model_1.n1940 ;
  wire \oc8051_golden_model_1.n1956 ;
  wire [7:0] \oc8051_golden_model_1.n1957 ;
  wire \oc8051_golden_model_1.n1973 ;
  wire [7:0] \oc8051_golden_model_1.n1974 ;
  wire \oc8051_golden_model_1.n2073 ;
  wire [7:0] \oc8051_golden_model_1.n2074 ;
  wire \oc8051_golden_model_1.n2090 ;
  wire [7:0] \oc8051_golden_model_1.n2091 ;
  wire \oc8051_golden_model_1.n2107 ;
  wire [7:0] \oc8051_golden_model_1.n2108 ;
  wire \oc8051_golden_model_1.n2124 ;
  wire [7:0] \oc8051_golden_model_1.n2125 ;
  wire \oc8051_golden_model_1.n2128 ;
  wire [6:0] \oc8051_golden_model_1.n2129 ;
  wire [7:0] \oc8051_golden_model_1.n2130 ;
  wire [6:0] \oc8051_golden_model_1.n2131 ;
  wire [7:0] \oc8051_golden_model_1.n2132 ;
  wire \oc8051_golden_model_1.n2147 ;
  wire [7:0] \oc8051_golden_model_1.n2148 ;
  wire \oc8051_golden_model_1.n2187 ;
  wire [7:0] \oc8051_golden_model_1.n2188 ;
  wire [6:0] \oc8051_golden_model_1.n2189 ;
  wire [7:0] \oc8051_golden_model_1.n2190 ;
  wire [3:0] \oc8051_golden_model_1.n2197 ;
  wire \oc8051_golden_model_1.n2198 ;
  wire [7:0] \oc8051_golden_model_1.n2199 ;
  wire [6:0] \oc8051_golden_model_1.n2200 ;
  wire \oc8051_golden_model_1.n2215 ;
  wire [7:0] \oc8051_golden_model_1.n2216 ;
  wire [7:0] \oc8051_golden_model_1.n2428 ;
  wire \oc8051_golden_model_1.n2431 ;
  wire \oc8051_golden_model_1.n2433 ;
  wire \oc8051_golden_model_1.n2439 ;
  wire [7:0] \oc8051_golden_model_1.n2440 ;
  wire [6:0] \oc8051_golden_model_1.n2441 ;
  wire \oc8051_golden_model_1.n2456 ;
  wire [7:0] \oc8051_golden_model_1.n2457 ;
  wire \oc8051_golden_model_1.n2461 ;
  wire \oc8051_golden_model_1.n2463 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire [6:0] \oc8051_golden_model_1.n2471 ;
  wire \oc8051_golden_model_1.n2486 ;
  wire [7:0] \oc8051_golden_model_1.n2487 ;
  wire \oc8051_golden_model_1.n2491 ;
  wire \oc8051_golden_model_1.n2493 ;
  wire \oc8051_golden_model_1.n2499 ;
  wire [7:0] \oc8051_golden_model_1.n2500 ;
  wire [6:0] \oc8051_golden_model_1.n2501 ;
  wire \oc8051_golden_model_1.n2516 ;
  wire [7:0] \oc8051_golden_model_1.n2517 ;
  wire \oc8051_golden_model_1.n2521 ;
  wire \oc8051_golden_model_1.n2523 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire [7:0] \oc8051_golden_model_1.n2530 ;
  wire [6:0] \oc8051_golden_model_1.n2531 ;
  wire \oc8051_golden_model_1.n2546 ;
  wire [7:0] \oc8051_golden_model_1.n2547 ;
  wire \oc8051_golden_model_1.n2549 ;
  wire [7:0] \oc8051_golden_model_1.n2550 ;
  wire [6:0] \oc8051_golden_model_1.n2551 ;
  wire [7:0] \oc8051_golden_model_1.n2552 ;
  wire [7:0] \oc8051_golden_model_1.n2553 ;
  wire [6:0] \oc8051_golden_model_1.n2554 ;
  wire [7:0] \oc8051_golden_model_1.n2555 ;
  wire [15:0] \oc8051_golden_model_1.n2559 ;
  wire \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [6:0] \oc8051_golden_model_1.n2567 ;
  wire \oc8051_golden_model_1.n2582 ;
  wire [7:0] \oc8051_golden_model_1.n2583 ;
  wire \oc8051_golden_model_1.n2586 ;
  wire [7:0] \oc8051_golden_model_1.n2587 ;
  wire [6:0] \oc8051_golden_model_1.n2588 ;
  wire [7:0] \oc8051_golden_model_1.n2589 ;
  wire \oc8051_golden_model_1.n2626 ;
  wire [7:0] \oc8051_golden_model_1.n2627 ;
  wire [6:0] \oc8051_golden_model_1.n2628 ;
  wire [7:0] \oc8051_golden_model_1.n2629 ;
  wire \oc8051_golden_model_1.n2634 ;
  wire [7:0] \oc8051_golden_model_1.n2635 ;
  wire [6:0] \oc8051_golden_model_1.n2636 ;
  wire [7:0] \oc8051_golden_model_1.n2637 ;
  wire \oc8051_golden_model_1.n2642 ;
  wire [7:0] \oc8051_golden_model_1.n2643 ;
  wire [6:0] \oc8051_golden_model_1.n2644 ;
  wire [7:0] \oc8051_golden_model_1.n2645 ;
  wire \oc8051_golden_model_1.n2650 ;
  wire [7:0] \oc8051_golden_model_1.n2651 ;
  wire [6:0] \oc8051_golden_model_1.n2652 ;
  wire [7:0] \oc8051_golden_model_1.n2653 ;
  wire \oc8051_golden_model_1.n2658 ;
  wire [7:0] \oc8051_golden_model_1.n2659 ;
  wire [6:0] \oc8051_golden_model_1.n2660 ;
  wire [7:0] \oc8051_golden_model_1.n2661 ;
  wire [7:0] \oc8051_golden_model_1.n2662 ;
  wire [6:0] \oc8051_golden_model_1.n2663 ;
  wire [7:0] \oc8051_golden_model_1.n2664 ;
  wire [3:0] \oc8051_golden_model_1.n2665 ;
  wire [7:0] \oc8051_golden_model_1.n2666 ;
  wire \oc8051_golden_model_1.n2667 ;
  wire \oc8051_golden_model_1.n2668 ;
  wire \oc8051_golden_model_1.n2669 ;
  wire \oc8051_golden_model_1.n2670 ;
  wire \oc8051_golden_model_1.n2671 ;
  wire \oc8051_golden_model_1.n2672 ;
  wire \oc8051_golden_model_1.n2673 ;
  wire \oc8051_golden_model_1.n2674 ;
  wire \oc8051_golden_model_1.n2681 ;
  wire [7:0] \oc8051_golden_model_1.n2682 ;
  wire [7:0] \oc8051_golden_model_1.n2702 ;
  wire [6:0] \oc8051_golden_model_1.n2703 ;
  wire [7:0] \oc8051_golden_model_1.n2719 ;
  wire \oc8051_golden_model_1.n2720 ;
  wire \oc8051_golden_model_1.n2721 ;
  wire \oc8051_golden_model_1.n2722 ;
  wire \oc8051_golden_model_1.n2723 ;
  wire \oc8051_golden_model_1.n2724 ;
  wire \oc8051_golden_model_1.n2725 ;
  wire \oc8051_golden_model_1.n2726 ;
  wire \oc8051_golden_model_1.n2727 ;
  wire \oc8051_golden_model_1.n2734 ;
  wire [7:0] \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2736 ;
  wire \oc8051_golden_model_1.n2737 ;
  wire \oc8051_golden_model_1.n2738 ;
  wire \oc8051_golden_model_1.n2739 ;
  wire \oc8051_golden_model_1.n2740 ;
  wire \oc8051_golden_model_1.n2741 ;
  wire \oc8051_golden_model_1.n2742 ;
  wire \oc8051_golden_model_1.n2743 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire [7:0] \oc8051_golden_model_1.n2751 ;
  wire [7:0] \oc8051_golden_model_1.n2784 ;
  wire [6:0] \oc8051_golden_model_1.n2785 ;
  wire [7:0] \oc8051_golden_model_1.n2786 ;
  wire \oc8051_golden_model_1.n2805 ;
  wire [7:0] \oc8051_golden_model_1.n2806 ;
  wire [6:0] \oc8051_golden_model_1.n2807 ;
  wire \oc8051_golden_model_1.n2822 ;
  wire [7:0] \oc8051_golden_model_1.n2823 ;
  wire [7:0] \oc8051_golden_model_1.n2827 ;
  wire [3:0] \oc8051_golden_model_1.n2828 ;
  wire [7:0] \oc8051_golden_model_1.n2829 ;
  wire \oc8051_golden_model_1.n2830 ;
  wire \oc8051_golden_model_1.n2831 ;
  wire \oc8051_golden_model_1.n2832 ;
  wire \oc8051_golden_model_1.n2833 ;
  wire \oc8051_golden_model_1.n2834 ;
  wire \oc8051_golden_model_1.n2835 ;
  wire \oc8051_golden_model_1.n2836 ;
  wire \oc8051_golden_model_1.n2837 ;
  wire \oc8051_golden_model_1.n2844 ;
  wire [7:0] \oc8051_golden_model_1.n2845 ;
  wire \oc8051_golden_model_1.n2863 ;
  wire [7:0] \oc8051_golden_model_1.n2864 ;
  wire \oc8051_golden_model_1.n2880 ;
  wire [7:0] \oc8051_golden_model_1.n2881 ;
  wire [7:0] \oc8051_golden_model_1.n2882 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff0 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff1 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff2 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff3 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_41894_, rst);
  not (_16086_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_16097_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_16108_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _16097_);
  and (_16119_, _16108_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_16130_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _16097_);
  and (_16141_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _16097_);
  nor (_16151_, _16141_, _16130_);
  and (_16162_, _16151_, _16119_);
  nor (_16173_, _16162_, _16086_);
  and (_16184_, _16086_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_16195_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_16206_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _16195_);
  nor (_16217_, _16206_, _16184_);
  not (_16228_, _16217_);
  and (_16239_, _16228_, _16162_);
  or (_16250_, _16239_, _16173_);
  and (_22329_, _16250_, _41894_);
  nor (_16271_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_16282_, _16271_);
  and (_16293_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_16304_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_16315_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_16326_, _16315_);
  not (_16337_, _16206_);
  nor (_16348_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_16359_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_16370_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _16359_);
  nor (_16381_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_16392_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_16403_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _16392_);
  nor (_16414_, _16403_, _16381_);
  nor (_16425_, _16414_, _16370_);
  not (_16436_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_16458_, _16370_, _16436_);
  nor (_16459_, _16458_, _16425_);
  and (_16470_, _16459_, _16348_);
  not (_16480_, _16470_);
  and (_16491_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16502_, _16491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_16513_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16524_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _16513_);
  and (_16535_, _16524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_16546_, _16535_, _16502_);
  and (_16557_, _16546_, _16480_);
  nor (_16568_, _16557_, _16337_);
  not (_16579_, _16184_);
  nor (_16590_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_16601_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _16392_);
  nor (_16612_, _16601_, _16590_);
  nor (_16623_, _16612_, _16370_);
  not (_16634_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_16645_, _16370_, _16634_);
  nor (_16656_, _16645_, _16623_);
  and (_16667_, _16656_, _16348_);
  not (_16678_, _16667_);
  and (_16689_, _16491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_16700_, _16524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_16711_, _16700_, _16689_);
  and (_16722_, _16711_, _16678_);
  nor (_16733_, _16722_, _16579_);
  nor (_16744_, _16733_, _16568_);
  nor (_16755_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_16766_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _16392_);
  nor (_16777_, _16766_, _16755_);
  nor (_16788_, _16777_, _16370_);
  not (_16799_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_16810_, _16370_, _16799_);
  nor (_16821_, _16810_, _16788_);
  and (_16831_, _16821_, _16348_);
  not (_16842_, _16831_);
  and (_16853_, _16491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_16864_, _16524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_16875_, _16864_, _16853_);
  and (_16886_, _16875_, _16842_);
  nor (_16897_, _16886_, _16228_);
  nor (_16908_, _16897_, _16271_);
  and (_16919_, _16908_, _16744_);
  nor (_16930_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_16941_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _16392_);
  nor (_16952_, _16941_, _16930_);
  nor (_16963_, _16952_, _16370_);
  not (_16974_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_16985_, _16370_, _16974_);
  nor (_16996_, _16985_, _16963_);
  and (_17007_, _16996_, _16348_);
  not (_17018_, _17007_);
  and (_17029_, _16491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_17040_, _16524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_17051_, _17040_, _17029_);
  and (_17062_, _17051_, _17018_);
  and (_17073_, _17062_, _16271_);
  nor (_17084_, _17073_, _16919_);
  not (_17095_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_17106_, _17095_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_17117_, _17106_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17128_, _17117_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_17139_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_17150_, _17139_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17160_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_17181_, _17160_, _17128_);
  not (_17182_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17203_, _17106_, _17182_);
  and (_17204_, _17203_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_17215_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17226_, _17215_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_17237_, _17226_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_17247_, _17237_, _17204_);
  and (_17258_, _17247_, _17181_);
  and (_17269_, _17139_, _17182_);
  and (_17280_, _17269_, _16996_);
  and (_17291_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_17302_, _17291_, _17182_);
  and (_17313_, _17302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_17324_, _17291_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_17334_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_17345_, _17334_, _17313_);
  not (_17356_, _17345_);
  nor (_17367_, _17356_, _17280_);
  and (_17378_, _17367_, _17258_);
  not (_17389_, _17378_);
  and (_17400_, _17389_, _17084_);
  not (_17411_, _17400_);
  nor (_17421_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_17432_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _16392_);
  nor (_17443_, _17432_, _17421_);
  nor (_17454_, _17443_, _16370_);
  not (_17465_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_17476_, _16370_, _17465_);
  nor (_17487_, _17476_, _17454_);
  and (_17498_, _17487_, _16348_);
  not (_17508_, _17498_);
  and (_17519_, _16491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_17530_, _16524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_17541_, _17530_, _17519_);
  and (_17552_, _17541_, _17508_);
  nor (_17563_, _17552_, _16337_);
  nor (_17574_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_17585_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _16392_);
  nor (_17595_, _17585_, _17574_);
  nor (_17606_, _17595_, _16370_);
  not (_17617_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_17628_, _16370_, _17617_);
  nor (_17639_, _17628_, _17606_);
  and (_17650_, _17639_, _16348_);
  not (_17661_, _17650_);
  and (_17672_, _16491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_17682_, _16524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17693_, _17682_, _17672_);
  and (_17704_, _17693_, _17661_);
  nor (_17715_, _17704_, _16579_);
  nor (_17726_, _17715_, _17563_);
  nor (_17737_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_17748_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _16392_);
  nor (_17759_, _17748_, _17737_);
  nor (_17769_, _17759_, _16370_);
  not (_17780_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_17791_, _16370_, _17780_);
  nor (_17802_, _17791_, _17769_);
  and (_17813_, _17802_, _16348_);
  not (_17824_, _17813_);
  and (_17835_, _16491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_17846_, _16524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_17857_, _17846_, _17835_);
  and (_17868_, _17857_, _17824_);
  nor (_17878_, _17868_, _16228_);
  nor (_17889_, _17878_, _16271_);
  and (_17900_, _17889_, _17726_);
  nor (_17911_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_17922_, _16392_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_17933_, _17922_, _17911_);
  nor (_17944_, _17933_, _16370_);
  not (_17955_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_17966_, _16370_, _17955_);
  nor (_17977_, _17966_, _17944_);
  and (_17987_, _17977_, _16348_);
  not (_17998_, _17987_);
  and (_18009_, _16491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_18020_, _16524_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_18031_, _18020_, _18009_);
  and (_18042_, _18031_, _17998_);
  and (_18053_, _18042_, _16271_);
  or (_18064_, _18053_, _17900_);
  and (_18075_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_18086_, _17117_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_18097_, _18086_, _18075_);
  and (_18107_, _17302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_18118_, _17226_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_18129_, _18118_, _18107_);
  and (_18140_, _18129_, _18097_);
  and (_18151_, _17977_, _17269_);
  and (_18162_, _17203_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_18173_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_18184_, _18173_, _18162_);
  not (_18195_, _18184_);
  nor (_18206_, _18195_, _18151_);
  and (_18216_, _18206_, _18140_);
  nor (_18227_, _18216_, _18064_);
  and (_18238_, _18227_, _17411_);
  not (_18249_, _18238_);
  and (_18260_, _17117_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_18271_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_18282_, _18271_, _18260_);
  and (_18293_, _17226_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_18304_, _17203_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_18315_, _18304_, _18293_);
  and (_18326_, _18315_, _18282_);
  and (_18336_, _17639_, _17269_);
  and (_18347_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_18358_, _17302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_18369_, _18358_, _18347_);
  not (_18380_, _18369_);
  nor (_18391_, _18380_, _18336_);
  and (_18402_, _18391_, _18326_);
  nor (_18413_, _18402_, _18064_);
  and (_18424_, _17117_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_18435_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_18445_, _18435_, _18424_);
  and (_18456_, _17226_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_18467_, _17203_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_18478_, _18467_, _18456_);
  and (_18489_, _18478_, _18445_);
  and (_18500_, _17269_, _16656_);
  and (_18511_, _17302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_18522_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_18533_, _18522_, _18511_);
  not (_18544_, _18533_);
  nor (_18555_, _18544_, _18500_);
  and (_18565_, _18555_, _18489_);
  not (_18576_, _18565_);
  and (_18587_, _18576_, _17084_);
  and (_18598_, _18413_, _18587_);
  and (_18609_, _17389_, _18598_);
  nor (_18620_, _17400_, _18598_);
  nor (_18631_, _18620_, _18609_);
  and (_18641_, _18631_, _18413_);
  and (_18652_, _18227_, _17400_);
  nor (_18663_, _17378_, _18064_);
  not (_18674_, _18216_);
  and (_18685_, _18674_, _17084_);
  nor (_18696_, _18685_, _18663_);
  nor (_18707_, _18696_, _18652_);
  and (_18718_, _18707_, _18641_);
  nor (_18729_, _18707_, _18641_);
  nor (_18739_, _18729_, _18718_);
  and (_18750_, _18739_, _18609_);
  nor (_18761_, _18750_, _18718_);
  nor (_18772_, _18761_, _18249_);
  nor (_18783_, _18064_, _18565_);
  and (_18794_, _17117_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_18805_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_18816_, _18805_, _18794_);
  and (_18826_, _17226_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_18837_, _17203_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_18848_, _18837_, _18826_);
  and (_18859_, _18848_, _18816_);
  and (_18870_, _17487_, _17269_);
  and (_18881_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_18892_, _17302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_18903_, _18892_, _18881_);
  not (_18913_, _18903_);
  nor (_18924_, _18913_, _18870_);
  and (_18935_, _18924_, _18859_);
  not (_18946_, _18935_);
  and (_18957_, _18946_, _17084_);
  and (_18968_, _18957_, _18783_);
  not (_18979_, _18402_);
  and (_18990_, _18979_, _17084_);
  nor (_19000_, _18990_, _18783_);
  nor (_19011_, _19000_, _18598_);
  and (_19022_, _19011_, _18968_);
  nor (_19033_, _17400_, _18413_);
  nor (_19044_, _19033_, _18641_);
  and (_19055_, _19044_, _19022_);
  nor (_19066_, _18739_, _18609_);
  nor (_19077_, _19066_, _18750_);
  and (_19087_, _19077_, _19055_);
  nor (_19098_, _19077_, _19055_);
  nor (_19109_, _19098_, _19087_);
  not (_19120_, _19109_);
  and (_19131_, _17117_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_19142_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_19153_, _19142_, _19131_);
  and (_19164_, _17226_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_19174_, _17203_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_19185_, _19174_, _19164_);
  and (_19196_, _19185_, _19153_);
  and (_19207_, _17802_, _17269_);
  and (_19218_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_19229_, _17302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_19240_, _19229_, _19218_);
  not (_19251_, _19240_);
  nor (_19262_, _19251_, _19207_);
  and (_19272_, _19262_, _19196_);
  nor (_19283_, _19272_, _18064_);
  and (_19294_, _17117_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_19305_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_19316_, _19305_, _19294_);
  and (_19327_, _17226_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_19338_, _17203_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_19349_, _19338_, _19327_);
  and (_19360_, _19349_, _19316_);
  and (_19371_, _17269_, _16459_);
  and (_19382_, _17302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_19392_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_19403_, _19392_, _19382_);
  not (_19414_, _19403_);
  nor (_19425_, _19414_, _19371_);
  and (_19436_, _19425_, _19360_);
  not (_19447_, _19436_);
  and (_19458_, _19447_, _17084_);
  and (_19469_, _19458_, _19283_);
  not (_19480_, _19272_);
  and (_19491_, _19480_, _17084_);
  not (_19501_, _19491_);
  nor (_19512_, _19436_, _18064_);
  and (_19523_, _19512_, _19501_);
  and (_19534_, _19523_, _18957_);
  nor (_19545_, _19534_, _19469_);
  nor (_19556_, _18935_, _18064_);
  nor (_19567_, _19556_, _18587_);
  nor (_19578_, _19567_, _18968_);
  not (_19589_, _19578_);
  nor (_19600_, _19589_, _19545_);
  nor (_19611_, _19011_, _18968_);
  nor (_19621_, _19611_, _19022_);
  and (_19632_, _19621_, _19600_);
  nor (_19643_, _19044_, _19022_);
  nor (_19654_, _19643_, _19055_);
  and (_19665_, _19654_, _19632_);
  and (_19676_, _17117_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_19687_, _17150_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_19698_, _19687_, _19676_);
  and (_19709_, _17226_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_19720_, _17203_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_19730_, _19720_, _19709_);
  and (_19741_, _19730_, _19698_);
  and (_19752_, _17269_, _16821_);
  and (_19763_, _17324_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_19774_, _17302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_19785_, _19774_, _19763_);
  not (_19796_, _19785_);
  nor (_19807_, _19796_, _19752_);
  and (_19818_, _19807_, _19741_);
  nor (_19829_, _19818_, _18064_);
  and (_19839_, _19829_, _19491_);
  nor (_19850_, _19458_, _19283_);
  nor (_19861_, _19850_, _19469_);
  and (_19872_, _19861_, _19839_);
  nor (_19883_, _19523_, _18957_);
  nor (_19894_, _19883_, _19534_);
  and (_19905_, _19894_, _19872_);
  and (_19916_, _19589_, _19545_);
  nor (_19927_, _19916_, _19600_);
  and (_19938_, _19927_, _19905_);
  nor (_19949_, _19621_, _19600_);
  nor (_19959_, _19949_, _19632_);
  and (_19970_, _19959_, _19938_);
  nor (_19981_, _19654_, _19632_);
  nor (_19992_, _19981_, _19665_);
  and (_20003_, _19992_, _19970_);
  nor (_20014_, _20003_, _19665_);
  nor (_20025_, _20014_, _19120_);
  nor (_20036_, _20025_, _19087_);
  and (_20046_, _18761_, _18249_);
  nor (_20057_, _20046_, _18772_);
  not (_20068_, _20057_);
  nor (_20079_, _20068_, _20036_);
  or (_20090_, _20079_, _18652_);
  nor (_20101_, _20090_, _18772_);
  nor (_20112_, _20101_, _16326_);
  and (_20123_, _20101_, _16326_);
  nor (_20133_, _20123_, _20112_);
  not (_20144_, _20133_);
  and (_20155_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_20166_, _20068_, _20036_);
  nor (_20177_, _20166_, _20079_);
  and (_20188_, _20177_, _20155_);
  and (_20199_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_20210_, _20014_, _19120_);
  nor (_20220_, _20210_, _20025_);
  and (_20231_, _20220_, _20199_);
  nor (_20242_, _20220_, _20199_);
  nor (_20253_, _20242_, _20231_);
  not (_20264_, _20253_);
  and (_20275_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_20286_, _19992_, _19970_);
  nor (_20297_, _20286_, _20003_);
  and (_20307_, _20297_, _20275_);
  nor (_20318_, _20297_, _20275_);
  nor (_20329_, _20318_, _20307_);
  not (_20340_, _20329_);
  and (_20351_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_20362_, _19959_, _19938_);
  nor (_20373_, _20362_, _19970_);
  and (_20384_, _20373_, _20351_);
  nor (_20394_, _20373_, _20351_);
  nor (_20405_, _20394_, _20384_);
  not (_20416_, _20405_);
  and (_20427_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_20438_, _19927_, _19905_);
  nor (_20449_, _20438_, _19938_);
  and (_20460_, _20449_, _20427_);
  and (_20471_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_20481_, _19894_, _19872_);
  nor (_20492_, _20481_, _19905_);
  and (_20503_, _20492_, _20471_);
  and (_20514_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_20525_, _19861_, _19839_);
  nor (_20536_, _20525_, _19872_);
  and (_20547_, _20536_, _20514_);
  nor (_20558_, _20492_, _20471_);
  nor (_20568_, _20558_, _20503_);
  and (_20579_, _20568_, _20547_);
  nor (_20590_, _20579_, _20503_);
  not (_20601_, _20590_);
  nor (_20612_, _20449_, _20427_);
  nor (_20623_, _20612_, _20460_);
  and (_20634_, _20623_, _20601_);
  nor (_20644_, _20634_, _20460_);
  nor (_20655_, _20644_, _20416_);
  nor (_20666_, _20655_, _20384_);
  nor (_20677_, _20666_, _20340_);
  nor (_20688_, _20677_, _20307_);
  nor (_20699_, _20688_, _20264_);
  nor (_20710_, _20699_, _20231_);
  nor (_20721_, _20177_, _20155_);
  nor (_20731_, _20721_, _20188_);
  not (_20742_, _20731_);
  nor (_20753_, _20742_, _20710_);
  nor (_20764_, _20753_, _20188_);
  nor (_20775_, _20764_, _20144_);
  nor (_20786_, _20775_, _20112_);
  not (_20797_, _20786_);
  and (_20808_, _20797_, _16304_);
  and (_20818_, _20808_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_20829_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_20840_, _20829_, _20818_);
  and (_20851_, _20840_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_20862_, _20851_, _16293_);
  and (_20873_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20884_, _20873_, _20862_);
  and (_20895_, _20862_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20905_, _20895_, _20884_);
  and (_24502_, _20905_, _41894_);
  nor (_20926_, _16162_, _16195_);
  and (_20937_, _16162_, _16195_);
  or (_20948_, _20937_, _20926_);
  and (_02425_, _20948_, _41894_);
  not (_20969_, _19818_);
  and (_20980_, _20969_, _17084_);
  and (_02620_, _20980_, _41894_);
  nor (_21000_, _19829_, _19491_);
  nor (_21011_, _21000_, _19839_);
  and (_02814_, _21011_, _41894_);
  nor (_21032_, _20536_, _20514_);
  nor (_21043_, _21032_, _20547_);
  and (_03012_, _21043_, _41894_);
  nor (_21064_, _20568_, _20547_);
  nor (_21074_, _21064_, _20579_);
  and (_03220_, _21074_, _41894_);
  nor (_21095_, _20623_, _20601_);
  nor (_21106_, _21095_, _20634_);
  and (_03421_, _21106_, _41894_);
  and (_21127_, _20644_, _20416_);
  nor (_21138_, _21127_, _20655_);
  and (_03622_, _21138_, _41894_);
  and (_21158_, _20666_, _20340_);
  nor (_21169_, _21158_, _20677_);
  and (_03823_, _21169_, _41894_);
  and (_21190_, _20688_, _20264_);
  nor (_21201_, _21190_, _20699_);
  and (_04024_, _21201_, _41894_);
  and (_21222_, _20742_, _20710_);
  nor (_21232_, _21222_, _20753_);
  and (_04125_, _21232_, _41894_);
  and (_21253_, _20764_, _20144_);
  nor (_21264_, _21253_, _20775_);
  and (_04226_, _21264_, _41894_);
  nor (_21285_, _20797_, _16304_);
  nor (_21296_, _21285_, _20808_);
  and (_04327_, _21296_, _41894_);
  and (_21316_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_21327_, _21316_, _20808_);
  nor (_21338_, _21327_, _20818_);
  and (_04428_, _21338_, _41894_);
  nor (_21359_, _20829_, _20818_);
  nor (_21370_, _21359_, _20840_);
  and (_04529_, _21370_, _41894_);
  and (_21403_, _16282_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_21414_, _21403_, _20840_);
  nor (_21426_, _21414_, _20851_);
  and (_04630_, _21426_, _41894_);
  nor (_21449_, _20851_, _16293_);
  nor (_21450_, _21449_, _20862_);
  and (_04731_, _21450_, _41894_);
  and (_21471_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _16097_);
  nor (_21482_, _21471_, _16108_);
  not (_21493_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_21503_, _16130_, _21493_);
  and (_21514_, _21503_, _21482_);
  and (_21525_, _21514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_21536_, _21525_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21547_, _21525_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21558_, _21547_, _21536_);
  and (_00839_, _21558_, _41894_);
  and (_00864_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _41894_);
  not (_21588_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_21599_, _17868_, _21588_);
  and (_21610_, _17552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21621_, _21610_, _21599_);
  nor (_21632_, _21621_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21643_, _17704_, _21588_);
  and (_21654_, _18042_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_21665_, _21654_, _21643_);
  and (_21675_, _21665_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21686_, _21675_, _21632_);
  nor (_21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_21708_, _21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and (_21719_, _21697_, _18216_);
  nor (_21730_, _21719_, _21708_);
  not (_21741_, _21730_);
  and (_21752_, _16886_, _21588_);
  and (_21762_, _16557_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21773_, _21762_, _21752_);
  nor (_21784_, _21773_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21795_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21806_, _16722_, _21588_);
  and (_21817_, _17062_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21828_, _21817_, _21806_);
  nor (_21838_, _21828_, _21795_);
  nor (_21849_, _21838_, _21784_);
  nor (_21860_, _21849_, _21741_);
  and (_21871_, _21849_, _21741_);
  nor (_21882_, _21871_, _21860_);
  and (_21893_, _21697_, _17378_);
  nor (_21904_, _21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor (_21915_, _21904_, _21893_);
  not (_21926_, _21915_);
  nor (_21936_, _17868_, _21588_);
  nor (_21957_, _21936_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21958_, _17552_, _21588_);
  and (_21969_, _17704_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21980_, _21969_, _21958_);
  nor (_21991_, _21980_, _21795_);
  nor (_22002_, _21991_, _21957_);
  nor (_22013_, _22002_, _21926_);
  and (_22023_, _22002_, _21926_);
  nor (_22034_, _22023_, _22013_);
  not (_22045_, _22034_);
  nor (_22056_, _21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_22067_, _21697_, _18402_);
  nor (_22078_, _22067_, _22056_);
  not (_22089_, _22078_);
  nor (_22100_, _16886_, _21588_);
  nor (_22110_, _22100_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_22121_, _16557_, _21588_);
  and (_22132_, _16722_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_22143_, _22132_, _22121_);
  nor (_22154_, _22143_, _21795_);
  nor (_22165_, _22154_, _22110_);
  nor (_22176_, _22165_, _22089_);
  and (_22187_, _22165_, _22089_);
  and (_22197_, _21621_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22219_, _22197_);
  nor (_22220_, _21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_22231_, _21697_, _18565_);
  nor (_22242_, _22231_, _22220_);
  and (_22253_, _22242_, _22219_);
  and (_22264_, _21773_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22275_, _22264_);
  and (_22285_, _21697_, _18935_);
  nor (_22296_, _21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_22307_, _22296_, _22285_);
  and (_22318_, _22307_, _22275_);
  nor (_22330_, _22307_, _22275_);
  nor (_22341_, _22330_, _22318_);
  not (_22352_, _22341_);
  and (_22363_, _21936_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22373_, _22363_);
  and (_22384_, _21697_, _19436_);
  nor (_22395_, _21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_22406_, _22395_, _22384_);
  and (_22417_, _22406_, _22373_);
  and (_22428_, _22100_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22439_, _22428_);
  and (_22449_, _21697_, _19272_);
  nor (_22460_, _21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  nor (_22471_, _22460_, _22449_);
  nor (_22482_, _22471_, _22439_);
  not (_22493_, _22482_);
  nor (_22504_, _22406_, _22373_);
  nor (_22515_, _22504_, _22417_);
  and (_22526_, _22515_, _22493_);
  nor (_22537_, _22526_, _22417_);
  nor (_22547_, _22537_, _22352_);
  nor (_22558_, _22547_, _22318_);
  nor (_22569_, _22242_, _22219_);
  nor (_22580_, _22569_, _22253_);
  not (_22591_, _22580_);
  nor (_22602_, _22591_, _22558_);
  nor (_22613_, _22602_, _22253_);
  nor (_22624_, _22613_, _22187_);
  nor (_22634_, _22624_, _22176_);
  nor (_22645_, _22634_, _22045_);
  nor (_22656_, _22645_, _22013_);
  not (_22667_, _22656_);
  and (_22678_, _22667_, _21882_);
  or (_22689_, _22678_, _21860_);
  and (_22700_, _18042_, _17062_);
  or (_22711_, _22700_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_22721_, _21828_);
  and (_22732_, _21665_, _22721_);
  nor (_22743_, _22143_, _21980_);
  and (_22754_, _22743_, _22732_);
  or (_22765_, _22754_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_22776_, _22765_, _22711_);
  and (_22787_, _22776_, _22689_);
  and (_22798_, _22787_, _21686_);
  nor (_22808_, _22667_, _21882_);
  or (_22819_, _22808_, _22678_);
  and (_22830_, _22819_, _22798_);
  nor (_22841_, _22798_, _21730_);
  nor (_22852_, _22841_, _22830_);
  not (_22863_, _22852_);
  and (_22874_, _22852_, _21686_);
  not (_22894_, _21849_);
  nor (_22895_, _22798_, _21926_);
  and (_22906_, _22634_, _22045_);
  nor (_22927_, _22906_, _22645_);
  and (_22928_, _22927_, _22798_);
  or (_22939_, _22928_, _22895_);
  and (_22960_, _22939_, _22894_);
  nor (_22961_, _22939_, _22894_);
  nor (_22972_, _22961_, _22960_);
  not (_22992_, _22972_);
  not (_22993_, _22002_);
  nor (_23004_, _22798_, _22089_);
  nor (_23025_, _22187_, _22176_);
  nor (_23026_, _23025_, _22613_);
  and (_23037_, _23025_, _22613_);
  or (_23058_, _23037_, _23026_);
  and (_23059_, _23058_, _22798_);
  or (_23070_, _23059_, _23004_);
  and (_23090_, _23070_, _22993_);
  nor (_23091_, _23070_, _22993_);
  not (_23102_, _22165_);
  and (_23113_, _22591_, _22558_);
  or (_23124_, _23113_, _22602_);
  and (_23135_, _23124_, _22798_);
  nor (_23146_, _22798_, _22242_);
  nor (_23157_, _23146_, _23135_);
  and (_23168_, _23157_, _23102_);
  and (_23179_, _22537_, _22352_);
  nor (_23190_, _23179_, _22547_);
  not (_23200_, _23190_);
  and (_23211_, _23200_, _22798_);
  nor (_23222_, _22798_, _22307_);
  nor (_23233_, _23222_, _23211_);
  and (_23244_, _23233_, _22219_);
  nor (_23255_, _23233_, _22219_);
  nor (_23266_, _23255_, _23244_);
  not (_23277_, _23266_);
  nor (_23288_, _22515_, _22493_);
  nor (_23299_, _23288_, _22526_);
  not (_23309_, _23299_);
  and (_23320_, _23309_, _22798_);
  nor (_23331_, _22798_, _22406_);
  nor (_23342_, _23331_, _23320_);
  and (_23353_, _23342_, _22275_);
  not (_23364_, _22471_);
  and (_23375_, _22798_, _22428_);
  or (_23386_, _23375_, _23364_);
  nand (_23397_, _22798_, _22428_);
  or (_23408_, _23397_, _22471_);
  and (_23419_, _23408_, _23386_);
  nor (_23429_, _23419_, _22363_);
  and (_23440_, _23419_, _22363_);
  nor (_23451_, _23440_, _23429_);
  and (_23462_, _21697_, _19818_);
  nor (_23473_, _21697_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_23484_, _23473_, _23462_);
  nor (_23495_, _23484_, _22439_);
  not (_23506_, _23495_);
  and (_23517_, _23506_, _23451_);
  nor (_23528_, _23517_, _23429_);
  nor (_23538_, _23342_, _22275_);
  nor (_23549_, _23538_, _23353_);
  not (_23560_, _23549_);
  nor (_23571_, _23560_, _23528_);
  nor (_23582_, _23571_, _23353_);
  nor (_23593_, _23582_, _23277_);
  nor (_23604_, _23593_, _23244_);
  nor (_23615_, _23157_, _23102_);
  nor (_23626_, _23615_, _23168_);
  not (_23637_, _23626_);
  nor (_23648_, _23637_, _23604_);
  nor (_23658_, _23648_, _23168_);
  nor (_23669_, _23658_, _23091_);
  nor (_23680_, _23669_, _23090_);
  nor (_23691_, _23680_, _22992_);
  or (_23702_, _23691_, _22960_);
  or (_23713_, _23702_, _22874_);
  and (_23724_, _23713_, _22776_);
  nor (_23735_, _23724_, _22863_);
  and (_23746_, _22874_, _22776_);
  and (_23757_, _23746_, _23702_);
  or (_23767_, _23757_, _23735_);
  and (_00882_, _23767_, _41894_);
  or (_23788_, _22852_, _21686_);
  and (_23799_, _23788_, _23724_);
  and (_02970_, _23799_, _41894_);
  and (_02981_, _22798_, _41894_);
  and (_03001_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _41894_);
  and (_03022_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _41894_);
  and (_03043_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _41894_);
  or (_23860_, _21514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23870_, _21525_, rst);
  and (_03053_, _23870_, _23860_);
  and (_23891_, _23799_, _22428_);
  or (_23902_, _23891_, _23484_);
  nand (_23913_, _23891_, _23484_);
  and (_23924_, _23913_, _23902_);
  and (_03064_, _23924_, _41894_);
  nor (_23945_, _23799_, _23419_);
  nor (_23956_, _23506_, _23451_);
  nor (_23967_, _23956_, _23517_);
  and (_23977_, _23967_, _23799_);
  or (_23988_, _23977_, _23945_);
  and (_03075_, _23988_, _41894_);
  and (_24009_, _23560_, _23528_);
  or (_24020_, _24009_, _23571_);
  nand (_24031_, _24020_, _23799_);
  or (_24042_, _23799_, _23342_);
  and (_24053_, _24042_, _24031_);
  and (_03085_, _24053_, _41894_);
  and (_24086_, _23582_, _23277_);
  or (_24097_, _24086_, _23593_);
  nand (_24109_, _24097_, _23799_);
  or (_24121_, _23799_, _23233_);
  and (_24133_, _24121_, _24109_);
  and (_03096_, _24133_, _41894_);
  and (_24145_, _23637_, _23604_);
  or (_24156_, _24145_, _23648_);
  nand (_24167_, _24156_, _23799_);
  or (_24178_, _23799_, _23157_);
  and (_24189_, _24178_, _24167_);
  and (_03107_, _24189_, _41894_);
  or (_24209_, _23091_, _23090_);
  and (_24220_, _24209_, _23658_);
  nor (_24231_, _24209_, _23658_);
  or (_24242_, _24231_, _24220_);
  nand (_24253_, _24242_, _23799_);
  or (_24264_, _23799_, _23070_);
  and (_24275_, _24264_, _24253_);
  and (_03118_, _24275_, _41894_);
  and (_24296_, _23680_, _22992_);
  or (_24307_, _24296_, _23691_);
  nand (_24317_, _24307_, _23799_);
  or (_24328_, _23799_, _22939_);
  and (_24339_, _24328_, _24317_);
  and (_03129_, _24339_, _41894_);
  not (_24360_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24371_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _16097_);
  and (_24382_, _24371_, _24360_);
  and (_24393_, _24382_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_24404_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24415_, _24404_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24426_, _24404_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24436_, _24426_, _24415_);
  and (_24447_, _24436_, _24393_);
  not (_24458_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_24469_, _24382_, _24458_);
  and (_24480_, _24469_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24491_, _24480_, _24447_);
  not (_24503_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_24514_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _16097_);
  and (_24525_, _24514_, _24503_);
  and (_24536_, _24525_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24546_, _24536_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_24557_, _24525_, _24360_);
  and (_24568_, _24557_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_24579_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24590_, _24579_, _16097_);
  nor (_24601_, _24590_, _24514_);
  and (_24612_, _24601_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_24623_, _24612_, _24568_);
  nor (_24633_, _24623_, _24546_);
  and (_24644_, _24633_, _24491_);
  and (_24655_, _24536_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_24666_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24677_, _24666_, _24404_);
  and (_24688_, _24677_, _24393_);
  nor (_24699_, _24688_, _24655_);
  and (_24710_, _24469_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_24721_, _24601_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_24731_, _24557_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_24742_, _24731_, _24721_);
  nor (_24753_, _24742_, _24710_);
  and (_24764_, _24753_, _24699_);
  and (_24775_, _24536_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_24786_, _24601_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_24797_, _24786_, _24775_);
  not (_24808_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24818_, _24393_, _24808_);
  not (_24829_, _24818_);
  and (_24840_, _24557_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_24851_, _24469_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_24862_, _24851_, _24840_);
  and (_24873_, _24862_, _24829_);
  and (_24884_, _24873_, _24797_);
  and (_24895_, _24884_, _24764_);
  and (_24906_, _24895_, _24644_);
  and (_24916_, _24415_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_24927_, _24916_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_24938_, _24927_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_24949_, _24938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_24960_, _24949_);
  not (_24971_, _24393_);
  nor (_24992_, _24938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_24993_, _24992_, _24971_);
  and (_25003_, _24993_, _24960_);
  not (_25014_, _25003_);
  and (_25035_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_25036_, _25035_, _24371_);
  and (_25047_, _24557_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_25068_, _25047_, _25036_);
  and (_25069_, _24469_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_25080_, _24536_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_25091_, _25080_, _25069_);
  and (_25101_, _25091_, _25068_);
  and (_25122_, _25101_, _25014_);
  nor (_25123_, _24927_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_25134_, _25123_);
  nor (_25145_, _24938_, _24971_);
  and (_25156_, _25145_, _25134_);
  not (_25167_, _25156_);
  and (_25178_, _24557_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_25188_, _25178_, _25036_);
  and (_25199_, _24469_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_25210_, _24536_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_25221_, _25210_, _25199_);
  and (_25232_, _25221_, _25188_);
  and (_25253_, _25232_, _25167_);
  nor (_25254_, _25253_, _25122_);
  not (_25265_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_25275_, _24949_, _25265_);
  and (_25286_, _24949_, _25265_);
  nor (_25297_, _25286_, _25275_);
  nor (_25308_, _25297_, _24971_);
  not (_25319_, _25308_);
  and (_25330_, _24557_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_25341_, _25330_, _25036_);
  and (_25352_, _24469_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_25363_, _24536_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_25373_, _25363_, _25352_);
  and (_25384_, _25373_, _25341_);
  and (_25395_, _25384_, _25319_);
  not (_25406_, _25395_);
  and (_25427_, _24536_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_25428_, _24557_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_25439_, _25428_, _25427_);
  not (_25450_, _24916_);
  nor (_25460_, _24415_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_25471_, _25460_, _24971_);
  and (_25482_, _25471_, _25450_);
  and (_25493_, _24601_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_25504_, _24469_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_25515_, _25504_, _25493_);
  not (_25526_, _25515_);
  nor (_25537_, _25526_, _25482_);
  and (_25548_, _25537_, _25439_);
  not (_25558_, _25548_);
  and (_25569_, _24469_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_25580_, _25569_, _25036_);
  and (_25591_, _24536_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_25602_, _25591_);
  and (_25623_, _25602_, _25580_);
  nor (_25624_, _24916_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_25635_, _25624_);
  nor (_25646_, _24927_, _24971_);
  and (_25656_, _25646_, _25635_);
  and (_25667_, _24557_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and (_25678_, _24601_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_25689_, _25678_, _25667_);
  not (_25700_, _25689_);
  nor (_25711_, _25700_, _25656_);
  and (_25722_, _25711_, _25623_);
  nor (_25733_, _25722_, _25558_);
  and (_25743_, _25733_, _25406_);
  and (_25754_, _25743_, _25254_);
  nand (_25765_, _25754_, _24906_);
  and (_25776_, _23767_, _21514_);
  not (_25787_, _25776_);
  and (_25798_, _20905_, _16162_);
  not (_25809_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_25820_, _16108_, _25809_);
  and (_25831_, _25820_, _16151_);
  not (_25841_, _25831_);
  nor (_25852_, _18216_, _18042_);
  and (_25863_, _18216_, _18042_);
  nor (_25874_, _25863_, _25852_);
  not (_25885_, _17062_);
  nor (_25896_, _17378_, _25885_);
  nor (_25907_, _17378_, _17062_);
  and (_25918_, _17378_, _17062_);
  nor (_25929_, _25918_, _25907_);
  not (_25940_, _17704_);
  nor (_25951_, _18402_, _25940_);
  nor (_25972_, _18402_, _17704_);
  and (_25973_, _18402_, _17704_);
  nor (_25984_, _25973_, _25972_);
  not (_25995_, _16722_);
  and (_26006_, _18565_, _25995_);
  nor (_26017_, _26006_, _25984_);
  nor (_26028_, _26017_, _25951_);
  nor (_26039_, _26028_, _25929_);
  nor (_26050_, _26039_, _25896_);
  and (_26061_, _26028_, _25929_);
  nor (_26082_, _26061_, _26039_);
  not (_26083_, _26082_);
  and (_26094_, _26006_, _25984_);
  nor (_26104_, _26094_, _26017_);
  not (_26115_, _26104_);
  nor (_26126_, _18565_, _16722_);
  and (_26137_, _18565_, _16722_);
  nor (_26148_, _26137_, _26126_);
  not (_26159_, _26148_);
  and (_26170_, _18935_, _17552_);
  nor (_26181_, _18935_, _17552_);
  nor (_26192_, _26181_, _26170_);
  nor (_26203_, _19436_, _16557_);
  and (_26214_, _19436_, _16557_);
  nor (_26225_, _26214_, _26203_);
  nor (_26236_, _19272_, _17868_);
  and (_26247_, _19272_, _17868_);
  nor (_26258_, _26247_, _26236_);
  not (_26269_, _16886_);
  and (_26280_, _19818_, _26269_);
  nor (_26291_, _26280_, _26258_);
  not (_26302_, _17868_);
  nor (_26313_, _19272_, _26302_);
  nor (_26324_, _26313_, _26291_);
  nor (_26335_, _26324_, _26225_);
  not (_26346_, _16557_);
  nor (_26357_, _19436_, _26346_);
  nor (_26368_, _26357_, _26335_);
  nor (_26379_, _26368_, _26192_);
  and (_26390_, _26368_, _26192_);
  nor (_26401_, _26390_, _26379_);
  not (_26412_, _26401_);
  and (_26423_, _26324_, _26225_);
  nor (_26434_, _26423_, _26335_);
  not (_26445_, _26434_);
  and (_26456_, _26280_, _26258_);
  nor (_26467_, _26456_, _26291_);
  not (_26478_, _26467_);
  nor (_26488_, _19818_, _16886_);
  and (_26499_, _19818_, _16886_);
  nor (_26510_, _26499_, _26488_);
  not (_26531_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_26532_, _16370_, _26531_);
  not (_26543_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_26554_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_26565_, _26554_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26576_, _26565_, _16952_);
  nor (_26587_, _26576_, _26543_);
  nor (_26598_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26609_, _26598_, _16612_);
  not (_26620_, _26609_);
  and (_26631_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26642_, _26631_, _17933_);
  not (_26653_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26664_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _26653_);
  and (_26675_, _26664_, _17595_);
  nor (_26686_, _26675_, _26642_);
  and (_26697_, _26686_, _26620_);
  and (_26708_, _26697_, _26587_);
  and (_26719_, _26565_, _16414_);
  nor (_26730_, _26719_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26741_, _26664_, _17759_);
  not (_26752_, _26741_);
  and (_26763_, _26631_, _17443_);
  and (_26774_, _26598_, _16777_);
  nor (_26785_, _26774_, _26763_);
  and (_26796_, _26785_, _26752_);
  and (_26807_, _26796_, _26730_);
  nor (_26828_, _26807_, _26708_);
  nor (_26829_, _26828_, _16370_);
  nor (_26840_, _26829_, _26532_);
  and (_26851_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_26861_, _26851_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_26872_, _26861_);
  and (_26883_, _26872_, _26840_);
  and (_26894_, _26872_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_26905_, _26894_, _26883_);
  nor (_26916_, _26905_, _26510_);
  and (_26937_, _26916_, _26478_);
  and (_26938_, _26937_, _26445_);
  and (_26949_, _26938_, _26412_);
  not (_26960_, _17552_);
  or (_26971_, _18935_, _26960_);
  and (_26982_, _18935_, _26960_);
  or (_26993_, _26368_, _26982_);
  and (_27004_, _26993_, _26971_);
  or (_27015_, _27004_, _26949_);
  and (_27026_, _27015_, _26159_);
  and (_27037_, _27026_, _26115_);
  and (_27048_, _27037_, _26083_);
  nor (_27059_, _27048_, _26050_);
  nor (_27070_, _27059_, _25874_);
  and (_27081_, _27059_, _25874_);
  nor (_27092_, _27081_, _27070_);
  nor (_27103_, _27092_, _25841_);
  not (_27114_, _27103_);
  not (_27125_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_27136_, _21471_, _27125_);
  and (_27157_, _27136_, _16151_);
  not (_27158_, _25874_);
  not (_27169_, _25929_);
  and (_27180_, _26126_, _25984_);
  nor (_27191_, _27180_, _25972_);
  nor (_27202_, _27191_, _27169_);
  not (_27212_, _26225_);
  and (_27223_, _26488_, _26258_);
  nor (_27234_, _27223_, _26236_);
  nor (_27245_, _27234_, _27212_);
  nor (_27256_, _27245_, _26203_);
  nor (_27267_, _27256_, _26192_);
  and (_27278_, _27256_, _26192_);
  nor (_27289_, _27278_, _27267_);
  not (_27300_, _26510_);
  nor (_27311_, _26905_, _27300_);
  and (_27322_, _27311_, _26258_);
  and (_27333_, _27234_, _27212_);
  nor (_27344_, _27333_, _27245_);
  and (_27355_, _27344_, _27322_);
  not (_27366_, _27355_);
  nor (_27377_, _27366_, _27289_);
  nor (_27388_, _27256_, _26170_);
  or (_27399_, _27388_, _26181_);
  or (_27420_, _27399_, _27377_);
  and (_27421_, _27420_, _26148_);
  nor (_27432_, _26126_, _25984_);
  nor (_27443_, _27432_, _27180_);
  and (_27454_, _27443_, _27421_);
  and (_27465_, _27191_, _27169_);
  nor (_27476_, _27465_, _27202_);
  and (_27487_, _27476_, _27454_);
  or (_27498_, _27487_, _27202_);
  nor (_27509_, _27498_, _25907_);
  nor (_27520_, _27509_, _27158_);
  and (_27531_, _27509_, _27158_);
  nor (_27542_, _27531_, _27520_);
  and (_27553_, _27542_, _27157_);
  and (_27563_, _16141_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27574_, _27563_, _25820_);
  nor (_27585_, _19818_, _19272_);
  and (_27596_, _27585_, _19447_);
  and (_27607_, _27596_, _18946_);
  and (_27618_, _27607_, _18576_);
  and (_27629_, _27618_, _18979_);
  and (_27640_, _27629_, _17389_);
  and (_27651_, _27640_, _26905_);
  not (_27662_, _26905_);
  and (_27673_, _17378_, _18402_);
  and (_27684_, _19436_, _19272_);
  and (_27705_, _27684_, _19818_);
  and (_27706_, _27705_, _18935_);
  and (_27717_, _27706_, _18565_);
  and (_27728_, _27717_, _27673_);
  and (_27739_, _27728_, _27662_);
  nor (_27750_, _27739_, _27651_);
  and (_27761_, _27750_, _18216_);
  nor (_27772_, _27750_, _18216_);
  nor (_27783_, _27772_, _27761_);
  and (_27794_, _27783_, _27574_);
  not (_27805_, _18042_);
  nor (_27816_, _26905_, _27805_);
  not (_27827_, _27816_);
  and (_27838_, _26905_, _18216_);
  and (_27849_, _27563_, _16119_);
  not (_27860_, _27849_);
  nor (_27871_, _27860_, _27838_);
  and (_27882_, _27871_, _27827_);
  nor (_27893_, _27882_, _27794_);
  and (_27904_, _27136_, _21503_);
  not (_27915_, _27673_);
  nor (_27925_, _27684_, _18935_);
  and (_27936_, _27925_, _27904_);
  and (_27947_, _27936_, _18576_);
  nor (_27958_, _27947_, _27915_);
  nor (_27969_, _27673_, _18216_);
  nor (_27980_, _27969_, _27936_);
  and (_27991_, _27980_, _26905_);
  nor (_28002_, _27991_, _27958_);
  nor (_28013_, _28002_, _18674_);
  and (_28024_, _28002_, _18674_);
  nor (_28035_, _28024_, _28013_);
  and (_28046_, _28035_, _27904_);
  and (_28057_, _27563_, _27136_);
  not (_28068_, _28057_);
  nor (_28079_, _28068_, _26905_);
  not (_28090_, _28079_);
  not (_28101_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_28112_, _16141_, _28101_);
  and (_28123_, _28112_, _27136_);
  not (_28144_, _28123_);
  nor (_28145_, _28144_, _25863_);
  and (_28156_, _28112_, _21482_);
  and (_28167_, _28156_, _25874_);
  nor (_28178_, _28167_, _28145_);
  and (_28189_, _21503_, _16119_);
  and (_28200_, _28189_, _25852_);
  and (_28211_, _25820_, _21503_);
  and (_28222_, _28211_, _18216_);
  nor (_28233_, _28222_, _28200_);
  and (_28244_, _28112_, _16108_);
  not (_28255_, _28244_);
  nor (_28266_, _28255_, _17378_);
  not (_28276_, _28266_);
  and (_28287_, _21482_, _16151_);
  not (_28298_, _28287_);
  nor (_28309_, _28298_, _18216_);
  and (_28330_, _27563_, _21482_);
  not (_28331_, _28330_);
  nor (_28342_, _28331_, _19818_);
  nor (_28353_, _28342_, _28309_);
  and (_28364_, _28353_, _28276_);
  and (_28375_, _28364_, _28233_);
  and (_28386_, _28375_, _28178_);
  and (_28397_, _28386_, _28090_);
  not (_28408_, _28397_);
  nor (_28419_, _28408_, _28046_);
  and (_28430_, _28419_, _27893_);
  not (_28441_, _28430_);
  nor (_28452_, _28441_, _27553_);
  and (_28463_, _28452_, _27114_);
  not (_28474_, _28463_);
  nor (_28485_, _28474_, _25798_);
  and (_28496_, _28485_, _25787_);
  not (_28507_, _28496_);
  or (_28518_, _28507_, _25765_);
  not (_28529_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_28540_, \oc8051_top_1.oc8051_decoder1.wr , _16097_);
  not (_28551_, _28540_);
  nor (_28562_, _28551_, _24382_);
  and (_28573_, _28562_, _28529_);
  not (_28584_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_28595_, _25765_, _28584_);
  and (_28606_, _28595_, _28573_);
  and (_28617_, _28606_, _28518_);
  nor (_28627_, _28562_, _28584_);
  not (_28638_, _27157_);
  nor (_28649_, _27520_, _25852_);
  nor (_28660_, _28649_, _28638_);
  not (_28671_, _28660_);
  and (_28682_, _18216_, _27805_);
  nor (_28693_, _28682_, _27070_);
  nor (_28704_, _28693_, _25841_);
  and (_28715_, _27958_, _26905_);
  nor (_28726_, _28715_, _27838_);
  not (_28737_, _27904_);
  nor (_28748_, _26905_, _18216_);
  not (_28759_, _28748_);
  nor (_28770_, _28759_, _27958_);
  nor (_28781_, _28770_, _28737_);
  and (_28792_, _28781_, _28726_);
  or (_28803_, _28792_, _27936_);
  nor (_28814_, _28287_, _26905_);
  nor (_28825_, _28211_, _27662_);
  nor (_28836_, _28825_, _28814_);
  not (_28847_, _28836_);
  nor (_28868_, _26894_, _26840_);
  not (_28869_, _28156_);
  nor (_28880_, _28869_, _26883_);
  not (_28891_, _28880_);
  nor (_28902_, _28331_, _26840_);
  nor (_28913_, _28902_, _28123_);
  and (_28924_, _28913_, _28891_);
  nor (_28935_, _28924_, _28868_);
  and (_28946_, _26861_, _26840_);
  and (_28956_, _28112_, _25820_);
  and (_28967_, _28189_, _26840_);
  nor (_28978_, _28967_, _28956_);
  nor (_28989_, _28978_, _28946_);
  nor (_29000_, _28068_, _19818_);
  and (_29011_, _28112_, _16119_);
  not (_29022_, _29011_);
  nor (_29033_, _29022_, _18216_);
  nor (_29044_, _29033_, _29000_);
  not (_29055_, _29044_);
  nor (_29066_, _29055_, _28989_);
  not (_29077_, _29066_);
  nor (_29088_, _29077_, _28935_);
  and (_29099_, _29088_, _28847_);
  not (_29110_, _29099_);
  nor (_29121_, _29110_, _28803_);
  not (_29132_, _29121_);
  nor (_29143_, _29132_, _28704_);
  and (_29154_, _29143_, _28671_);
  not (_29165_, _24644_);
  nor (_29176_, _24884_, _24764_);
  and (_29187_, _29176_, _29165_);
  and (_29198_, _29187_, _25754_);
  nand (_29209_, _29198_, _29154_);
  or (_29220_, _29198_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_29231_, _28562_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_29242_, _29231_, _29220_);
  and (_29253_, _29242_, _29209_);
  or (_29264_, _29253_, _28627_);
  or (_29275_, _29264_, _28617_);
  and (_06647_, _29275_, _41894_);
  and (_29295_, _23924_, _21514_);
  not (_29306_, _29295_);
  and (_29317_, _21232_, _16162_);
  nor (_29328_, _28869_, _26488_);
  nor (_29339_, _29328_, _28123_);
  or (_29350_, _29339_, _26499_);
  and (_29361_, _27563_, _27125_);
  not (_29372_, _29361_);
  nor (_29383_, _29372_, _19272_);
  and (_29394_, _28956_, _18674_);
  nor (_29415_, _29394_, _29383_);
  and (_29416_, _29415_, _29350_);
  nor (_29427_, _29022_, _26905_);
  nor (_29438_, _27860_, _16886_);
  and (_29449_, _27574_, _19818_);
  nor (_29460_, _29449_, _29438_);
  nor (_29471_, _28287_, _27904_);
  nor (_29482_, _29471_, _19818_);
  not (_29493_, _29482_);
  nand (_29504_, _29493_, _29460_);
  nor (_29515_, _29504_, _29427_);
  and (_29526_, _29515_, _29416_);
  and (_29537_, _26905_, _27300_);
  nor (_29548_, _29537_, _27311_);
  not (_29559_, _29548_);
  nor (_29570_, _27157_, _25831_);
  nor (_29581_, _29570_, _29559_);
  not (_29592_, _29581_);
  and (_29603_, _28189_, _26488_);
  and (_29613_, _28211_, _19818_);
  nor (_29624_, _29613_, _29603_);
  and (_29635_, _29624_, _29592_);
  and (_29646_, _29635_, _29526_);
  not (_29657_, _29646_);
  nor (_29678_, _29657_, _29317_);
  and (_29679_, _29678_, _29306_);
  not (_29690_, _29679_);
  or (_29701_, _29690_, _25765_);
  not (_29712_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_29723_, _25765_, _29712_);
  and (_29734_, _29723_, _28573_);
  and (_29745_, _29734_, _29701_);
  nor (_29756_, _28562_, _29712_);
  not (_29767_, _29154_);
  or (_29778_, _29767_, _25765_);
  and (_29789_, _29723_, _29231_);
  and (_29800_, _29789_, _29778_);
  or (_29811_, _29800_, _29756_);
  or (_29822_, _29811_, _29745_);
  and (_08885_, _29822_, _41894_);
  and (_29843_, _21264_, _16162_);
  not (_29854_, _29843_);
  and (_29865_, _23988_, _21514_);
  nor (_29876_, _27860_, _17868_);
  and (_29887_, _19818_, _19272_);
  nor (_29898_, _29887_, _27585_);
  not (_29909_, _29898_);
  nor (_29920_, _29909_, _26905_);
  and (_29931_, _29909_, _26905_);
  nor (_29941_, _29931_, _29920_);
  and (_29952_, _29941_, _27574_);
  nor (_29963_, _29952_, _29876_);
  nor (_29984_, _27925_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_29985_, _29984_, _19480_);
  nor (_29996_, _29984_, _19480_);
  nor (_30007_, _29996_, _29985_);
  nor (_30018_, _30007_, _28737_);
  not (_30029_, _30018_);
  and (_30040_, _28156_, _26258_);
  and (_30051_, _28189_, _26236_);
  nor (_30062_, _28144_, _26247_);
  and (_30073_, _28211_, _19272_);
  or (_30084_, _30073_, _30062_);
  or (_30095_, _30084_, _30051_);
  nor (_30106_, _30095_, _30040_);
  nor (_30117_, _28255_, _19818_);
  not (_30128_, _30117_);
  nor (_30139_, _28298_, _19272_);
  nor (_30150_, _29372_, _19436_);
  nor (_30161_, _30150_, _30139_);
  and (_30172_, _30161_, _30128_);
  and (_30183_, _30172_, _30106_);
  and (_30194_, _30183_, _30029_);
  and (_30205_, _30194_, _29963_);
  nor (_30216_, _26488_, _26258_);
  or (_30227_, _30216_, _27223_);
  and (_30238_, _30227_, _27311_);
  nor (_30248_, _30227_, _27311_);
  or (_30259_, _30248_, _30238_);
  and (_30270_, _30259_, _27157_);
  nor (_30281_, _26916_, _26478_);
  nor (_30292_, _30281_, _26937_);
  nor (_30313_, _30292_, _25841_);
  nor (_30314_, _30313_, _30270_);
  and (_30325_, _30314_, _30205_);
  not (_30336_, _30325_);
  nor (_30347_, _30336_, _29865_);
  and (_30358_, _30347_, _29854_);
  not (_30369_, _30358_);
  or (_30381_, _30369_, _25765_);
  not (_30402_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_30413_, _25765_, _30402_);
  and (_30424_, _30413_, _28573_);
  and (_30435_, _30424_, _30381_);
  nor (_30446_, _28562_, _30402_);
  nand (_30457_, _25754_, _24644_);
  not (_30468_, _24884_);
  and (_30479_, _30468_, _24764_);
  not (_30490_, _30479_);
  nor (_30501_, _30490_, _30457_);
  nand (_30512_, _30501_, _29154_);
  or (_30523_, _30501_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_30534_, _30523_, _29231_);
  and (_30545_, _30534_, _30512_);
  or (_30556_, _30545_, _30446_);
  or (_30567_, _30556_, _30435_);
  and (_08896_, _30567_, _41894_);
  and (_30587_, _21296_, _16162_);
  not (_30598_, _30587_);
  and (_30609_, _24053_, _21514_);
  nor (_30620_, _27860_, _16557_);
  nor (_30631_, _29887_, _26905_);
  nor (_30642_, _27585_, _27662_);
  nor (_30653_, _30642_, _30631_);
  and (_30664_, _30653_, _19447_);
  not (_30675_, _30664_);
  not (_30686_, _27574_);
  nor (_30697_, _30653_, _19447_);
  nor (_30708_, _30697_, _30686_);
  and (_30719_, _30708_, _30675_);
  nor (_30730_, _30719_, _30620_);
  nor (_30741_, _26937_, _26445_);
  nor (_30752_, _30741_, _26938_);
  nor (_30763_, _30752_, _25841_);
  not (_30774_, _30763_);
  nor (_30785_, _29372_, _18935_);
  and (_30806_, _28189_, _26203_);
  and (_30807_, _28211_, _19436_);
  nor (_30818_, _30807_, _30806_);
  nor (_30829_, _28144_, _26214_);
  and (_30840_, _28156_, _26225_);
  nor (_30851_, _30840_, _30829_);
  nor (_30862_, _28298_, _19436_);
  nor (_30873_, _28255_, _19272_);
  nor (_30884_, _30873_, _30862_);
  and (_30894_, _30884_, _30851_);
  nand (_30905_, _30894_, _30818_);
  nor (_30916_, _30905_, _30785_);
  and (_30927_, _30916_, _30774_);
  nor (_30938_, _27344_, _27322_);
  nor (_30949_, _30938_, _28638_);
  and (_30960_, _30949_, _27366_);
  nor (_30971_, _29996_, _19436_);
  and (_30982_, _27684_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_30993_, _30982_, _30971_);
  nor (_31004_, _30993_, _28737_);
  nor (_31015_, _31004_, _30960_);
  and (_31035_, _31015_, _30927_);
  and (_31036_, _31035_, _30730_);
  not (_31047_, _31036_);
  nor (_31058_, _31047_, _30609_);
  and (_31069_, _31058_, _30598_);
  not (_31080_, _31069_);
  or (_31091_, _31080_, _25765_);
  not (_31102_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_31113_, _25765_, _31102_);
  and (_31124_, _31113_, _28573_);
  and (_31135_, _31124_, _31091_);
  nor (_31146_, _28562_, _31102_);
  or (_31157_, _29176_, _30457_);
  and (_31168_, _31157_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_31178_, _24764_);
  and (_31189_, _24644_, _24884_);
  and (_31200_, _31189_, _31178_);
  not (_31211_, _31200_);
  nor (_31222_, _31211_, _29154_);
  and (_31233_, _24644_, _24764_);
  and (_31244_, _31233_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_31255_, _31244_, _31222_);
  and (_31266_, _31255_, _25754_);
  or (_31277_, _31266_, _31168_);
  and (_31288_, _31277_, _29231_);
  or (_31299_, _31288_, _31146_);
  or (_31310_, _31299_, _31135_);
  and (_08907_, _31310_, _41894_);
  and (_31330_, _21338_, _16162_);
  not (_31341_, _31330_);
  and (_31352_, _24133_, _21514_);
  nor (_31363_, _26938_, _26412_);
  nor (_31374_, _31363_, _26949_);
  nor (_31385_, _31374_, _25841_);
  not (_31396_, _31385_);
  not (_31407_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_31418_, _27684_, _31407_);
  nor (_31429_, _31418_, _18946_);
  or (_31440_, _31429_, _28737_);
  or (_31451_, _31440_, _27925_);
  and (_31462_, _27366_, _27289_);
  or (_31473_, _31462_, _28638_);
  nor (_31483_, _31473_, _27377_);
  nor (_31494_, _27860_, _17552_);
  and (_31505_, _27596_, _26905_);
  and (_31516_, _27705_, _27662_);
  nor (_31527_, _31516_, _31505_);
  nor (_31538_, _31527_, _18935_);
  not (_31549_, _31538_);
  and (_31560_, _31527_, _18935_);
  nor (_31571_, _31560_, _30686_);
  and (_31582_, _31571_, _31549_);
  nor (_31593_, _31582_, _31494_);
  and (_31614_, _28189_, _26181_);
  and (_31615_, _28211_, _18935_);
  nor (_31626_, _31615_, _31614_);
  nor (_31636_, _29372_, _18565_);
  not (_31647_, _31636_);
  and (_31658_, _31647_, _31626_);
  nor (_31669_, _28144_, _26170_);
  and (_31680_, _28156_, _26192_);
  nor (_31691_, _31680_, _31669_);
  nor (_31702_, _28298_, _18935_);
  nor (_31713_, _28255_, _19436_);
  nor (_31724_, _31713_, _31702_);
  and (_31735_, _31724_, _31691_);
  and (_31746_, _31735_, _31658_);
  nand (_31757_, _31746_, _31593_);
  nor (_31768_, _31757_, _31483_);
  and (_31779_, _31768_, _31451_);
  and (_31789_, _31779_, _31396_);
  not (_31800_, _31789_);
  nor (_31811_, _31800_, _31352_);
  and (_31822_, _31811_, _31341_);
  not (_31833_, _31822_);
  or (_31844_, _31833_, _25765_);
  not (_31855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_31866_, _25765_, _31855_);
  and (_31877_, _31866_, _28573_);
  and (_31888_, _31877_, _31844_);
  nor (_31899_, _28562_, _31855_);
  and (_31910_, _30457_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_31921_, _29176_, _24644_);
  not (_31932_, _31921_);
  nor (_31942_, _31932_, _29154_);
  nor (_31953_, _31233_, _31189_);
  nor (_31964_, _31953_, _31855_);
  or (_31975_, _31964_, _31942_);
  and (_31986_, _31975_, _25754_);
  or (_31997_, _31986_, _31910_);
  and (_32008_, _31997_, _29231_);
  or (_32019_, _32008_, _31899_);
  or (_32030_, _32019_, _31888_);
  and (_08918_, _32030_, _41894_);
  and (_32050_, _24189_, _21514_);
  not (_32061_, _32050_);
  and (_32072_, _21370_, _16162_);
  nor (_32083_, _27015_, _26148_);
  and (_32094_, _27015_, _26148_);
  nor (_32105_, _32094_, _32083_);
  and (_32116_, _32105_, _25831_);
  not (_32127_, _32116_);
  nor (_32138_, _27420_, _26148_);
  nor (_32148_, _32138_, _27421_);
  and (_32159_, _32148_, _27157_);
  nor (_32170_, _26905_, _16722_);
  and (_32181_, _26905_, _18576_);
  nor (_32192_, _32181_, _32170_);
  nor (_32203_, _32192_, _27860_);
  and (_32214_, _27607_, _26905_);
  and (_32225_, _27706_, _27662_);
  nor (_32246_, _32225_, _32214_);
  and (_32247_, _32246_, _18565_);
  nor (_32257_, _32246_, _18565_);
  nor (_32268_, _32257_, _32247_);
  and (_32279_, _32268_, _27574_);
  nor (_32290_, _32279_, _32203_);
  nor (_32301_, _27936_, _18576_);
  not (_32312_, _32301_);
  nor (_32323_, _27947_, _28737_);
  and (_32334_, _32323_, _32312_);
  not (_32345_, _32334_);
  and (_32356_, _28156_, _26148_);
  and (_32366_, _28189_, _26126_);
  nor (_32377_, _28144_, _26137_);
  and (_32388_, _28211_, _18565_);
  or (_32399_, _32388_, _32377_);
  or (_32410_, _32399_, _32366_);
  nor (_32421_, _32410_, _32356_);
  nor (_32432_, _28298_, _18565_);
  not (_32443_, _32432_);
  nor (_32454_, _29372_, _18402_);
  nor (_32465_, _28255_, _18935_);
  nor (_32476_, _32465_, _32454_);
  and (_32486_, _32476_, _32443_);
  and (_32497_, _32486_, _32421_);
  and (_32508_, _32497_, _32345_);
  and (_32519_, _32508_, _32290_);
  not (_32530_, _32519_);
  nor (_32551_, _32530_, _32159_);
  and (_32552_, _32551_, _32127_);
  not (_32563_, _32552_);
  nor (_32574_, _32563_, _32072_);
  and (_32585_, _32574_, _32061_);
  not (_32595_, _32585_);
  or (_32606_, _32595_, _25765_);
  not (_32617_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_32628_, _25765_, _32617_);
  and (_32639_, _32628_, _28573_);
  and (_32650_, _32639_, _32606_);
  nor (_32661_, _28562_, _32617_);
  not (_32672_, _25754_);
  and (_32683_, _24895_, _29165_);
  nor (_32694_, _24895_, _29165_);
  nor (_32704_, _32694_, _32683_);
  or (_32715_, _32704_, _32672_);
  and (_32726_, _32715_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_32737_, _32683_, _29767_);
  and (_32748_, _32694_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_32759_, _32748_, _32737_);
  and (_32770_, _32759_, _25754_);
  or (_32781_, _32770_, _32726_);
  and (_32792_, _32781_, _29231_);
  or (_32802_, _32792_, _32661_);
  or (_32813_, _32802_, _32650_);
  and (_08929_, _32813_, _41894_);
  and (_32834_, _24275_, _21514_);
  not (_32845_, _32834_);
  and (_32856_, _21426_, _16162_);
  nor (_32867_, _27443_, _27421_);
  nor (_32878_, _32867_, _27454_);
  and (_32899_, _32878_, _27157_);
  not (_32900_, _32899_);
  nor (_32910_, _27026_, _26115_);
  nor (_32921_, _32910_, _27037_);
  nor (_32932_, _32921_, _25841_);
  nor (_32943_, _26905_, _17704_);
  and (_32954_, _26905_, _18979_);
  nor (_32965_, _32954_, _32943_);
  nor (_32976_, _32965_, _27860_);
  and (_32987_, _27618_, _26905_);
  and (_32998_, _27717_, _27662_);
  nor (_33009_, _32998_, _32987_);
  and (_33019_, _33009_, _18402_);
  nor (_33030_, _33009_, _18402_);
  or (_33041_, _33030_, _30686_);
  nor (_33052_, _33041_, _33019_);
  nor (_33063_, _33052_, _32976_);
  nor (_33074_, _27991_, _27947_);
  nor (_33085_, _33074_, _18402_);
  and (_33096_, _33074_, _18402_);
  nor (_33107_, _33096_, _33085_);
  nor (_33118_, _33107_, _28737_);
  and (_33129_, _28156_, _25984_);
  nor (_33139_, _28144_, _25973_);
  not (_33150_, _33139_);
  and (_33161_, _28189_, _25972_);
  and (_33172_, _28211_, _18402_);
  nor (_33183_, _33172_, _33161_);
  nand (_33194_, _33183_, _33150_);
  nor (_33205_, _33194_, _33129_);
  nor (_33216_, _28255_, _18565_);
  not (_33227_, _33216_);
  nor (_33238_, _28298_, _18402_);
  nor (_33248_, _29372_, _17378_);
  nor (_33269_, _33248_, _33238_);
  and (_33270_, _33269_, _33227_);
  and (_33281_, _33270_, _33205_);
  not (_33292_, _33281_);
  nor (_33303_, _33292_, _33118_);
  and (_33314_, _33303_, _33063_);
  not (_33325_, _33314_);
  nor (_33336_, _33325_, _32932_);
  and (_33347_, _33336_, _32900_);
  not (_33357_, _33347_);
  nor (_33368_, _33357_, _32856_);
  and (_33379_, _33368_, _32845_);
  not (_33390_, _33379_);
  or (_33401_, _33390_, _25765_);
  not (_33412_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_33423_, _25765_, _33412_);
  and (_33434_, _33423_, _28573_);
  and (_33445_, _33434_, _33401_);
  nor (_33456_, _28562_, _33412_);
  and (_33466_, _30479_, _29165_);
  and (_33477_, _33466_, _25754_);
  nand (_33488_, _33477_, _29154_);
  or (_33499_, _33477_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_33510_, _33499_, _29231_);
  and (_33521_, _33510_, _33488_);
  or (_33532_, _33521_, _33456_);
  or (_33543_, _33532_, _33445_);
  and (_08940_, _33543_, _41894_);
  and (_33563_, _24339_, _21514_);
  not (_33574_, _33563_);
  and (_33585_, _21450_, _16162_);
  nor (_33596_, _27037_, _26083_);
  nor (_33607_, _33596_, _27048_);
  nor (_33618_, _33607_, _25841_);
  not (_33629_, _33618_);
  nor (_33640_, _27476_, _27454_);
  not (_33651_, _33640_);
  nor (_33662_, _28638_, _27487_);
  and (_33672_, _33662_, _33651_);
  and (_33683_, _26905_, _17389_);
  nor (_33694_, _26905_, _17062_);
  or (_33705_, _33694_, _33683_);
  and (_33716_, _33705_, _27849_);
  or (_33727_, _26905_, _18402_);
  or (_33738_, _32998_, _27629_);
  and (_33749_, _33738_, _33727_);
  nor (_33760_, _33749_, _17389_);
  and (_33771_, _33749_, _17389_);
  or (_33791_, _33771_, _30686_);
  nor (_33792_, _33791_, _33760_);
  nor (_33803_, _33792_, _33716_);
  and (_33814_, _33096_, _17378_);
  nor (_33825_, _33096_, _17378_);
  nor (_33836_, _33825_, _33814_);
  nor (_33847_, _33836_, _28737_);
  and (_33858_, _28156_, _25929_);
  and (_33869_, _28189_, _25907_);
  nor (_33880_, _28144_, _25918_);
  and (_33891_, _28211_, _17378_);
  or (_33901_, _33891_, _33880_);
  or (_33912_, _33901_, _33869_);
  nor (_33923_, _33912_, _33858_);
  nor (_33934_, _28298_, _17378_);
  not (_33945_, _33934_);
  nor (_33956_, _29372_, _18216_);
  nor (_33967_, _28255_, _18402_);
  nor (_33978_, _33967_, _33956_);
  and (_33989_, _33978_, _33945_);
  and (_34000_, _33989_, _33923_);
  not (_34010_, _34000_);
  nor (_34021_, _34010_, _33847_);
  and (_34032_, _34021_, _33803_);
  not (_34043_, _34032_);
  nor (_34064_, _34043_, _33672_);
  and (_34065_, _34064_, _33629_);
  not (_34076_, _34065_);
  nor (_34087_, _34076_, _33585_);
  and (_34098_, _34087_, _33574_);
  not (_34109_, _34098_);
  or (_34119_, _34109_, _25765_);
  not (_34130_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_34141_, _25765_, _34130_);
  and (_34152_, _34141_, _28573_);
  and (_34163_, _34152_, _34119_);
  nor (_34174_, _28562_, _34130_);
  nor (_34185_, _24644_, _24764_);
  and (_34196_, _34185_, _24884_);
  and (_34207_, _34196_, _25754_);
  nand (_34218_, _34207_, _29154_);
  or (_34228_, _34207_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_34239_, _34228_, _29231_);
  and (_34250_, _34239_, _34218_);
  or (_34261_, _34250_, _34174_);
  or (_34272_, _34261_, _34163_);
  and (_08950_, _34272_, _41894_);
  and (_34293_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_34303_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_34314_, _34303_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_34325_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_34336_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_34347_, _34336_, _34325_);
  and (_34358_, _34303_, _16097_);
  and (_34369_, _34358_, _34347_);
  not (_34380_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_34391_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_34402_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34413_, _34402_, _34391_);
  and (_34423_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_34434_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34445_, _34434_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_34456_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_34467_, _34456_, _34423_);
  and (_34478_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_34489_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34500_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _34489_);
  and (_34511_, _34500_, _34391_);
  and (_34522_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_34533_, _34522_, _34478_);
  and (_34543_, _34533_, _34467_);
  not (_34554_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_34565_, _34554_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34576_, _34565_, _34391_);
  and (_34587_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_34598_, _34587_);
  and (_34609_, _34434_, _34391_);
  and (_34620_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_34631_, _34434_, _34391_);
  and (_34642_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_34653_, _34642_, _34620_);
  and (_34663_, _34653_, _34598_);
  and (_34684_, _34663_, _34543_);
  and (_34685_, _34684_, _34380_);
  nor (_34696_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _34380_);
  or (_34707_, _34696_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34718_, _34707_, _34685_);
  and (_34729_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_34740_, _34729_, _34718_);
  and (_34751_, _34740_, _34369_);
  not (_34762_, _34369_);
  and (_34773_, _34347_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_34783_, _34773_, _34762_);
  nor (_34794_, _34783_, _34751_);
  and (_34805_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34816_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34827_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_34838_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_34849_, _34838_, _34827_);
  and (_34860_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34871_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_34882_, _34871_, _34860_);
  and (_34893_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_34904_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_34914_, _34904_, _34893_);
  and (_34925_, _34914_, _34882_);
  and (_34936_, _34925_, _34849_);
  nor (_34947_, _34936_, _34478_);
  and (_34958_, _34947_, _34380_);
  nor (_34969_, _34958_, _34816_);
  nor (_34980_, _34969_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34991_, _34980_, _34805_);
  nor (_35002_, _34991_, _34762_);
  and (_35013_, _34347_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_35024_, _35013_, _34762_);
  nor (_35034_, _35024_, _35002_);
  not (_35045_, _35034_);
  and (_35056_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_35067_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  or (_35078_, _34478_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35089_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_35100_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_35111_, _35100_, _35089_);
  and (_35122_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_35133_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_35144_, _35133_, _35122_);
  and (_35155_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_35166_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_35177_, _35166_, _35155_);
  and (_35188_, _35177_, _35144_);
  and (_35199_, _35188_, _35111_);
  nor (_35210_, _35199_, _35078_);
  nor (_35221_, _35210_, _35067_);
  nor (_35232_, _35221_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35243_, _35232_, _35056_);
  nor (_35254_, _35243_, _34762_);
  and (_35265_, _34347_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_35276_, _35265_, _34762_);
  nor (_35287_, _35276_, _35254_);
  not (_35298_, _35287_);
  and (_35309_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35320_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35331_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_35342_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_35353_, _35342_, _35331_);
  and (_35364_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_35375_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_35397_, _35375_, _35364_);
  and (_35398_, _35397_, _35353_);
  and (_35420_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_35421_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_35443_, _35421_, _35420_);
  and (_35444_, _35443_, _35398_);
  nor (_35466_, _35444_, _35078_);
  nor (_35467_, _35466_, _35320_);
  nor (_35478_, _35467_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35489_, _35478_, _35309_);
  nor (_35500_, _35489_, _34762_);
  and (_35511_, _34347_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_35522_, _35511_, _34762_);
  nor (_35533_, _35522_, _35500_);
  and (_35544_, _35533_, _35298_);
  and (_35555_, _35544_, _35045_);
  and (_35566_, _35555_, _34794_);
  and (_35577_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35588_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35599_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_35610_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_35621_, _35610_, _35599_);
  and (_35632_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_35643_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_35654_, _35643_, _35632_);
  and (_35665_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_35676_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_35687_, _35676_, _35665_);
  and (_35698_, _35687_, _35654_);
  and (_35709_, _35698_, _35621_);
  nor (_35720_, _35709_, _34478_);
  and (_35731_, _35720_, _34380_);
  nor (_35742_, _35731_, _35588_);
  nor (_35753_, _35742_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35764_, _35753_, _35577_);
  nor (_35775_, _35764_, _34762_);
  and (_35786_, _34347_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_35797_, _35786_, _34762_);
  nor (_35808_, _35797_, _35775_);
  not (_35819_, _35808_);
  not (_35830_, _34478_);
  and (_35841_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_35852_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_35863_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_35874_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_35885_, _35874_, _35863_);
  and (_35896_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_35907_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_35918_, _35907_, _35896_);
  nand (_35929_, _35918_, _35885_);
  or (_35940_, _35929_, _35852_);
  nor (_35951_, _35940_, _35841_);
  and (_35962_, _35951_, _35830_);
  and (_35973_, _35962_, _34380_);
  nor (_35984_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _34380_);
  nor (_35995_, _35984_, _35973_);
  nor (_36006_, _35995_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_36017_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_36028_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _36017_);
  nor (_36039_, _36028_, _36006_);
  and (_36050_, _36039_, _34369_);
  and (_36061_, _34347_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_36072_, _36061_, _34762_);
  nor (_36083_, _36072_, _36050_);
  and (_36094_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_36105_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_36116_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_36127_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_36138_, _36127_, _36116_);
  and (_36149_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_36160_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_36171_, _36160_, _36149_);
  and (_36182_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_36193_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_36204_, _36193_, _36182_);
  and (_36215_, _36204_, _36171_);
  and (_36226_, _36215_, _36138_);
  nor (_36237_, _36226_, _34478_);
  and (_36248_, _36237_, _34380_);
  or (_36259_, _36248_, _36105_);
  and (_36270_, _36259_, _36017_);
  nor (_36281_, _36270_, _36094_);
  nor (_36292_, _36281_, _34762_);
  and (_36303_, _34347_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_36314_, _36303_, _34762_);
  nor (_36325_, _36314_, _36292_);
  and (_36336_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_36347_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_36358_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_36369_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_36380_, _36369_, _36358_);
  and (_36391_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_36402_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_36413_, _36402_, _36391_);
  and (_36424_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_36435_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_36446_, _36435_, _36424_);
  and (_36457_, _36446_, _36413_);
  and (_36468_, _36457_, _36380_);
  nor (_36479_, _36468_, _34478_);
  and (_36490_, _36479_, _34380_);
  or (_36501_, _36490_, _36347_);
  and (_36512_, _36501_, _36017_);
  nor (_36523_, _36512_, _36336_);
  nor (_36534_, _36523_, _34762_);
  and (_36545_, _34347_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_36555_, _36545_, _34762_);
  nor (_36566_, _36555_, _36534_);
  and (_36577_, _36566_, _36325_);
  not (_36588_, _36577_);
  nor (_36599_, _36588_, _36083_);
  and (_36610_, _36599_, _35819_);
  and (_36621_, _36610_, _35566_);
  not (_36632_, _34794_);
  and (_36643_, _35544_, _35034_);
  and (_36654_, _36643_, _36632_);
  nor (_36665_, _35533_, _35034_);
  and (_36675_, _36665_, _35287_);
  and (_36686_, _36675_, _36632_);
  or (_36697_, _36686_, _36654_);
  and (_36708_, _36697_, _36610_);
  nor (_36719_, _36708_, _36621_);
  nor (_36730_, _36719_, _34314_);
  not (_36741_, _36730_);
  not (_36752_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_36763_, _16097_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_36774_, _36763_, _36752_);
  nor (_36785_, _35533_, _35298_);
  and (_36796_, _36083_, _35808_);
  and (_36807_, _36796_, _36577_);
  and (_36818_, _36807_, _36785_);
  and (_36829_, _36818_, _36774_);
  not (_36840_, _36829_);
  and (_36851_, _36643_, _34794_);
  not (_36862_, _36566_);
  and (_36873_, _36862_, _36325_);
  and (_36884_, _36796_, _36873_);
  and (_36895_, _36884_, _36851_);
  and (_36906_, _36884_, _35566_);
  nor (_36916_, _36906_, _36895_);
  and (_36927_, _36916_, _36840_);
  and (_36938_, _36927_, _36741_);
  nor (_36949_, _36938_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36960_, _36949_, _34293_);
  and (_36971_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_36982_, _36599_, _35808_);
  and (_36993_, _35533_, _35287_);
  and (_37004_, _36993_, _35045_);
  and (_37015_, _37004_, _36982_);
  not (_37026_, _37015_);
  and (_37036_, _36083_, _35819_);
  and (_37047_, _37036_, _36873_);
  and (_37058_, _35555_, _36632_);
  or (_37069_, _37058_, _36654_);
  nand (_37080_, _37069_, _37047_);
  and (_37091_, _37080_, _37026_);
  and (_37102_, _36665_, _35298_);
  and (_37113_, _37102_, _34794_);
  and (_37124_, _37113_, _37047_);
  and (_37135_, _36675_, _34794_);
  and (_37145_, _37135_, _36599_);
  nor (_37156_, _35533_, _35045_);
  and (_37167_, _37156_, _35298_);
  and (_37178_, _36807_, _37167_);
  nor (_37189_, _37178_, _37145_);
  not (_37200_, _37189_);
  nor (_37211_, _37200_, _37124_);
  and (_37222_, _37211_, _37091_);
  and (_37233_, _37135_, _37047_);
  and (_37244_, _37167_, _34794_);
  and (_37254_, _37244_, _37047_);
  nor (_37265_, _37254_, _37233_);
  nor (_37276_, _36566_, _36083_);
  and (_37287_, _37276_, _36325_);
  nand (_37298_, _37287_, _35566_);
  nor (_37309_, _36632_, _36325_);
  and (_37320_, _37309_, _35555_);
  and (_37331_, _36993_, _35034_);
  and (_37342_, _37331_, _34794_);
  and (_37353_, _37342_, _37047_);
  nor (_37364_, _37353_, _37320_);
  and (_37375_, _37364_, _37298_);
  and (_37386_, _37375_, _37265_);
  not (_37397_, _37047_);
  and (_37408_, _37156_, _35287_);
  and (_37419_, _37408_, _36632_);
  nor (_37427_, _37419_, _37004_);
  nor (_37435_, _37427_, _37397_);
  not (_37443_, _37435_);
  and (_37450_, _36654_, _36982_);
  and (_37458_, _36851_, _37047_);
  nor (_37466_, _37458_, _37450_);
  and (_37473_, _37466_, _37443_);
  and (_37481_, _37473_, _37386_);
  and (_37487_, _37481_, _37222_);
  and (_37488_, _37331_, _36632_);
  and (_37489_, _37488_, _37047_);
  and (_37494_, _37167_, _36632_);
  and (_37505_, _37494_, _37047_);
  nor (_37516_, _37505_, _37489_);
  and (_37527_, _36807_, _35555_);
  and (_37538_, _37408_, _34794_);
  and (_37549_, _37538_, _37047_);
  nor (_37560_, _37549_, _37527_);
  and (_37571_, _37560_, _37516_);
  and (_37582_, _37058_, _36982_);
  and (_37593_, _37244_, _36982_);
  nor (_37604_, _37593_, _37582_);
  and (_37615_, _36686_, _36982_);
  and (_37626_, _37538_, _36599_);
  nor (_37637_, _37626_, _37615_);
  and (_37648_, _37637_, _37604_);
  and (_37659_, _37648_, _37571_);
  and (_37670_, _34794_, _37004_);
  and (_37681_, _37670_, _36807_);
  not (_37692_, _36807_);
  and (_37698_, _36632_, _37004_);
  nor (_37709_, _37698_, _37488_);
  nor (_37720_, _37709_, _37692_);
  nor (_37731_, _37720_, _37681_);
  and (_37742_, _36851_, _36982_);
  and (_37753_, _37419_, _36599_);
  nor (_37764_, _37753_, _37742_);
  and (_37775_, _35566_, _36982_);
  and (_37786_, _37494_, _36982_);
  nor (_37797_, _37786_, _37775_);
  and (_37808_, _37797_, _37764_);
  and (_37819_, _37808_, _37731_);
  and (_37830_, _37819_, _37659_);
  and (_37841_, _37830_, _37487_);
  nor (_37852_, _37841_, _34314_);
  and (_37863_, _37488_, _36807_);
  nor (_37874_, _37863_, _37681_);
  not (_37885_, _36774_);
  nor (_37896_, _37885_, _37874_);
  nor (_37907_, _37896_, _36829_);
  and (_37918_, _37015_, _36763_);
  and (_37929_, _37918_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_37940_, _37929_);
  nand (_37951_, _37940_, _37907_);
  nor (_37962_, _37951_, _37852_);
  nor (_37973_, _37962_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37984_, _37973_, _36971_);
  and (_37995_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38006_, _34794_, _36325_);
  and (_38017_, _38006_, _37276_);
  and (_38028_, _37408_, _38017_);
  and (_38039_, _38017_, _37102_);
  nor (_38050_, _38039_, _38028_);
  and (_38061_, _36632_, _36325_);
  and (_38072_, _38061_, _37276_);
  and (_38083_, _37408_, _38072_);
  and (_38094_, _37287_, _37004_);
  or (_38105_, _38094_, _38083_);
  not (_38116_, _38105_);
  and (_38127_, _38072_, _36643_);
  and (_38138_, _37287_, _37167_);
  nor (_38149_, _38138_, _38127_);
  and (_38160_, _36851_, _37287_);
  and (_38171_, _37287_, _37135_);
  nor (_38182_, _38171_, _38160_);
  and (_38193_, _38182_, _38149_);
  and (_38204_, _38193_, _38116_);
  and (_38215_, _38204_, _38050_);
  and (_38226_, _37494_, _36807_);
  not (_38237_, _38226_);
  and (_38248_, _37331_, _37287_);
  and (_38259_, _38072_, _35555_);
  nor (_38270_, _38259_, _38248_);
  and (_38281_, _38270_, _37026_);
  and (_38292_, _38281_, _38237_);
  and (_38303_, _38292_, _36719_);
  and (_38314_, _38303_, _38215_);
  nor (_38325_, _38314_, _34314_);
  and (_38336_, _36774_, _36675_);
  and (_38346_, _38336_, _36807_);
  or (_38357_, _38346_, _37929_);
  nor (_38368_, _38357_, _38325_);
  nor (_38379_, _38368_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38389_, _38379_, _37995_);
  nor (_38400_, _38389_, _37984_);
  and (_38411_, _38400_, _36960_);
  and (_09495_, _38411_, _41894_);
  and (_38432_, _25253_, _25122_);
  not (_38443_, _25722_);
  nor (_38449_, _38443_, _25395_);
  and (_38450_, _38449_, _38432_);
  and (_38451_, _30479_, _24644_);
  and (_38452_, _38451_, _25548_);
  and (_38453_, _38452_, _38450_);
  and (_38454_, _38453_, _28562_);
  and (_38455_, _38454_, _28529_);
  not (_38456_, _38455_);
  and (_38457_, _38456_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_38458_, _38450_, _25548_);
  and (_38459_, _38458_, _24644_);
  and (_38460_, _38459_, _30479_);
  and (_38461_, _38460_, _28573_);
  not (_38462_, _38461_);
  nor (_38463_, _21514_, _16162_);
  and (_38464_, _27136_, _21493_);
  nor (_38465_, _28287_, _38464_);
  and (_38466_, _38465_, _28255_);
  and (_38467_, _38466_, _38463_);
  and (_38468_, _38467_, _29372_);
  nor (_38469_, _38468_, _17378_);
  not (_38470_, _38469_);
  and (_38471_, _38470_, _33923_);
  and (_38472_, _38471_, _33803_);
  nor (_38473_, _38472_, _38462_);
  nor (_38474_, _38473_, _38457_);
  and (_38475_, _38456_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38476_, _38468_, _18402_);
  not (_38477_, _38476_);
  and (_38478_, _38477_, _33205_);
  and (_38479_, _38478_, _33063_);
  nor (_38480_, _38479_, _38462_);
  nor (_38481_, _38480_, _38475_);
  and (_38482_, _38456_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38483_, _38468_, _18565_);
  not (_38484_, _38483_);
  and (_38485_, _38484_, _32421_);
  and (_38486_, _38485_, _32290_);
  nor (_38487_, _38486_, _38462_);
  nor (_38488_, _38487_, _38482_);
  and (_38489_, _38456_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38490_, _38468_, _18935_);
  not (_38491_, _38490_);
  and (_38492_, _38491_, _31626_);
  and (_38493_, _38492_, _31691_);
  and (_38494_, _38493_, _31593_);
  nor (_38495_, _38494_, _38462_);
  nor (_38496_, _38495_, _38489_);
  and (_38497_, _38456_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38498_, _38468_, _19436_);
  not (_38499_, _38498_);
  and (_38500_, _38499_, _30818_);
  and (_38501_, _38500_, _30851_);
  and (_38502_, _38501_, _30730_);
  nor (_38503_, _38502_, _38462_);
  nor (_38504_, _38503_, _38497_);
  and (_38505_, _38456_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38506_, _38468_, _19272_);
  not (_38507_, _38506_);
  and (_38508_, _38507_, _30106_);
  and (_38509_, _38508_, _29963_);
  not (_38510_, _38509_);
  and (_38511_, _38510_, _38461_);
  nor (_38512_, _38511_, _38505_);
  nor (_38513_, _38455_, _24808_);
  nor (_38514_, _38468_, _19818_);
  not (_38515_, _38514_);
  and (_38516_, _38515_, _29460_);
  and (_38517_, _38516_, _29624_);
  and (_38518_, _38517_, _29350_);
  not (_38519_, _38518_);
  and (_38520_, _38519_, _38461_);
  nor (_38521_, _38520_, _38513_);
  and (_38522_, _38521_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38523_, _38522_, _38512_);
  and (_38524_, _38523_, _38504_);
  and (_38525_, _38524_, _38496_);
  and (_38526_, _38525_, _38488_);
  and (_38527_, _38526_, _38481_);
  and (_38528_, _38527_, _38474_);
  nor (_38529_, _38455_, _25265_);
  nand (_38530_, _38529_, _38528_);
  or (_38531_, _38529_, _38528_);
  and (_38532_, _38531_, _24971_);
  and (_38533_, _38532_, _38530_);
  or (_38534_, _38455_, _25308_);
  or (_38535_, _38534_, _38533_);
  nor (_38536_, _38468_, _18216_);
  not (_38537_, _38536_);
  and (_38538_, _38537_, _28233_);
  and (_38539_, _38538_, _28178_);
  and (_38540_, _38539_, _27893_);
  nand (_38541_, _38540_, _38455_);
  and (_38542_, _38541_, _38535_);
  and (_09516_, _38542_, _41894_);
  not (_38543_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38544_, _38521_, _38543_);
  nor (_38545_, _38521_, _38543_);
  nor (_38546_, _38545_, _38544_);
  and (_38547_, _38546_, _24971_);
  nor (_38548_, _38547_, _24818_);
  nor (_38549_, _38548_, _38461_);
  nor (_38550_, _38549_, _38520_);
  nand (_10641_, _38550_, _41894_);
  nor (_38551_, _38522_, _38512_);
  nor (_38552_, _38551_, _38523_);
  nor (_38553_, _38552_, _24393_);
  nor (_38554_, _38553_, _24688_);
  nor (_38555_, _38554_, _38461_);
  nor (_38556_, _38555_, _38511_);
  nand (_10652_, _38556_, _41894_);
  nor (_38557_, _38523_, _38504_);
  nor (_38558_, _38557_, _38524_);
  nor (_38559_, _38558_, _24393_);
  nor (_38560_, _38559_, _24447_);
  nor (_38561_, _38560_, _38461_);
  nor (_38562_, _38561_, _38503_);
  nand (_10663_, _38562_, _41894_);
  nor (_38563_, _38524_, _38496_);
  nor (_38564_, _38563_, _38525_);
  nor (_38565_, _38564_, _24393_);
  nor (_38566_, _38565_, _25482_);
  nor (_38567_, _38566_, _38461_);
  nor (_38568_, _38567_, _38495_);
  nor (_10674_, _38568_, rst);
  nor (_38569_, _38525_, _38488_);
  nor (_38570_, _38569_, _38526_);
  nor (_38571_, _38570_, _24393_);
  nor (_38572_, _38571_, _25656_);
  nor (_38573_, _38572_, _38461_);
  nor (_38574_, _38573_, _38487_);
  nor (_10685_, _38574_, rst);
  nor (_38575_, _38526_, _38481_);
  nor (_38576_, _38575_, _38527_);
  nor (_38577_, _38576_, _24393_);
  nor (_38578_, _38577_, _25156_);
  nor (_38579_, _38578_, _38461_);
  nor (_38580_, _38579_, _38480_);
  nor (_10696_, _38580_, rst);
  nor (_38581_, _38527_, _38474_);
  nor (_38582_, _38581_, _38528_);
  nor (_38583_, _38582_, _24393_);
  nor (_38584_, _38583_, _25003_);
  nor (_38585_, _38584_, _38461_);
  nor (_38586_, _38585_, _38473_);
  nor (_10707_, _38586_, rst);
  and (_38587_, _28573_, _25548_);
  and (_38588_, _38587_, _31921_);
  nand (_38589_, _38588_, _38450_);
  nor (_38590_, _38589_, _28496_);
  and (_38591_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _16097_);
  and (_38592_, _38591_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38593_, _38589_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38594_, _38593_, _38592_);
  or (_38595_, _38594_, _38590_);
  nor (_38596_, _28298_, _18042_);
  nor (_38597_, _29022_, _18935_);
  and (_38598_, _27640_, _18674_);
  and (_38599_, _38598_, _26269_);
  and (_38600_, _38599_, _26302_);
  and (_38601_, _38600_, _26346_);
  and (_38602_, _38601_, _26960_);
  nor (_38603_, _38602_, _27662_);
  and (_38604_, _26905_, _16722_);
  nor (_38605_, _38604_, _38603_);
  and (_38606_, _27728_, _18216_);
  and (_38607_, _17552_, _16557_);
  and (_38608_, _17868_, _16886_);
  and (_38609_, _38608_, _38607_);
  and (_38610_, _38609_, _38606_);
  and (_38611_, _17704_, _16722_);
  and (_38612_, _38611_, _38610_);
  nor (_38613_, _38612_, _26905_);
  and (_38614_, _26905_, _17704_);
  nor (_38615_, _38614_, _38613_);
  and (_38616_, _38615_, _38605_);
  and (_38617_, _26905_, _17062_);
  nor (_38618_, _38617_, _33694_);
  and (_38619_, _38618_, _38616_);
  and (_38620_, _38619_, _27805_);
  nor (_38621_, _38619_, _27805_);
  nor (_38622_, _38621_, _38620_);
  and (_38623_, _38622_, _27574_);
  and (_38624_, _26905_, _27805_);
  nor (_38625_, _38624_, _28748_);
  nor (_38626_, _38625_, _27860_);
  or (_38627_, _38626_, _38623_);
  or (_38628_, _38627_, _38597_);
  and (_38629_, _21514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_38630_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38631_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38632_, _38631_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38633_, _38632_, _38630_);
  nor (_38634_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38635_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38636_, _38635_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38637_, _38636_, _38634_);
  nor (_38638_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38639_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38640_, _38639_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38641_, _38640_, _38638_);
  not (_38642_, _38641_);
  nor (_38643_, _38642_, _28649_);
  nor (_38644_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38645_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38646_, _38645_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38647_, _38646_, _38644_);
  and (_38648_, _38647_, _38643_);
  nor (_38649_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38650_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38651_, _38650_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38652_, _38651_, _38649_);
  and (_38653_, _38652_, _38648_);
  and (_38654_, _38653_, _38637_);
  nor (_38655_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38656_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38657_, _38656_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38658_, _38657_, _38655_);
  and (_38659_, _38658_, _38654_);
  and (_38660_, _38659_, _38633_);
  nor (_38661_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38662_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38663_, _38662_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38664_, _38663_, _38661_);
  and (_38665_, _38664_, _38660_);
  nor (_38666_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38667_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38668_, _38667_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38669_, _38668_, _38666_);
  nand (_38670_, _38669_, _38665_);
  or (_38671_, _38669_, _38665_);
  and (_38672_, _38671_, _27157_);
  and (_38673_, _38672_, _38670_);
  and (_38674_, _21201_, _16162_);
  or (_38675_, _38674_, _38673_);
  or (_38676_, _38675_, _38629_);
  or (_38677_, _38676_, _38628_);
  nor (_38678_, _38677_, _38596_);
  nand (_38679_, _38678_, _38592_);
  and (_38680_, _38679_, _41894_);
  and (_12654_, _38680_, _38595_);
  and (_38681_, _38587_, _31200_);
  and (_38682_, _38681_, _38450_);
  nor (_38683_, _38682_, _38592_);
  not (_38684_, _38683_);
  nand (_38685_, _38684_, _28496_);
  or (_38686_, _38684_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38687_, _38686_, _41894_);
  and (_12675_, _38687_, _38685_);
  nor (_38688_, _38589_, _29679_);
  and (_38689_, _38589_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38690_, _38689_, _38592_);
  or (_38691_, _38690_, _38688_);
  nor (_38692_, _28298_, _16886_);
  nor (_38693_, _29022_, _18565_);
  nor (_38694_, _28748_, _27838_);
  not (_38695_, _38694_);
  nor (_38696_, _38695_, _27750_);
  nor (_38697_, _38696_, _26269_);
  and (_38698_, _38696_, _26269_);
  nor (_38699_, _38698_, _38697_);
  and (_38700_, _38699_, _27574_);
  nor (_38701_, _27860_, _19818_);
  or (_38702_, _38701_, _38700_);
  or (_38703_, _38702_, _38693_);
  and (_38704_, _23799_, _21514_);
  and (_38705_, _38642_, _28649_);
  nor (_38706_, _38705_, _38643_);
  and (_38707_, _38706_, _27157_);
  and (_38708_, _20980_, _16162_);
  or (_38709_, _38708_, _38707_);
  or (_38710_, _38709_, _38704_);
  or (_38711_, _38710_, _38703_);
  nor (_38712_, _38711_, _38692_);
  nand (_38713_, _38712_, _38592_);
  and (_38714_, _38713_, _41894_);
  and (_13577_, _38714_, _38691_);
  nor (_38715_, _38589_, _30358_);
  and (_38716_, _38589_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38717_, _38716_, _38592_);
  or (_38718_, _38717_, _38715_);
  nor (_38719_, _28298_, _17868_);
  nor (_38720_, _29022_, _18402_);
  nor (_38721_, _38599_, _27662_);
  and (_38722_, _38606_, _16886_);
  nor (_38723_, _38722_, _26905_);
  or (_38724_, _38723_, _38721_);
  and (_38725_, _38724_, _17868_);
  nor (_38726_, _38724_, _17868_);
  or (_38727_, _38726_, _30686_);
  nor (_38728_, _38727_, _38725_);
  nor (_38729_, _27860_, _19272_);
  or (_38730_, _38729_, _38728_);
  or (_38731_, _38730_, _38720_);
  and (_38732_, _22798_, _21514_);
  nor (_38733_, _38647_, _38643_);
  nor (_38734_, _38733_, _38648_);
  and (_38735_, _38734_, _27157_);
  and (_38736_, _21011_, _16162_);
  or (_38737_, _38736_, _38735_);
  or (_38738_, _38737_, _38732_);
  or (_38739_, _38738_, _38731_);
  nor (_38740_, _38739_, _38719_);
  nand (_38741_, _38740_, _38592_);
  and (_38742_, _38741_, _41894_);
  and (_13587_, _38742_, _38718_);
  nor (_38743_, _38589_, _31069_);
  and (_38744_, _38589_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38745_, _38744_, _38592_);
  or (_38746_, _38745_, _38743_);
  nor (_38747_, _28298_, _16557_);
  nor (_38748_, _29022_, _17378_);
  and (_38749_, _38722_, _17868_);
  and (_38750_, _38749_, _27662_);
  and (_38751_, _38600_, _26905_);
  nor (_38752_, _38751_, _38750_);
  and (_38753_, _38752_, _16557_);
  nor (_38754_, _38752_, _16557_);
  nor (_38755_, _38754_, _38753_);
  and (_38756_, _38755_, _27574_);
  nor (_38757_, _27860_, _19436_);
  or (_38758_, _38757_, _38756_);
  or (_38759_, _38758_, _38748_);
  and (_38760_, _21514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38761_, _38652_, _38648_);
  nor (_38762_, _38761_, _38653_);
  and (_38763_, _38762_, _27157_);
  and (_38764_, _21043_, _16162_);
  or (_38765_, _38764_, _38763_);
  or (_38766_, _38765_, _38760_);
  or (_38767_, _38766_, _38759_);
  nor (_38768_, _38767_, _38747_);
  nand (_38769_, _38768_, _38592_);
  and (_38770_, _38769_, _41894_);
  and (_13597_, _38770_, _38746_);
  nor (_38771_, _38589_, _31822_);
  and (_38772_, _38589_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38773_, _38772_, _38592_);
  or (_38774_, _38773_, _38771_);
  nor (_38775_, _28298_, _17552_);
  nor (_38776_, _38601_, _26960_);
  not (_38777_, _38776_);
  and (_38778_, _38777_, _38603_);
  and (_38779_, _38749_, _16557_);
  nor (_38780_, _38779_, _17552_);
  nor (_38781_, _38780_, _38610_);
  nor (_38782_, _38781_, _26905_);
  nor (_38783_, _38782_, _38778_);
  nor (_38784_, _38783_, _30686_);
  nor (_38785_, _27860_, _18935_);
  or (_38786_, _38785_, _38784_);
  or (_38787_, _38786_, _29033_);
  and (_38788_, _21514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_38789_, _38653_, _38637_);
  nor (_38790_, _38789_, _38654_);
  and (_38791_, _38790_, _27157_);
  and (_38792_, _21074_, _16162_);
  or (_38793_, _38792_, _38791_);
  or (_38794_, _38793_, _38788_);
  or (_38795_, _38794_, _38787_);
  nor (_38796_, _38795_, _38775_);
  nand (_38797_, _38796_, _38592_);
  and (_38798_, _38797_, _41894_);
  and (_13607_, _38798_, _38774_);
  nor (_38799_, _38589_, _32585_);
  and (_38800_, _38589_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38801_, _38800_, _38592_);
  or (_38802_, _38801_, _38799_);
  nor (_38803_, _28298_, _16722_);
  nor (_38804_, _29022_, _19818_);
  nor (_38805_, _38610_, _26905_);
  nor (_38806_, _38805_, _38603_);
  nor (_38807_, _38806_, _25995_);
  and (_38808_, _38806_, _25995_);
  nor (_38809_, _38808_, _38807_);
  and (_38810_, _38809_, _27574_);
  nor (_38811_, _26905_, _18576_);
  or (_38812_, _38811_, _27860_);
  nor (_38813_, _38812_, _38604_);
  or (_38814_, _38813_, _38810_);
  or (_38815_, _38814_, _38804_);
  and (_38816_, _21514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38817_, _38658_, _38654_);
  nor (_38818_, _38817_, _38659_);
  and (_38819_, _38818_, _27157_);
  and (_38820_, _21106_, _16162_);
  or (_38821_, _38820_, _38819_);
  or (_38822_, _38821_, _38816_);
  or (_38823_, _38822_, _38815_);
  nor (_38824_, _38823_, _38803_);
  nand (_38825_, _38824_, _38592_);
  and (_38826_, _38825_, _41894_);
  and (_13616_, _38826_, _38802_);
  nor (_38827_, _38589_, _33379_);
  and (_38828_, _38589_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38829_, _38828_, _38592_);
  or (_38830_, _38829_, _38827_);
  nor (_38831_, _28298_, _17704_);
  nor (_38832_, _29022_, _19272_);
  and (_38833_, _38610_, _16722_);
  nor (_38834_, _38833_, _26905_);
  not (_38835_, _38834_);
  and (_38836_, _38835_, _38605_);
  and (_38837_, _38836_, _17704_);
  nor (_38838_, _38836_, _17704_);
  nor (_38839_, _38838_, _38837_);
  nor (_38840_, _38839_, _30686_);
  nor (_38841_, _26905_, _18979_);
  or (_38842_, _38841_, _27860_);
  nor (_38843_, _38842_, _38614_);
  or (_38844_, _38843_, _38840_);
  or (_38845_, _38844_, _38832_);
  and (_38846_, _21514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_38847_, _38659_, _38633_);
  nor (_38848_, _38847_, _38660_);
  and (_38849_, _38848_, _27157_);
  and (_38850_, _21138_, _16162_);
  or (_38851_, _38850_, _38849_);
  or (_38852_, _38851_, _38846_);
  or (_38853_, _38852_, _38845_);
  nor (_38854_, _38853_, _38831_);
  nand (_38855_, _38854_, _38592_);
  and (_38856_, _38855_, _41894_);
  and (_13625_, _38856_, _38830_);
  nor (_38857_, _38589_, _34098_);
  and (_38858_, _38589_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38859_, _38858_, _38592_);
  or (_38860_, _38859_, _38857_);
  nor (_38861_, _28298_, _17062_);
  nor (_38862_, _29022_, _19436_);
  nor (_38863_, _38616_, _17062_);
  and (_38865_, _38616_, _17062_);
  nor (_38868_, _38865_, _38863_);
  nor (_38869_, _38868_, _30686_);
  nor (_38870_, _26905_, _17389_);
  or (_38871_, _38870_, _27860_);
  nor (_38872_, _38871_, _38617_);
  or (_38873_, _38872_, _38869_);
  or (_38874_, _38873_, _38862_);
  and (_38875_, _21514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_38876_, _38664_, _38660_);
  not (_38877_, _38876_);
  nor (_38878_, _38665_, _28638_);
  and (_38887_, _38878_, _38877_);
  and (_38893_, _21169_, _16162_);
  or (_38899_, _38893_, _38887_);
  or (_38903_, _38899_, _38875_);
  or (_38904_, _38903_, _38874_);
  nor (_38905_, _38904_, _38861_);
  nand (_38906_, _38905_, _38592_);
  and (_38907_, _38906_, _41894_);
  and (_13635_, _38907_, _38860_);
  nand (_38908_, _38684_, _29679_);
  or (_38909_, _38684_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_38910_, _38909_, _41894_);
  and (_13644_, _38910_, _38908_);
  nand (_38911_, _38684_, _30358_);
  or (_38912_, _38684_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38913_, _38912_, _41894_);
  and (_13654_, _38913_, _38911_);
  nand (_38914_, _38684_, _31069_);
  or (_38915_, _38684_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38916_, _38915_, _41894_);
  and (_13664_, _38916_, _38914_);
  nand (_38917_, _38684_, _31822_);
  or (_38918_, _38684_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38919_, _38918_, _41894_);
  and (_13674_, _38919_, _38917_);
  nand (_38920_, _38684_, _32585_);
  or (_38921_, _38684_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38922_, _38921_, _41894_);
  and (_13683_, _38922_, _38920_);
  nand (_38925_, _38684_, _33379_);
  or (_38926_, _38684_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38927_, _38926_, _41894_);
  and (_13692_, _38927_, _38925_);
  nand (_38928_, _38684_, _34098_);
  or (_38929_, _38684_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38930_, _38929_, _41894_);
  and (_13702_, _38930_, _38928_);
  and (_38931_, _28573_, _24906_);
  nor (_38932_, _25122_, _25395_);
  and (_38933_, _25733_, _25253_);
  and (_38934_, _38933_, _38932_);
  and (_38935_, _38934_, _38931_);
  nand (_38936_, _38935_, _38540_);
  and (_38937_, _38934_, _29231_);
  not (_38938_, _29187_);
  nor (_38939_, _38938_, _29154_);
  not (_38940_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38941_, _29187_, _38940_);
  or (_38942_, _38941_, _38939_);
  and (_38943_, _38942_, _38937_);
  nor (_38944_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_38945_, _38944_);
  nand (_38946_, _38945_, _29154_);
  and (_38947_, _38944_, _38940_);
  nor (_38948_, _38947_, _38937_);
  and (_38949_, _38948_, _38946_);
  or (_38950_, _38949_, _38935_);
  or (_38951_, _38950_, _38943_);
  and (_38952_, _38951_, _38936_);
  and (_16447_, _38952_, _41894_);
  not (_38953_, _38935_);
  nor (_38954_, _38953_, _38509_);
  not (_38955_, _25122_);
  and (_38956_, _38933_, _38955_);
  and (_38957_, _29231_, _25406_);
  and (_38958_, _38957_, _38956_);
  and (_38960_, _38958_, _38451_);
  or (_38963_, _38960_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_38969_, _38963_, _38953_);
  nand (_38974_, _38960_, _29154_);
  and (_38981_, _38974_, _38969_);
  or (_38988_, _38981_, _38954_);
  and (_21381_, _38988_, _41894_);
  nor (_38998_, _38953_, _38502_);
  or (_38999_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_39000_, _21264_, _21232_);
  or (_39001_, _39000_, _21296_);
  or (_39002_, _39001_, _21338_);
  or (_39003_, _39002_, _21370_);
  or (_39004_, _39003_, _21426_);
  or (_39005_, _39004_, _20905_);
  and (_39006_, _39005_, _16162_);
  not (_39007_, _25852_);
  nand (_39008_, _27509_, _39007_);
  or (_39009_, _27509_, _25863_);
  and (_39010_, _27157_, _39009_);
  and (_39011_, _39010_, _39008_);
  and (_39012_, _38611_, _22700_);
  and (_39013_, _38609_, _21514_);
  nand (_39014_, _39013_, _39012_);
  nand (_39015_, _39014_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_39016_, _39015_, _39011_);
  or (_39017_, _28693_, _27059_);
  not (_39018_, _28682_);
  nand (_39019_, _39018_, _27059_);
  and (_39020_, _39019_, _25831_);
  and (_39021_, _39020_, _39017_);
  or (_39022_, _39021_, _39016_);
  or (_39023_, _39022_, _33585_);
  or (_39024_, _39023_, _39006_);
  and (_39025_, _39024_, _38999_);
  or (_39026_, _39025_, _38937_);
  nand (_39027_, _31211_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand (_39028_, _39027_, _38937_);
  or (_39029_, _39028_, _31222_);
  and (_39030_, _39029_, _38953_);
  and (_39031_, _39030_, _39026_);
  or (_39032_, _39031_, _38998_);
  and (_21392_, _39032_, _41894_);
  not (_39033_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_39037_, _38937_, _31921_);
  nand (_39048_, _39037_, _39033_);
  and (_39051_, _39048_, _38953_);
  or (_39052_, _39037_, _29767_);
  and (_39053_, _39052_, _39051_);
  nor (_39062_, _38953_, _38494_);
  or (_39070_, _39062_, _39053_);
  and (_21404_, _39070_, _41894_);
  not (_39071_, _38958_);
  or (_39072_, _39071_, _32704_);
  and (_39073_, _39072_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_39074_, _32694_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_39075_, _39074_, _32737_);
  and (_39076_, _39075_, _38937_);
  or (_39077_, _39076_, _39073_);
  and (_39078_, _39077_, _38953_);
  nor (_39079_, _38953_, _38486_);
  or (_39080_, _39079_, _39078_);
  and (_21415_, _39080_, _41894_);
  nor (_39081_, _38953_, _38479_);
  and (_39082_, _38958_, _33466_);
  or (_39083_, _39082_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_39084_, _39083_, _38953_);
  nand (_39085_, _39082_, _29154_);
  and (_39086_, _39085_, _39084_);
  or (_39087_, _39086_, _39081_);
  and (_21427_, _39087_, _41894_);
  nor (_39088_, _38953_, _38472_);
  and (_39089_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_39090_, _27157_, _27420_);
  and (_39091_, _27015_, _25831_);
  or (_39092_, _39091_, _39090_);
  and (_39093_, _39092_, _39089_);
  nand (_39094_, _39089_, _28298_);
  and (_39095_, _39094_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_39096_, _39095_, _38937_);
  or (_39097_, _39096_, _39093_);
  not (_39098_, _34196_);
  nor (_39099_, _39098_, _29154_);
  nor (_39100_, _34196_, _31407_);
  or (_39101_, _39100_, _39099_);
  or (_39102_, _39101_, _39071_);
  and (_39103_, _39102_, _39097_);
  and (_39104_, _39103_, _38953_);
  or (_39105_, _39104_, _39088_);
  and (_21438_, _39105_, _41894_);
  not (_39106_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39107_, _38591_, _39106_);
  and (_39108_, _39107_, _38678_);
  nor (_39109_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_39110_, _39109_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39111_, _24906_, _25548_);
  not (_39112_, _25253_);
  and (_39113_, _25722_, _39112_);
  and (_39114_, _39113_, _28573_);
  and (_39115_, _39114_, _39111_);
  and (_39116_, _39115_, _38932_);
  nor (_39117_, _39116_, _39110_);
  nor (_39118_, _39117_, _28496_);
  and (_39119_, _25722_, _25548_);
  and (_39120_, _39119_, _25254_);
  and (_39121_, _39120_, _38957_);
  and (_39122_, _39121_, _29187_);
  and (_39123_, _39122_, _29154_);
  nor (_39124_, _39122_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_39125_, _39124_);
  not (_39126_, _39107_);
  and (_39127_, _39117_, _39126_);
  and (_39128_, _39127_, _39125_);
  not (_39129_, _39128_);
  nor (_39130_, _39129_, _39123_);
  nor (_39131_, _39130_, _39107_);
  not (_39132_, _39131_);
  nor (_39133_, _39132_, _39118_);
  nor (_39134_, _39133_, _39108_);
  and (_22208_, _39134_, _41894_);
  nor (_39135_, _39117_, _29679_);
  and (_39136_, _39121_, _24906_);
  and (_39137_, _39136_, _29154_);
  nor (_39138_, _39136_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not (_39139_, _39138_);
  and (_39140_, _39139_, _39127_);
  not (_39141_, _39140_);
  nor (_39142_, _39141_, _39137_);
  or (_39143_, _39142_, _39135_);
  and (_39144_, _39143_, _39126_);
  nor (_39145_, _39126_, _38712_);
  or (_39146_, _39145_, _39144_);
  and (_24064_, _39146_, _41894_);
  and (_39147_, _39107_, _38740_);
  nor (_39148_, _39117_, _30358_);
  and (_39149_, _39121_, _38451_);
  and (_39150_, _39149_, _29154_);
  nor (_39151_, _39149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not (_39152_, _39151_);
  and (_39153_, _39152_, _39127_);
  not (_39154_, _39153_);
  nor (_39155_, _39154_, _39150_);
  nor (_39156_, _39155_, _39107_);
  not (_39157_, _39156_);
  nor (_39158_, _39157_, _39148_);
  nor (_39159_, _39158_, _39147_);
  and (_24075_, _39159_, _41894_);
  nor (_39160_, _39117_, _31069_);
  and (_39161_, _39121_, _31200_);
  and (_39162_, _39161_, _29154_);
  nor (_39163_, _39161_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_39164_, _39163_);
  and (_39165_, _39164_, _39127_);
  not (_39166_, _39165_);
  nor (_39167_, _39166_, _39162_);
  or (_39168_, _39167_, _39160_);
  and (_39169_, _39168_, _39126_);
  nor (_39170_, _39126_, _38768_);
  or (_39171_, _39170_, _39169_);
  and (_24087_, _39171_, _41894_);
  nor (_39172_, _39117_, _31822_);
  not (_39173_, _39121_);
  and (_39174_, _39127_, _39173_);
  and (_39175_, _39174_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_39176_, _31932_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39177_, _39176_, _31942_);
  and (_39178_, _39121_, _39126_);
  not (_39179_, _39178_);
  nor (_39180_, _39179_, _39177_);
  and (_39181_, _39180_, _39127_);
  nor (_39182_, _39181_, _39175_);
  and (_39183_, _39182_, _39126_);
  not (_39184_, _39183_);
  nor (_39185_, _39184_, _39172_);
  and (_39186_, _39107_, _38796_);
  or (_39187_, _39186_, _39185_);
  nor (_24098_, _39187_, rst);
  nor (_39188_, _39117_, _32585_);
  and (_39189_, _39121_, _32683_);
  and (_39190_, _39189_, _29154_);
  nor (_39191_, _39189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_39192_, _39191_);
  and (_39193_, _39192_, _39127_);
  not (_39194_, _39193_);
  nor (_39195_, _39194_, _39190_);
  or (_39196_, _39195_, _39188_);
  and (_39197_, _39196_, _39126_);
  nor (_39198_, _39126_, _38824_);
  or (_39199_, _39198_, _39197_);
  and (_24110_, _39199_, _41894_);
  nor (_39200_, _39117_, _33379_);
  and (_39201_, _39121_, _33466_);
  and (_39202_, _39201_, _29154_);
  nor (_39203_, _39201_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_39204_, _39203_);
  and (_39205_, _39204_, _39127_);
  not (_39206_, _39205_);
  nor (_39207_, _39206_, _39202_);
  or (_39208_, _39207_, _39200_);
  and (_39209_, _39208_, _39126_);
  nor (_39210_, _39126_, _38854_);
  or (_39211_, _39210_, _39209_);
  and (_24122_, _39211_, _41894_);
  nor (_39212_, _39117_, _34098_);
  and (_39213_, _39121_, _34196_);
  and (_39214_, _39213_, _29154_);
  nor (_39215_, _39213_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not (_39216_, _39215_);
  and (_39217_, _39216_, _39127_);
  not (_39218_, _39217_);
  nor (_39219_, _39218_, _39214_);
  or (_39220_, _39219_, _39212_);
  and (_39221_, _39220_, _39126_);
  nor (_39222_, _39126_, _38905_);
  or (_39223_, _39222_, _39221_);
  and (_24134_, _39223_, _41894_);
  and (_39224_, _38458_, _29187_);
  nand (_39225_, _39224_, _29154_);
  or (_39226_, _39224_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39227_, _39226_, _29231_);
  and (_39228_, _39227_, _39225_);
  and (_39229_, _38450_, _39111_);
  nand (_39230_, _39229_, _38540_);
  or (_39231_, _39229_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39232_, _39231_, _28573_);
  and (_39233_, _39232_, _39230_);
  not (_39234_, _28562_);
  and (_39235_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_39236_, _39235_, rst);
  or (_39237_, _39236_, _39233_);
  or (_35386_, _39237_, _39228_);
  nor (_39238_, _38955_, _25395_);
  and (_39239_, _38933_, _39238_);
  and (_39240_, _39239_, _29187_);
  nand (_39241_, _39240_, _29154_);
  or (_39242_, _39240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39243_, _39242_, _29231_);
  and (_39244_, _39243_, _39241_);
  and (_39251_, _39239_, _24906_);
  not (_39262_, _39251_);
  nor (_39273_, _39262_, _38540_);
  and (_39283_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_39289_, _39283_, _39273_);
  and (_39299_, _39289_, _28573_);
  and (_39310_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_39321_, _39310_, rst);
  or (_39332_, _39321_, _39299_);
  or (_35409_, _39332_, _39244_);
  and (_39353_, _39112_, _25122_);
  and (_39364_, _39353_, _39119_);
  and (_39375_, _39364_, _25406_);
  and (_39386_, _39375_, _29187_);
  nand (_39397_, _39386_, _29154_);
  or (_39408_, _39386_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39419_, _39408_, _29231_);
  and (_39430_, _39419_, _39397_);
  and (_39441_, _39113_, _39238_);
  and (_39452_, _39441_, _39111_);
  not (_39458_, _39452_);
  nor (_39459_, _39458_, _38540_);
  and (_39460_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_39461_, _39460_, _39459_);
  and (_39462_, _39461_, _28573_);
  and (_39463_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_39464_, _39463_, rst);
  or (_39465_, _39464_, _39462_);
  or (_35432_, _39465_, _39430_);
  and (_39466_, _39353_, _25743_);
  and (_39467_, _39466_, _29187_);
  nand (_39468_, _39467_, _29154_);
  or (_39469_, _39467_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_39470_, _39469_, _29231_);
  and (_39471_, _39470_, _39468_);
  nor (_39472_, _25722_, _25253_);
  and (_39473_, _39238_, _39472_);
  and (_39474_, _39473_, _39111_);
  not (_39475_, _39474_);
  nor (_39476_, _39475_, _38540_);
  and (_39477_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_39478_, _39477_, _39476_);
  and (_39479_, _39478_, _28573_);
  and (_39480_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_39481_, _39480_, rst);
  or (_39482_, _39481_, _39479_);
  or (_35455_, _39482_, _39471_);
  not (_39483_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39484_, _39229_, _39483_);
  nand (_39485_, _38458_, _24906_);
  nor (_39486_, _39485_, _29154_);
  or (_39487_, _39486_, _39484_);
  and (_39488_, _39487_, _29231_);
  and (_39489_, _39229_, _38519_);
  or (_39490_, _39489_, _39484_);
  and (_39491_, _39490_, _28573_);
  nor (_39492_, _28562_, _39483_);
  or (_39493_, _39492_, rst);
  or (_39494_, _39493_, _39491_);
  or (_41298_, _39494_, _39488_);
  or (_39495_, _38453_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39496_, _39495_, _29231_);
  nand (_39497_, _38460_, _29154_);
  and (_39498_, _39497_, _39496_);
  nand (_39499_, _39229_, _38509_);
  or (_39500_, _39229_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39501_, _39500_, _28573_);
  and (_39502_, _39501_, _39499_);
  and (_39503_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_39504_, _39503_, rst);
  or (_39505_, _39504_, _39502_);
  or (_41300_, _39505_, _39498_);
  not (_39506_, _31953_);
  nand (_39507_, _38458_, _39506_);
  and (_39508_, _39507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39509_, _31233_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39510_, _39509_, _31222_);
  and (_39511_, _39510_, _38458_);
  or (_39512_, _39511_, _39508_);
  and (_39513_, _39512_, _29231_);
  nand (_39514_, _39229_, _38502_);
  or (_39515_, _39229_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39516_, _39515_, _28573_);
  and (_39517_, _39516_, _39514_);
  and (_39518_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39519_, _39518_, rst);
  or (_39520_, _39519_, _39517_);
  or (_41302_, _39520_, _39513_);
  not (_39521_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_39522_, _38459_, _39521_);
  nor (_39523_, _31953_, _39521_);
  or (_39524_, _39523_, _31942_);
  and (_39525_, _39524_, _38458_);
  or (_39526_, _39525_, _39522_);
  and (_39527_, _39526_, _29231_);
  nand (_39528_, _39229_, _38494_);
  or (_39529_, _39229_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39530_, _39529_, _28573_);
  and (_39531_, _39530_, _39528_);
  nor (_39532_, _28562_, _39521_);
  or (_39533_, _39532_, rst);
  or (_39534_, _39533_, _39531_);
  or (_41303_, _39534_, _39527_);
  not (_39535_, _38458_);
  or (_39536_, _39535_, _32704_);
  and (_39537_, _39536_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39538_, _32694_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39539_, _39538_, _32737_);
  and (_39540_, _39539_, _38458_);
  or (_39541_, _39540_, _39537_);
  and (_39542_, _39541_, _29231_);
  nand (_39543_, _39229_, _38486_);
  or (_39544_, _39229_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39545_, _39544_, _28573_);
  and (_39546_, _39545_, _39543_);
  and (_39547_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39548_, _39547_, rst);
  or (_39549_, _39548_, _39546_);
  or (_41305_, _39549_, _39542_);
  and (_39550_, _38458_, _33466_);
  nand (_39551_, _39550_, _29154_);
  or (_39552_, _39550_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39553_, _39552_, _29231_);
  and (_39554_, _39553_, _39551_);
  nand (_39555_, _39229_, _38479_);
  or (_39556_, _39229_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39557_, _39556_, _28573_);
  and (_39558_, _39557_, _39555_);
  and (_39559_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39560_, _39559_, rst);
  or (_39561_, _39560_, _39558_);
  or (_41307_, _39561_, _39554_);
  and (_39562_, _38458_, _34196_);
  nand (_39563_, _39562_, _29154_);
  or (_39564_, _39562_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39565_, _39564_, _29231_);
  and (_39566_, _39565_, _39563_);
  nand (_39567_, _39229_, _38472_);
  or (_39568_, _39229_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39569_, _39568_, _28573_);
  and (_39570_, _39569_, _39567_);
  and (_39571_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39572_, _39571_, rst);
  or (_39573_, _39572_, _39570_);
  or (_41309_, _39573_, _39566_);
  nand (_39574_, _39251_, _29154_);
  or (_39575_, _39251_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39576_, _39575_, _29231_);
  and (_39577_, _39576_, _39574_);
  and (_39578_, _39251_, _38519_);
  and (_39579_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_39580_, _39579_, _39578_);
  and (_39581_, _39580_, _28573_);
  and (_39582_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_39583_, _39582_, rst);
  or (_39584_, _39583_, _39581_);
  or (_41310_, _39584_, _39577_);
  and (_39585_, _39239_, _38451_);
  nand (_39586_, _39585_, _29154_);
  or (_39587_, _39585_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39588_, _39587_, _29231_);
  and (_39589_, _39588_, _39586_);
  nor (_39590_, _39262_, _38509_);
  and (_39591_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39592_, _39591_, _39590_);
  and (_39593_, _39592_, _28573_);
  and (_39594_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39595_, _39594_, rst);
  or (_39596_, _39595_, _39593_);
  or (_41312_, _39596_, _39589_);
  and (_39597_, _39239_, _31200_);
  nand (_39598_, _39597_, _29154_);
  or (_39599_, _39597_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39600_, _39599_, _29231_);
  and (_39601_, _39600_, _39598_);
  nor (_39602_, _39262_, _38502_);
  and (_39603_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39604_, _39603_, _39602_);
  and (_39605_, _39604_, _28573_);
  and (_39606_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39607_, _39606_, rst);
  or (_39608_, _39607_, _39605_);
  or (_41314_, _39608_, _39601_);
  and (_39609_, _39239_, _31921_);
  nand (_39610_, _39609_, _29154_);
  or (_39611_, _39609_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39612_, _39611_, _29231_);
  and (_39613_, _39612_, _39610_);
  nor (_39614_, _39262_, _38494_);
  and (_39615_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39616_, _39615_, _39614_);
  and (_39617_, _39616_, _28573_);
  and (_39618_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39619_, _39618_, rst);
  or (_39620_, _39619_, _39617_);
  or (_41316_, _39620_, _39613_);
  and (_39621_, _39239_, _32683_);
  nand (_39622_, _39621_, _29154_);
  or (_39623_, _39621_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39624_, _39623_, _29231_);
  and (_39625_, _39624_, _39622_);
  nor (_39626_, _39262_, _38486_);
  and (_39627_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39628_, _39627_, _39626_);
  and (_39629_, _39628_, _28573_);
  and (_39630_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39631_, _39630_, rst);
  or (_39632_, _39631_, _39629_);
  or (_41317_, _39632_, _39625_);
  and (_39633_, _39239_, _33466_);
  nand (_39634_, _39633_, _29154_);
  or (_39635_, _39633_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39636_, _39635_, _29231_);
  and (_39637_, _39636_, _39634_);
  nor (_39638_, _39262_, _38479_);
  and (_39639_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39640_, _39639_, _39638_);
  and (_39641_, _39640_, _28573_);
  and (_39642_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39643_, _39642_, rst);
  or (_39644_, _39643_, _39641_);
  or (_41319_, _39644_, _39637_);
  and (_39645_, _39239_, _34196_);
  nand (_39646_, _39645_, _29154_);
  or (_39647_, _39645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39648_, _39647_, _29231_);
  and (_39649_, _39648_, _39646_);
  nor (_39650_, _39262_, _38472_);
  and (_39651_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39652_, _39651_, _39650_);
  and (_39653_, _39652_, _28573_);
  and (_39654_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39655_, _39654_, rst);
  or (_39656_, _39655_, _39653_);
  or (_41321_, _39656_, _39649_);
  nand (_39657_, _39452_, _29154_);
  or (_39658_, _39452_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39659_, _39658_, _29231_);
  and (_39660_, _39659_, _39657_);
  and (_39661_, _39452_, _38519_);
  and (_39662_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_39663_, _39662_, _39661_);
  and (_39664_, _39663_, _28573_);
  and (_39665_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_39666_, _39665_, rst);
  or (_39667_, _39666_, _39664_);
  or (_41323_, _39667_, _39660_);
  and (_39671_, _39375_, _38451_);
  nand (_39674_, _39671_, _29154_);
  or (_39675_, _39671_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39676_, _39675_, _29231_);
  and (_39677_, _39676_, _39674_);
  nor (_39678_, _39458_, _38509_);
  and (_39679_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39680_, _39679_, _39678_);
  and (_39681_, _39680_, _28573_);
  and (_39682_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39683_, _39682_, rst);
  or (_39684_, _39683_, _39681_);
  or (_41324_, _39684_, _39677_);
  and (_39685_, _39375_, _31200_);
  nand (_39686_, _39685_, _29154_);
  or (_39687_, _39685_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39688_, _39687_, _29231_);
  and (_39689_, _39688_, _39686_);
  nor (_39690_, _39458_, _38502_);
  and (_39691_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39692_, _39691_, _39690_);
  and (_39693_, _39692_, _28573_);
  and (_39694_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39695_, _39694_, rst);
  or (_39696_, _39695_, _39693_);
  or (_41326_, _39696_, _39689_);
  and (_39697_, _39375_, _31921_);
  nand (_39698_, _39697_, _29154_);
  or (_39699_, _39697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39700_, _39699_, _29231_);
  and (_39706_, _39700_, _39698_);
  nor (_39717_, _39458_, _38494_);
  and (_39728_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39732_, _39728_, _39717_);
  and (_39733_, _39732_, _28573_);
  and (_39734_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39735_, _39734_, rst);
  or (_39736_, _39735_, _39733_);
  or (_41328_, _39736_, _39706_);
  and (_39737_, _39375_, _32683_);
  nand (_39738_, _39737_, _29154_);
  or (_39739_, _39737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39740_, _39739_, _29231_);
  and (_39741_, _39740_, _39738_);
  nor (_39742_, _39458_, _38486_);
  and (_39743_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39744_, _39743_, _39742_);
  and (_39745_, _39744_, _28573_);
  and (_39746_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39747_, _39746_, rst);
  or (_39748_, _39747_, _39745_);
  or (_41329_, _39748_, _39741_);
  and (_39749_, _39375_, _33466_);
  nand (_39750_, _39749_, _29154_);
  or (_39751_, _39749_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39752_, _39751_, _29231_);
  and (_39753_, _39752_, _39750_);
  nor (_39754_, _39458_, _38479_);
  and (_39755_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39756_, _39755_, _39754_);
  and (_39757_, _39756_, _28573_);
  and (_39758_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39759_, _39758_, rst);
  or (_39760_, _39759_, _39757_);
  or (_41331_, _39760_, _39753_);
  and (_39765_, _39375_, _34196_);
  nand (_39766_, _39765_, _29154_);
  or (_39767_, _39765_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39768_, _39767_, _29231_);
  and (_39769_, _39768_, _39766_);
  nor (_39770_, _39458_, _38472_);
  and (_39771_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39772_, _39771_, _39770_);
  and (_39773_, _39772_, _28573_);
  and (_39774_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39775_, _39774_, rst);
  or (_39776_, _39775_, _39773_);
  or (_41333_, _39776_, _39769_);
  and (_39777_, _39466_, _24906_);
  nand (_39778_, _39777_, _29154_);
  or (_39779_, _39777_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39780_, _39779_, _29231_);
  and (_39781_, _39780_, _39778_);
  and (_39782_, _39474_, _38519_);
  and (_39783_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_39784_, _39783_, _39782_);
  and (_39785_, _39784_, _28573_);
  and (_39786_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_39787_, _39786_, rst);
  or (_39788_, _39787_, _39785_);
  or (_41335_, _39788_, _39781_);
  and (_39789_, _39466_, _38451_);
  nand (_39790_, _39789_, _29154_);
  or (_39791_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39792_, _39791_, _29231_);
  and (_39793_, _39792_, _39790_);
  nor (_39794_, _39475_, _38509_);
  and (_39795_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39796_, _39795_, _39794_);
  and (_39797_, _39796_, _28573_);
  and (_39798_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39799_, _39798_, rst);
  or (_39800_, _39799_, _39797_);
  or (_41337_, _39800_, _39793_);
  and (_39801_, _39466_, _31200_);
  nand (_39802_, _39801_, _29154_);
  or (_39803_, _39801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39804_, _39803_, _29231_);
  and (_39805_, _39804_, _39802_);
  nor (_39806_, _39475_, _38502_);
  and (_39807_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39808_, _39807_, _39806_);
  and (_39809_, _39808_, _28573_);
  and (_39810_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39811_, _39810_, rst);
  or (_39812_, _39811_, _39809_);
  or (_41338_, _39812_, _39805_);
  and (_39813_, _39466_, _31921_);
  nand (_39814_, _39813_, _29154_);
  or (_39815_, _39813_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39816_, _39815_, _29231_);
  and (_39817_, _39816_, _39814_);
  nor (_39818_, _39475_, _38494_);
  and (_39819_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39820_, _39819_, _39818_);
  and (_39821_, _39820_, _28573_);
  and (_39822_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39823_, _39822_, rst);
  or (_39824_, _39823_, _39821_);
  or (_41340_, _39824_, _39817_);
  and (_39827_, _39466_, _32683_);
  nand (_39833_, _39827_, _29154_);
  or (_39834_, _39827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39835_, _39834_, _29231_);
  and (_39836_, _39835_, _39833_);
  nor (_39837_, _39475_, _38486_);
  and (_39838_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39839_, _39838_, _39837_);
  and (_39840_, _39839_, _28573_);
  and (_39841_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39842_, _39841_, rst);
  or (_39843_, _39842_, _39840_);
  or (_41342_, _39843_, _39836_);
  and (_39844_, _39466_, _33466_);
  nand (_39845_, _39844_, _29154_);
  or (_39846_, _39844_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39847_, _39846_, _29231_);
  and (_39848_, _39847_, _39845_);
  nor (_39849_, _39475_, _38479_);
  and (_39850_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39851_, _39850_, _39849_);
  and (_39852_, _39851_, _28573_);
  and (_39853_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39854_, _39853_, rst);
  or (_39855_, _39854_, _39852_);
  or (_41344_, _39855_, _39848_);
  and (_39856_, _39466_, _34196_);
  nand (_39857_, _39856_, _29154_);
  or (_39858_, _39856_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39859_, _39858_, _29231_);
  and (_39860_, _39859_, _39857_);
  nor (_39861_, _39475_, _38472_);
  and (_39862_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39863_, _39862_, _39861_);
  and (_39864_, _39863_, _28573_);
  and (_39865_, _39234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39866_, _39865_, rst);
  or (_39867_, _39866_, _39864_);
  or (_41345_, _39867_, _39860_);
  nor (_39868_, _25722_, _25548_);
  and (_39869_, _39868_, _39353_);
  and (_39870_, _39869_, _38957_);
  and (_39871_, _39870_, _29187_);
  nand (_39872_, _39871_, _29154_);
  and (_39873_, _38931_, _25558_);
  and (_39874_, _39873_, _39473_);
  not (_39875_, _39874_);
  or (_39877_, _39871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_39881_, _39877_, _39875_);
  and (_39882_, _39881_, _39872_);
  nor (_39883_, _39875_, _38540_);
  or (_39884_, _39883_, _39882_);
  and (_41836_, _39884_, _41894_);
  and (_39885_, _25722_, _25558_);
  and (_39886_, _39885_, _38957_);
  and (_39887_, _39886_, _39353_);
  and (_39888_, _39887_, _29187_);
  nand (_39889_, _39888_, _29154_);
  and (_39890_, _39873_, _39441_);
  not (_39891_, _39890_);
  or (_39892_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_39893_, _39892_, _39891_);
  and (_39894_, _39893_, _39889_);
  nor (_39898_, _39891_, _38540_);
  or (_39905_, _39898_, _39894_);
  and (_41839_, _39905_, _41894_);
  or (_39906_, _24895_, _31189_);
  and (_39907_, _39906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39908_, _39907_, _39099_);
  and (_39909_, _39886_, _38432_);
  and (_39910_, _39909_, _39908_);
  and (_39911_, _39873_, _38450_);
  nand (_39912_, _39909_, _24884_);
  and (_39913_, _39912_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39914_, _39913_, _39911_);
  or (_39915_, _39914_, _39910_);
  nand (_39916_, _39911_, _38472_);
  and (_39917_, _39916_, _41894_);
  and (_41841_, _39917_, _39915_);
  and (_39918_, _29231_, _29176_);
  nor (_39919_, _24644_, _25548_);
  and (_39920_, _39919_, _38450_);
  and (_39921_, _39920_, _39918_);
  nand (_39922_, _39921_, _29154_);
  not (_39923_, _39911_);
  not (_39924_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_39925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_39926_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_39927_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _39926_);
  and (_39928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39929_, _39928_, _39927_);
  nor (_39930_, _39929_, _39925_);
  or (_39931_, _39930_, _39924_);
  and (_39932_, _39926_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_39933_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_39934_, _39933_, _39932_);
  nor (_39935_, _39934_, _39925_);
  and (_39936_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _39926_);
  and (_39937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39938_, _39937_, _39936_);
  nand (_39939_, _39938_, _39935_);
  or (_39940_, _39939_, _39931_);
  and (_39941_, _39940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_39942_, _39941_, _39921_);
  and (_39943_, _39942_, _39923_);
  and (_39944_, _39943_, _39922_);
  nor (_39945_, _39923_, _38540_);
  or (_39946_, _39945_, _39944_);
  and (_41844_, _39946_, _41894_);
  and (_39947_, _29231_, _30479_);
  and (_39948_, _39947_, _39920_);
  nand (_39949_, _39948_, _29154_);
  nor (_39950_, _39938_, _39925_);
  nand (_39951_, _39950_, _39934_);
  or (_39952_, _39951_, _39931_);
  and (_39953_, _39952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_39954_, _39953_, _39948_);
  and (_39955_, _39954_, _39923_);
  and (_39956_, _39955_, _39949_);
  nor (_39957_, _39923_, _38479_);
  or (_39958_, _39957_, _39956_);
  and (_41845_, _39958_, _41894_);
  nor (_39959_, _29165_, _25548_);
  and (_39960_, _39959_, _38450_);
  and (_39961_, _39960_, _39947_);
  nand (_39962_, _39961_, _29154_);
  not (_39963_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_39964_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _39963_);
  nand (_39965_, _39930_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_39966_, _39950_, _39935_);
  or (_39967_, _39966_, _39965_);
  and (_39968_, _39967_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_39969_, _39968_, _39964_);
  or (_39970_, _39969_, _39961_);
  and (_39971_, _39970_, _39923_);
  and (_39972_, _39971_, _39962_);
  nor (_39973_, _39923_, _38509_);
  or (_39974_, _39973_, _39972_);
  and (_41847_, _39974_, _41894_);
  and (_39975_, _39960_, _39918_);
  nand (_39976_, _39975_, _29154_);
  and (_39977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_39978_, _39965_, _39951_);
  and (_39979_, _39978_, _39977_);
  or (_39980_, _39979_, _39975_);
  and (_39981_, _39980_, _39923_);
  and (_39982_, _39981_, _39976_);
  nor (_39983_, _39923_, _38494_);
  or (_39984_, _39983_, _39982_);
  and (_41849_, _39984_, _41894_);
  and (_39985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_39986_, _39985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_39987_, _39986_);
  and (_39988_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_39989_, _39988_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_39990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_39991_, _39990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_39992_, _39991_, _39989_);
  and (_39993_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_39994_, _39993_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  not (_39995_, _39994_);
  and (_39996_, _39995_, _39992_);
  and (_39997_, _39996_, _39987_);
  not (_39998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_39999_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40000_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _39926_);
  or (_40001_, _40000_, _39999_);
  nor (_40002_, _40001_, _39998_);
  nor (_40003_, _40002_, _39925_);
  nor (_40004_, _40003_, _39997_);
  and (_40005_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_40006_, _40005_, _39926_);
  and (_40007_, _40006_, _40004_);
  and (_40008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _39925_);
  not (_40009_, _40008_);
  not (_40010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40011_, _39988_, _40010_);
  not (_40012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40013_, _39990_, _40012_);
  nor (_40014_, _40013_, _40011_);
  not (_40015_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40016_, _39993_, _40015_);
  not (_40017_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40018_, _39985_, _40017_);
  nor (_40019_, _40018_, _40016_);
  and (_40020_, _40019_, _40014_);
  nor (_40021_, _40020_, _40009_);
  nand (_40022_, _40021_, _40006_);
  and (_40023_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41894_);
  nand (_40024_, _40023_, _40022_);
  nor (_41881_, _40024_, _40007_);
  nor (_40025_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40026_, _40025_);
  nor (_40027_, _40021_, _40004_);
  nor (_40028_, _40027_, _40026_);
  nand (_40029_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41894_);
  nor (_41883_, _40029_, _40028_);
  and (_40030_, _39986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40031_, _39992_);
  or (_40032_, _40031_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_40033_, _40032_, _40030_);
  or (_40034_, _39996_, _39932_);
  and (_40035_, _40034_, _40033_);
  and (_40036_, _40035_, _40004_);
  or (_40037_, _40036_, _40005_);
  and (_40038_, _40027_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_40039_, _40004_);
  and (_40040_, _40021_, _40039_);
  and (_40041_, _40018_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40042_, _40041_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_40043_, _40014_);
  and (_40044_, _40016_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40045_, _40044_, _40043_);
  and (_40046_, _40045_, _40042_);
  and (_40047_, _40043_, _39932_);
  or (_40048_, _40047_, _40046_);
  and (_40049_, _40048_, _40040_);
  or (_40050_, _40049_, _40038_);
  or (_40051_, _40050_, _40037_);
  not (_40052_, _40005_);
  or (_40053_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40054_, _40053_, _41894_);
  and (_41885_, _40054_, _40051_);
  and (_40055_, _39986_, _39926_);
  or (_40056_, _40031_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_40057_, _40056_, _40055_);
  or (_40058_, _39996_, _39933_);
  and (_40059_, _40058_, _40057_);
  and (_40060_, _40059_, _40004_);
  or (_40061_, _40060_, _40005_);
  and (_40062_, _40027_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40063_, _40018_, _39926_);
  or (_40064_, _40063_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40065_, _40016_, _39926_);
  nor (_40066_, _40065_, _40043_);
  and (_40067_, _40066_, _40064_);
  and (_40068_, _40043_, _39933_);
  or (_40069_, _40068_, _40067_);
  and (_40070_, _40069_, _40040_);
  or (_40071_, _40070_, _40062_);
  or (_40072_, _40071_, _40061_);
  or (_40073_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40074_, _40073_, _41894_);
  and (_41886_, _40074_, _40072_);
  nand (_40075_, _40027_, _39925_);
  nor (_40076_, _39926_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_40077_, _40076_, _40005_);
  and (_40078_, _40077_, _41894_);
  and (_41888_, _40078_, _40075_);
  and (_40079_, _40027_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_40080_, _39926_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_40081_, _40080_, _40076_);
  nor (_40082_, _40081_, _40039_);
  or (_40083_, _40082_, _40005_);
  or (_40084_, _40083_, _40079_);
  or (_40085_, _40081_, _40052_);
  and (_40086_, _40085_, _41894_);
  and (_41890_, _40086_, _40084_);
  and (_40087_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41894_);
  and (_41892_, _40087_, _40005_);
  nor (_40088_, _40027_, _40005_);
  and (_40089_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_40090_, _40089_, _40088_);
  and (_42811_, _40090_, _41894_);
  and (_40091_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_40092_, _40091_, _40088_);
  and (_42813_, _40092_, _41894_);
  and (_40093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _41894_);
  and (_42815_, _40093_, _40005_);
  not (_40094_, _40011_);
  nor (_40095_, _40018_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_40096_, _40095_, _40016_);
  or (_40097_, _40096_, _40013_);
  and (_40098_, _40097_, _40094_);
  and (_40099_, _40098_, _40040_);
  not (_40100_, _39989_);
  or (_40101_, _39986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40102_, _40101_, _39995_);
  or (_40103_, _40102_, _39991_);
  and (_40104_, _40103_, _40100_);
  and (_40105_, _40104_, _40004_);
  or (_40106_, _40105_, _40005_);
  or (_40107_, _40106_, _40099_);
  or (_40108_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40109_, _40108_, _41894_);
  and (_42817_, _40109_, _40107_);
  nand (_40110_, _40014_, _40008_);
  nor (_40111_, _40110_, _40019_);
  or (_40112_, _40111_, _40004_);
  nand (_40113_, _40004_, _40031_);
  and (_40114_, _40113_, _40112_);
  or (_40115_, _40114_, _40005_);
  or (_40116_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_40117_, _40116_, _41894_);
  and (_42818_, _40117_, _40115_);
  and (_40118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _41894_);
  and (_42820_, _40118_, _40005_);
  and (_40119_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _41894_);
  and (_42822_, _40119_, _40005_);
  nand (_40120_, _40027_, _40025_);
  nor (_40121_, _40005_, _40004_);
  or (_40122_, _40121_, _39926_);
  and (_40123_, _40122_, _41894_);
  and (_42824_, _40123_, _40120_);
  not (_40124_, _40088_);
  and (_40125_, _40124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_40126_, _40055_);
  and (_40127_, _40126_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_40128_, _39994_, _39926_);
  or (_40129_, _40128_, _39991_);
  or (_40130_, _40129_, _40127_);
  not (_40131_, _39991_);
  or (_40132_, _40131_, _39928_);
  and (_40133_, _40132_, _40130_);
  or (_40134_, _40133_, _39989_);
  or (_40135_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _39926_);
  or (_40136_, _40135_, _40100_);
  and (_40137_, _40136_, _40004_);
  and (_40138_, _40137_, _40134_);
  not (_40139_, _40063_);
  and (_40140_, _40139_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_40141_, _40065_, _40013_);
  or (_40142_, _40141_, _40140_);
  not (_40143_, _40013_);
  or (_40144_, _40143_, _39928_);
  and (_40145_, _40144_, _40094_);
  and (_40146_, _40145_, _40142_);
  and (_40147_, _40135_, _40011_);
  or (_40148_, _40147_, _40146_);
  and (_40149_, _40148_, _40040_);
  or (_40150_, _40149_, _40138_);
  and (_40151_, _40150_, _40052_);
  or (_40152_, _40151_, _40125_);
  and (_42826_, _40152_, _41894_);
  and (_40153_, _40124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40154_, _40126_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40155_, _40154_, _40129_);
  or (_40156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _39926_);
  or (_40157_, _40156_, _40131_);
  and (_40158_, _40157_, _40100_);
  and (_40159_, _40158_, _40155_);
  and (_40160_, _39989_, _39937_);
  or (_40161_, _40160_, _40159_);
  and (_40162_, _40161_, _40004_);
  and (_40163_, _40139_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40164_, _40163_, _40141_);
  or (_40165_, _40156_, _40143_);
  and (_40166_, _40165_, _40094_);
  and (_40167_, _40166_, _40164_);
  and (_40168_, _40011_, _39937_);
  or (_40169_, _40168_, _40167_);
  and (_40170_, _40169_, _40040_);
  or (_40171_, _40170_, _40162_);
  and (_40172_, _40171_, _40052_);
  or (_40173_, _40172_, _40153_);
  and (_42827_, _40173_, _41894_);
  and (_40174_, _40124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_40175_, _40030_);
  and (_40176_, _40175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_40177_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40178_, _40177_, _39991_);
  or (_40179_, _40178_, _40176_);
  or (_40180_, _40131_, _39927_);
  and (_40181_, _40180_, _40179_);
  or (_40182_, _40181_, _39989_);
  or (_40183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40184_, _40183_, _40100_);
  and (_40185_, _40184_, _40004_);
  and (_40186_, _40185_, _40182_);
  not (_40187_, _40041_);
  and (_40188_, _40187_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_40189_, _40044_, _40013_);
  or (_40190_, _40189_, _40188_);
  or (_40191_, _40143_, _39927_);
  and (_40192_, _40191_, _40094_);
  and (_40193_, _40192_, _40190_);
  and (_40194_, _40183_, _40011_);
  or (_40195_, _40194_, _40193_);
  and (_40196_, _40195_, _40040_);
  or (_40197_, _40196_, _40186_);
  and (_40198_, _40197_, _40052_);
  or (_40199_, _40198_, _40174_);
  and (_42829_, _40199_, _41894_);
  and (_40200_, _40124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40201_, _40175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40202_, _40201_, _40178_);
  or (_40203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40204_, _40203_, _40131_);
  and (_40205_, _40204_, _40100_);
  and (_40206_, _40205_, _40202_);
  and (_40207_, _39989_, _39936_);
  or (_40208_, _40207_, _40206_);
  and (_40209_, _40208_, _40004_);
  and (_40210_, _40187_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40211_, _40210_, _40189_);
  or (_40212_, _40203_, _40143_);
  and (_40213_, _40212_, _40094_);
  and (_40214_, _40213_, _40211_);
  and (_40215_, _40011_, _39936_);
  or (_40216_, _40215_, _40214_);
  and (_40217_, _40216_, _40040_);
  or (_40218_, _40217_, _40209_);
  and (_40219_, _40218_, _40052_);
  or (_40220_, _40219_, _40200_);
  and (_42831_, _40220_, _41894_);
  and (_40221_, _40025_, _40004_);
  nand (_40222_, _40025_, _40021_);
  and (_40223_, _40222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_40224_, _40223_, _40221_);
  and (_42833_, _40224_, _41894_);
  and (_40225_, _40022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_40226_, _40225_, _40007_);
  and (_42835_, _40226_, _41894_);
  and (_40227_, _39909_, _24906_);
  or (_40228_, _40227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_40229_, _40228_, _39923_);
  nand (_40230_, _40227_, _29154_);
  and (_40231_, _40230_, _40229_);
  and (_40232_, _39911_, _38519_);
  or (_40233_, _40232_, _40231_);
  and (_42837_, _40233_, _41894_);
  and (_40234_, _39909_, _31200_);
  nand (_40235_, _40234_, _29154_);
  or (_40236_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_40237_, _40236_, _39923_);
  and (_40238_, _40237_, _40235_);
  nor (_40239_, _39923_, _38502_);
  or (_40240_, _40239_, _40238_);
  and (_42839_, _40240_, _41894_);
  and (_40241_, _39909_, _32683_);
  nand (_40242_, _40241_, _29154_);
  or (_40243_, _40241_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_40244_, _40243_, _39923_);
  and (_40245_, _40244_, _40242_);
  nor (_40246_, _39923_, _38486_);
  or (_40247_, _40246_, _40245_);
  and (_42841_, _40247_, _41894_);
  and (_40248_, _39887_, _24906_);
  nand (_40249_, _40248_, _29154_);
  or (_40250_, _40248_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40251_, _40250_, _39891_);
  and (_40252_, _40251_, _40249_);
  and (_40253_, _39890_, _38519_);
  or (_40254_, _40253_, _40252_);
  and (_42843_, _40254_, _41894_);
  and (_40255_, _39887_, _38451_);
  nand (_40256_, _40255_, _29154_);
  or (_40257_, _40255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40258_, _40257_, _40256_);
  or (_40259_, _40258_, _39890_);
  nand (_40260_, _39890_, _38509_);
  and (_40261_, _40260_, _41894_);
  and (_42844_, _40261_, _40259_);
  and (_40262_, _31233_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40263_, _40262_, _31222_);
  and (_40264_, _40263_, _39887_);
  nand (_40265_, _39887_, _39506_);
  and (_40266_, _40265_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40267_, _40266_, _39890_);
  or (_40268_, _40267_, _40264_);
  nand (_40269_, _39890_, _38502_);
  and (_40270_, _40269_, _41894_);
  and (_42846_, _40270_, _40268_);
  and (_40271_, _39887_, _31921_);
  nand (_40272_, _40271_, _29154_);
  or (_40273_, _40271_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40274_, _40273_, _39891_);
  and (_40275_, _40274_, _40272_);
  nor (_40276_, _39891_, _38494_);
  or (_40277_, _40276_, _40275_);
  and (_42848_, _40277_, _41894_);
  and (_40278_, _39887_, _32683_);
  nand (_40279_, _40278_, _29154_);
  or (_40280_, _40278_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_40281_, _40280_, _39891_);
  and (_40282_, _40281_, _40279_);
  nor (_40283_, _39891_, _38486_);
  or (_40284_, _40283_, _40282_);
  and (_42850_, _40284_, _41894_);
  and (_40285_, _39887_, _33466_);
  nand (_40286_, _40285_, _29154_);
  or (_40287_, _40285_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_40288_, _40287_, _39891_);
  and (_40289_, _40288_, _40286_);
  nor (_40290_, _39891_, _38479_);
  or (_40291_, _40290_, _40289_);
  and (_42852_, _40291_, _41894_);
  and (_40292_, _39887_, _34196_);
  nand (_40293_, _40292_, _29154_);
  or (_40294_, _40292_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_40295_, _40294_, _39891_);
  and (_40296_, _40295_, _40293_);
  nor (_40297_, _39891_, _38472_);
  or (_40298_, _40297_, _40296_);
  and (_42854_, _40298_, _41894_);
  and (_40299_, _39870_, _24906_);
  nand (_40300_, _40299_, _29154_);
  or (_40301_, _40299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40302_, _40301_, _39875_);
  and (_40303_, _40302_, _40300_);
  and (_40304_, _39874_, _38519_);
  or (_40305_, _40304_, _40303_);
  and (_42856_, _40305_, _41894_);
  and (_40306_, _39870_, _38451_);
  nand (_40307_, _40306_, _29154_);
  or (_40308_, _40306_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40309_, _40308_, _39875_);
  and (_40310_, _40309_, _40307_);
  nor (_40311_, _39875_, _38509_);
  or (_40312_, _40311_, _40310_);
  and (_42858_, _40312_, _41894_);
  and (_40313_, _31233_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40314_, _40313_, _31222_);
  and (_40315_, _40314_, _39870_);
  nand (_40316_, _39870_, _39506_);
  and (_40317_, _40316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40318_, _40317_, _39874_);
  or (_40319_, _40318_, _40315_);
  nand (_40320_, _39874_, _38502_);
  and (_40321_, _40320_, _41894_);
  and (_42860_, _40321_, _40319_);
  and (_40322_, _39870_, _31921_);
  nand (_40323_, _40322_, _29154_);
  or (_40324_, _40322_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40325_, _40324_, _39875_);
  and (_40326_, _40325_, _40323_);
  nor (_40327_, _39875_, _38494_);
  or (_40328_, _40327_, _40326_);
  and (_42862_, _40328_, _41894_);
  and (_40329_, _39870_, _32683_);
  nand (_40330_, _40329_, _29154_);
  or (_40331_, _40329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40332_, _40331_, _40330_);
  or (_40333_, _40332_, _39874_);
  nand (_40334_, _39874_, _38486_);
  and (_40335_, _40334_, _41894_);
  and (_42864_, _40335_, _40333_);
  and (_40336_, _39870_, _33466_);
  nand (_40337_, _40336_, _29154_);
  or (_40338_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40339_, _40338_, _39875_);
  and (_40340_, _40339_, _40337_);
  nor (_40341_, _39875_, _38479_);
  or (_40342_, _40341_, _40340_);
  and (_42866_, _40342_, _41894_);
  and (_40343_, _39870_, _34196_);
  nand (_40344_, _40343_, _29154_);
  or (_40345_, _40343_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_40346_, _40345_, _40344_);
  or (_40347_, _40346_, _39874_);
  nand (_40348_, _39874_, _38472_);
  and (_40349_, _40348_, _41894_);
  and (_42868_, _40349_, _40347_);
  and (_40350_, _38542_, _38411_);
  not (_40351_, _40350_);
  not (_40352_, _38389_);
  and (_40353_, _40352_, _37984_);
  and (_40354_, _40353_, _36960_);
  not (_40355_, _38540_);
  and (_40356_, _35808_, _30468_);
  nor (_40357_, _35808_, _30468_);
  not (_40358_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_40359_, _28540_, _40358_);
  and (_40360_, _40359_, _31233_);
  nand (_40361_, _40360_, _25395_);
  or (_40362_, _40361_, _40357_);
  nor (_40363_, _40362_, _40356_);
  nor (_40364_, _38935_, _39033_);
  nor (_40365_, _40364_, _39062_);
  and (_40366_, _40365_, _25558_);
  nor (_40367_, _40365_, _25558_);
  nor (_40368_, _40367_, _40366_);
  and (_40369_, _40368_, _40363_);
  and (_40370_, _40369_, _40355_);
  and (_40371_, _40365_, _35819_);
  and (_40372_, _40371_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_40373_, _40365_, _35819_);
  and (_40374_, _40373_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_40375_, _40374_, _40372_);
  nor (_40376_, _40365_, _35808_);
  and (_40377_, _40376_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_40378_, _40365_, _35808_);
  and (_40379_, _40378_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_40380_, _40379_, _40377_);
  and (_40381_, _40380_, _40375_);
  nor (_40382_, _40381_, _40369_);
  nor (_40383_, _40382_, _40370_);
  not (_40384_, _40383_);
  and (_40385_, _40384_, _40354_);
  not (_40386_, _40385_);
  not (_40387_, _36960_);
  nor (_40388_, _40352_, _37984_);
  not (_40389_, _34358_);
  and (_40390_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_40391_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_40392_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_40393_, _40392_, _40391_);
  and (_40394_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_40395_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_40396_, _40395_, _40394_);
  and (_40397_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_40398_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_40399_, _40398_, _40397_);
  and (_40400_, _40399_, _40396_);
  and (_40401_, _40400_, _40393_);
  and (_40402_, _35830_, _34358_);
  not (_40403_, _40402_);
  nor (_40404_, _40403_, _40401_);
  nor (_40405_, _40404_, _40390_);
  not (_40406_, _40405_);
  and (_40407_, _40406_, _40388_);
  nor (_40408_, _40407_, _40387_);
  and (_40409_, _40408_, _40386_);
  and (_40410_, _40409_, _40351_);
  not (_40411_, _37450_);
  and (_40412_, _37604_, _40411_);
  and (_40413_, _35566_, _36807_);
  nor (_40414_, _40413_, _37615_);
  and (_40415_, _36807_, _37058_);
  nor (_40416_, _40415_, _37742_);
  and (_40417_, _40416_, _40414_);
  and (_40418_, _37797_, _37731_);
  and (_40419_, _40418_, _40417_);
  and (_40420_, _40419_, _40412_);
  nor (_40421_, _40420_, _34314_);
  and (_40422_, _37698_, _36807_);
  nor (_40423_, _37863_, _40422_);
  nor (_40424_, _37885_, _40423_);
  nor (_40425_, _40424_, _40421_);
  not (_40426_, _40425_);
  and (_40427_, _40426_, _40410_);
  and (_40428_, _40388_, _36960_);
  and (_40429_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_40430_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_40431_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_40432_, _40431_, _40430_);
  and (_40433_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_40434_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_40435_, _40434_, _40433_);
  and (_40436_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_40437_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_40438_, _40437_, _40436_);
  and (_40439_, _40438_, _40435_);
  and (_40440_, _40439_, _40432_);
  nor (_40441_, _40440_, _40403_);
  nor (_40442_, _40441_, _40429_);
  not (_40443_, _40442_);
  and (_40444_, _40443_, _40428_);
  not (_40445_, _40444_);
  and (_40446_, _40387_, _38389_);
  and (_40447_, _40446_, _37984_);
  not (_40448_, _38580_);
  and (_40449_, _40448_, _38411_);
  nor (_40450_, _40449_, _40447_);
  and (_40451_, _40450_, _40445_);
  and (_40452_, _38400_, _40387_);
  and (_40453_, _40376_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  not (_40454_, _40453_);
  and (_40455_, _40373_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_40456_, _40371_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_40457_, _40456_, _40455_);
  and (_40458_, _40457_, _40454_);
  and (_40459_, _40378_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_40460_, _40459_, _40369_);
  and (_40461_, _40460_, _40458_);
  and (_40462_, _40369_, _38479_);
  or (_40463_, _40462_, _40461_);
  not (_40464_, _40463_);
  and (_40465_, _40464_, _40354_);
  nor (_40466_, _40465_, _40452_);
  and (_40467_, _40466_, _40451_);
  not (_40468_, _40467_);
  and (_40469_, _40468_, _40427_);
  not (_40470_, _38562_);
  and (_40471_, _40470_, _38411_);
  and (_40472_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_40473_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_40474_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_40475_, _40474_, _40473_);
  and (_40476_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_40477_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_40478_, _40477_, _40476_);
  and (_40479_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_40480_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_40481_, _40480_, _40479_);
  and (_40482_, _40481_, _40478_);
  and (_40483_, _40482_, _40475_);
  nor (_40484_, _40483_, _40403_);
  nor (_40485_, _40484_, _40472_);
  not (_40486_, _40485_);
  and (_40487_, _40486_, _40428_);
  nor (_40488_, _40487_, _40471_);
  and (_40489_, _38389_, _37984_);
  and (_40490_, _40489_, _36960_);
  and (_40491_, _40490_, _36862_);
  not (_40492_, _40369_);
  nor (_40493_, _40492_, _38502_);
  and (_40494_, _40371_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_40495_, _40373_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_40496_, _40495_, _40494_);
  and (_40497_, _40376_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_40498_, _40378_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_40499_, _40498_, _40497_);
  and (_40500_, _40499_, _40496_);
  nor (_40501_, _40500_, _40369_);
  nor (_40502_, _40501_, _40493_);
  not (_40503_, _40502_);
  and (_40504_, _40503_, _40354_);
  nor (_40505_, _40504_, _40491_);
  and (_40506_, _40505_, _40488_);
  nor (_40507_, _40506_, _40426_);
  nor (_40508_, _40507_, _40469_);
  and (_40509_, _25395_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40510_, _40509_, _39112_);
  nor (_40511_, _24644_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40512_, _40511_, _40510_);
  not (_40513_, _40512_);
  and (_40514_, _40513_, _40508_);
  not (_40515_, _38568_);
  and (_40516_, _40515_, _38411_);
  and (_40517_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_40518_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_40519_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_40520_, _40519_, _40518_);
  and (_40521_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_40522_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_40523_, _40522_, _40521_);
  and (_40524_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_40525_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_40526_, _40525_, _40524_);
  and (_40527_, _40526_, _40523_);
  and (_40528_, _40527_, _40520_);
  nor (_40529_, _40528_, _40403_);
  nor (_40530_, _40529_, _40517_);
  not (_40531_, _40530_);
  and (_40532_, _40531_, _40428_);
  nor (_40533_, _40532_, _40516_);
  not (_40534_, _40365_);
  and (_40535_, _40490_, _40534_);
  and (_40536_, _40373_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_40537_, _40371_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_40538_, _40537_, _40536_);
  and (_40539_, _40378_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  not (_40540_, _40539_);
  and (_40541_, _40540_, _40538_);
  and (_40542_, _40376_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_40543_, _40542_, _40369_);
  and (_40544_, _40543_, _40541_);
  and (_40545_, _40369_, _38494_);
  or (_40546_, _40545_, _40544_);
  not (_40547_, _40546_);
  and (_40548_, _40547_, _40354_);
  nor (_40549_, _40548_, _40535_);
  and (_40550_, _40549_, _40533_);
  not (_40551_, _40550_);
  and (_40552_, _40551_, _40427_);
  not (_40553_, _38550_);
  and (_40554_, _40553_, _38411_);
  and (_40555_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_40556_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_40557_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_40558_, _40557_, _40556_);
  and (_40559_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_40560_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_40561_, _40560_, _40559_);
  and (_40562_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_40563_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_40564_, _40563_, _40562_);
  and (_40565_, _40564_, _40561_);
  and (_40566_, _40565_, _40558_);
  nor (_40567_, _40566_, _40403_);
  nor (_40568_, _40567_, _40555_);
  not (_40569_, _40568_);
  and (_40570_, _40569_, _40428_);
  nor (_40571_, _40570_, _40554_);
  and (_40572_, _40490_, _35819_);
  and (_40573_, _40371_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_40574_, _40373_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_40575_, _40574_, _40573_);
  and (_40576_, _40376_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_40577_, _40378_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_40578_, _40577_, _40576_);
  and (_40579_, _40578_, _40575_);
  nor (_40580_, _40579_, _40369_);
  and (_40581_, _40369_, _38519_);
  nor (_40582_, _40581_, _40580_);
  not (_40583_, _40582_);
  and (_40584_, _40583_, _40354_);
  nor (_40585_, _40584_, _40572_);
  and (_40586_, _40585_, _40571_);
  nor (_40587_, _40586_, _40426_);
  nor (_40588_, _40587_, _40552_);
  and (_40589_, _40509_, _25558_);
  nor (_40590_, _24884_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40591_, _40590_, _40589_);
  not (_40592_, _40591_);
  nor (_40593_, _40592_, _40588_);
  nor (_40594_, _40593_, _40514_);
  nor (_40595_, _40513_, _40508_);
  not (_40596_, _40595_);
  nor (_40597_, _40551_, _40427_);
  not (_40598_, _38472_);
  and (_40599_, _40369_, _40598_);
  and (_40600_, _40371_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_40601_, _40373_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_40602_, _40601_, _40600_);
  and (_40603_, _40376_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_40604_, _40378_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_40605_, _40604_, _40603_);
  and (_40606_, _40605_, _40602_);
  nor (_40607_, _40606_, _40369_);
  nor (_40608_, _40607_, _40599_);
  not (_40609_, _40608_);
  and (_40610_, _40609_, _40354_);
  and (_40611_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_40612_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_40613_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_40614_, _40613_, _40612_);
  and (_40615_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_40616_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_40617_, _40616_, _40615_);
  and (_40618_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_40619_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_40620_, _40619_, _40618_);
  and (_40621_, _40620_, _40617_);
  and (_40622_, _40621_, _40614_);
  nor (_40623_, _40622_, _40403_);
  nor (_40624_, _40623_, _40611_);
  not (_40625_, _40624_);
  and (_40626_, _40625_, _40388_);
  nor (_40627_, _40626_, _40610_);
  nor (_40628_, _40353_, _36960_);
  not (_40629_, _38586_);
  and (_40630_, _40629_, _38411_);
  nor (_40631_, _40630_, _40628_);
  and (_40632_, _40631_, _40627_);
  and (_40633_, _40632_, _40427_);
  nor (_40634_, _40633_, _40597_);
  nor (_40635_, _40509_, _25558_);
  and (_40636_, _40509_, _25122_);
  nor (_40637_, _40636_, _40635_);
  not (_40638_, _40637_);
  and (_40639_, _40638_, _40634_);
  nor (_40640_, _40638_, _40634_);
  nor (_40641_, _40640_, _40639_);
  and (_40642_, _40641_, _40596_);
  not (_40643_, _38574_);
  and (_40644_, _40643_, _38411_);
  nor (_40645_, _40644_, _40446_);
  and (_40646_, _38953_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_40647_, _40646_, _39079_);
  not (_40648_, _40647_);
  and (_40649_, _40648_, _40490_);
  and (_40650_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_40651_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_40652_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_40653_, _40652_, _40651_);
  and (_40654_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_40655_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_40656_, _40655_, _40654_);
  and (_40657_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_40658_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_40659_, _40658_, _40657_);
  and (_40660_, _40659_, _40656_);
  and (_40661_, _40660_, _40653_);
  nor (_40662_, _40661_, _40403_);
  nor (_40663_, _40662_, _40650_);
  not (_40664_, _40663_);
  and (_40665_, _40664_, _40428_);
  and (_40666_, _40378_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_40667_, _40373_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_40668_, _40667_, _40666_);
  and (_40669_, _40376_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_40670_, _40371_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_40671_, _40670_, _40669_);
  and (_40672_, _40671_, _40668_);
  and (_40673_, _40672_, _40492_);
  and (_40674_, _40369_, _38486_);
  nor (_40675_, _40674_, _40673_);
  and (_40676_, _40675_, _40354_);
  or (_40677_, _40676_, _40665_);
  nor (_40678_, _40677_, _40649_);
  and (_40682_, _40678_, _40645_);
  not (_40688_, _40682_);
  and (_40694_, _40688_, _40427_);
  and (_40700_, _40353_, _40387_);
  not (_40706_, _38556_);
  and (_40711_, _40706_, _38411_);
  nor (_40712_, _40711_, _40700_);
  not (_40713_, _36083_);
  and (_40714_, _40490_, _40713_);
  and (_40715_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_40716_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_40717_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_40718_, _40717_, _40716_);
  and (_40719_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_40720_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_40721_, _40720_, _40719_);
  and (_40722_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_40723_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_40724_, _40723_, _40722_);
  and (_40725_, _40724_, _40721_);
  and (_40728_, _40725_, _40718_);
  nor (_40732_, _40728_, _40403_);
  nor (_40736_, _40732_, _40715_);
  not (_40737_, _40736_);
  and (_40738_, _40737_, _40428_);
  and (_40739_, _40371_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_40744_, _40373_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_40749_, _40744_, _40739_);
  and (_40750_, _40376_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_40751_, _40378_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_40753_, _40751_, _40750_);
  and (_40759_, _40753_, _40749_);
  nor (_40762_, _40759_, _40369_);
  and (_40763_, _40369_, _38510_);
  nor (_40764_, _40763_, _40762_);
  not (_40769_, _40764_);
  and (_40774_, _40769_, _40354_);
  or (_40775_, _40774_, _40738_);
  nor (_40776_, _40775_, _40714_);
  and (_40778_, _40776_, _40712_);
  nor (_40784_, _40778_, _40426_);
  nor (_40787_, _40784_, _40694_);
  and (_40788_, _40509_, _38443_);
  nor (_40789_, _24764_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40795_, _40789_, _40788_);
  nand (_40799_, _40795_, _40787_);
  or (_40800_, _40795_, _40787_);
  and (_40801_, _40800_, _40799_);
  not (_40807_, _40801_);
  nor (_40811_, _25395_, _24382_);
  nor (_40812_, _40811_, _28551_);
  not (_40813_, _40812_);
  and (_40818_, _40592_, _40588_);
  nor (_40823_, _40818_, _40813_);
  and (_40824_, _40823_, _40807_);
  and (_40825_, _40824_, _40642_);
  and (_40827_, _40825_, _40594_);
  not (_40833_, _40508_);
  and (_40836_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_40837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_40838_, _40588_, _40837_);
  or (_40844_, _40838_, _40836_);
  and (_40848_, _40844_, _40787_);
  not (_40849_, _40787_);
  not (_40850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_40856_, _40588_, _40850_);
  and (_40860_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_40861_, _40860_, _40856_);
  and (_40862_, _40861_, _40849_);
  or (_40867_, _40862_, _40848_);
  or (_40872_, _40867_, _40833_);
  not (_40873_, _40634_);
  and (_40874_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not (_40878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_40884_, _40588_, _40878_);
  or (_40885_, _40884_, _40874_);
  and (_40886_, _40885_, _40787_);
  not (_40889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_40895_, _40588_, _40889_);
  and (_40897_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_40898_, _40897_, _40895_);
  and (_40901_, _40898_, _40849_);
  or (_40907_, _40901_, _40886_);
  or (_40909_, _40907_, _40508_);
  and (_40910_, _40909_, _40873_);
  and (_40913_, _40910_, _40872_);
  not (_40919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_40920_, _40588_, _40919_);
  or (_40921_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_40922_, _40921_, _40920_);
  and (_40923_, _40922_, _40787_);
  or (_40924_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_40925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_40926_, _40588_, _40925_);
  and (_40927_, _40926_, _40924_);
  and (_40928_, _40927_, _40849_);
  or (_40929_, _40928_, _40923_);
  or (_40930_, _40929_, _40833_);
  not (_40931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_40932_, _40588_, _40931_);
  or (_40933_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_40934_, _40933_, _40932_);
  and (_40935_, _40934_, _40787_);
  or (_40936_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_40937_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_40938_, _40588_, _40937_);
  and (_40939_, _40938_, _40936_);
  and (_40940_, _40939_, _40849_);
  or (_40941_, _40940_, _40935_);
  or (_40942_, _40941_, _40508_);
  and (_40943_, _40942_, _40634_);
  and (_40944_, _40943_, _40930_);
  or (_40945_, _40944_, _40913_);
  or (_40946_, _40945_, _40827_);
  not (_40947_, _40827_);
  or (_40948_, _40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_40949_, _40948_, _41894_);
  and (_42947_, _40949_, _40946_);
  nor (_40950_, _40591_, _40813_);
  nor (_40951_, _40813_, _40795_);
  and (_40952_, _40951_, _40950_);
  and (_40953_, _40637_, _40812_);
  nor (_40954_, _40813_, _40512_);
  and (_40955_, _40954_, _40953_);
  and (_40956_, _40955_, _40952_);
  and (_40957_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_40958_, _40957_, _26631_);
  nor (_40959_, _40958_, _29154_);
  nand (_40960_, _26631_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40961_, _17933_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40962_, _40961_, _40960_);
  nor (_40963_, _38540_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_40964_, _40963_, _40962_);
  or (_40965_, _40964_, _40959_);
  and (_40966_, _40965_, _40812_);
  and (_40967_, _40966_, _40956_);
  not (_40968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_40969_, _40956_, _40968_);
  or (_42959_, _40969_, _40967_);
  nor (_40970_, _40954_, _40953_);
  nor (_40971_, _40951_, _40950_);
  and (_40972_, _40971_, _40812_);
  and (_40973_, _40972_, _40970_);
  and (_40974_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _26543_);
  and (_40975_, _40974_, _26598_);
  nand (_40976_, _40975_, _29154_);
  not (_40977_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40978_, _38518_, _40977_);
  or (_40979_, _16777_, _40977_);
  and (_40980_, _40979_, _40978_);
  or (_40981_, _40980_, _40975_);
  and (_40982_, _40981_, _40976_);
  and (_40983_, _40982_, _40973_);
  not (_40984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_40985_, _40973_, _40984_);
  or (_43214_, _40985_, _40983_);
  not (_40986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_40987_, _40973_, _40986_);
  nand (_40988_, _40974_, _26664_);
  nor (_40989_, _40988_, _29154_);
  nor (_40990_, _38509_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40991_, _40974_, _26554_);
  and (_40992_, _40974_, _26631_);
  or (_40993_, _40992_, _40957_);
  or (_40994_, _40993_, _40991_);
  and (_40995_, _40994_, _17759_);
  or (_40996_, _40995_, _40990_);
  or (_40997_, _40996_, _40989_);
  and (_40998_, _40997_, _40973_);
  or (_43220_, _40998_, _40987_);
  not (_40999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_41000_, _40973_, _40999_);
  nand (_41001_, _40974_, _26565_);
  nor (_41002_, _41001_, _29154_);
  nor (_41003_, _38502_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41004_, _40974_, _26653_);
  or (_41005_, _41004_, _40993_);
  and (_41006_, _41005_, _16414_);
  or (_41007_, _41006_, _41003_);
  or (_41008_, _41007_, _41002_);
  and (_41009_, _41008_, _40973_);
  or (_43226_, _41009_, _41000_);
  and (_41010_, _40992_, _29767_);
  nor (_41011_, _38494_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_41012_, _40991_, _40957_);
  or (_41013_, _41012_, _41004_);
  and (_41014_, _41013_, _17443_);
  or (_41015_, _41014_, _41011_);
  or (_41016_, _41015_, _41010_);
  and (_41017_, _41016_, _40973_);
  not (_41018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_41019_, _40973_, _41018_);
  or (_43232_, _41019_, _41017_);
  nand (_41020_, _40957_, _26598_);
  nor (_41021_, _41020_, _29154_);
  nor (_41022_, _38486_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41023_, _26598_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41024_, _16612_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41025_, _41024_, _41023_);
  or (_41026_, _41025_, _41022_);
  or (_41027_, _41026_, _41021_);
  and (_41028_, _41027_, _40973_);
  not (_41029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_41030_, _40973_, _41029_);
  or (_43238_, _41030_, _41028_);
  nand (_41031_, _40957_, _26664_);
  nor (_41032_, _41031_, _29154_);
  nor (_41033_, _38479_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41034_, _26664_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41035_, _17595_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41036_, _41035_, _41034_);
  or (_41037_, _41036_, _41033_);
  or (_41038_, _41037_, _41032_);
  and (_41039_, _41038_, _40973_);
  not (_41040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_41041_, _40973_, _41040_);
  or (_43244_, _41041_, _41039_);
  nand (_41042_, _40957_, _26565_);
  nor (_41043_, _41042_, _29154_);
  nor (_41044_, _38472_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41045_, _26565_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41046_, _16952_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41047_, _41046_, _41045_);
  or (_41048_, _41047_, _41044_);
  or (_41049_, _41048_, _41043_);
  and (_41050_, _41049_, _40973_);
  not (_41051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_41052_, _40973_, _41051_);
  or (_43250_, _41052_, _41050_);
  not (_41053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_41054_, _40973_, _41053_);
  and (_41055_, _40973_, _40965_);
  or (_43253_, _41055_, _41054_);
  and (_41056_, _40982_, _40812_);
  and (_41057_, _40950_, _40795_);
  and (_41058_, _41057_, _40970_);
  and (_41059_, _41058_, _41056_);
  not (_41060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_41061_, _41058_, _41060_);
  or (_43261_, _41061_, _41059_);
  and (_41062_, _40997_, _40812_);
  and (_41063_, _41058_, _41062_);
  not (_41064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_41065_, _41058_, _41064_);
  or (_43265_, _41065_, _41063_);
  and (_41066_, _41008_, _40812_);
  and (_41067_, _41058_, _41066_);
  not (_41068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_41069_, _41058_, _41068_);
  or (_43269_, _41069_, _41067_);
  and (_41070_, _41016_, _40812_);
  and (_41071_, _41058_, _41070_);
  not (_41072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_41073_, _41058_, _41072_);
  or (_43273_, _41073_, _41071_);
  and (_41074_, _41027_, _40812_);
  and (_41075_, _41058_, _41074_);
  not (_41076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_41077_, _41058_, _41076_);
  or (_43277_, _41077_, _41075_);
  and (_41078_, _41038_, _40812_);
  and (_41079_, _41058_, _41078_);
  not (_41080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_41081_, _41058_, _41080_);
  or (_43279_, _41081_, _41079_);
  and (_41082_, _41049_, _40812_);
  and (_41083_, _41058_, _41082_);
  not (_41084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_41085_, _41058_, _41084_);
  or (_43282_, _41085_, _41083_);
  and (_41086_, _41058_, _40966_);
  nor (_41087_, _41058_, _40837_);
  or (_43285_, _41087_, _41086_);
  and (_41088_, _40951_, _40591_);
  and (_41089_, _41088_, _40970_);
  and (_41090_, _41089_, _41056_);
  not (_41091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_41092_, _41089_, _41091_);
  or (_43293_, _41092_, _41090_);
  and (_41093_, _41089_, _41062_);
  not (_41094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_41095_, _41089_, _41094_);
  or (_43297_, _41095_, _41093_);
  and (_41096_, _41089_, _41066_);
  not (_41097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_41098_, _41089_, _41097_);
  or (_43301_, _41098_, _41096_);
  and (_41099_, _41089_, _41070_);
  not (_41100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_41101_, _41089_, _41100_);
  or (_43305_, _41101_, _41099_);
  and (_41102_, _41089_, _41074_);
  not (_41103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_41104_, _41089_, _41103_);
  or (_43309_, _41104_, _41102_);
  and (_41105_, _41089_, _41078_);
  not (_41106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_41107_, _41089_, _41106_);
  or (_43313_, _41107_, _41105_);
  and (_41108_, _41089_, _41082_);
  not (_41109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_41110_, _41089_, _41109_);
  or (_43317_, _41110_, _41108_);
  and (_41111_, _41089_, _40966_);
  not (_41112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_41113_, _41089_, _41112_);
  or (_43320_, _41113_, _41111_);
  and (_41114_, _40970_, _40952_);
  and (_41115_, _41114_, _41056_);
  not (_41116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_41117_, _41114_, _41116_);
  or (_43326_, _41117_, _41115_);
  and (_41118_, _41114_, _41062_);
  not (_41119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_41120_, _41114_, _41119_);
  or (_43330_, _41120_, _41118_);
  and (_41121_, _41114_, _41066_);
  not (_41122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_41123_, _41114_, _41122_);
  or (_43334_, _41123_, _41121_);
  and (_41124_, _41114_, _41070_);
  not (_41125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_41126_, _41114_, _41125_);
  or (_43338_, _41126_, _41124_);
  and (_41127_, _41114_, _41074_);
  not (_41128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_41129_, _41114_, _41128_);
  or (_43342_, _41129_, _41127_);
  and (_41130_, _41114_, _41078_);
  not (_41131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_41132_, _41114_, _41131_);
  or (_43346_, _41132_, _41130_);
  and (_41133_, _41114_, _41082_);
  not (_41134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_41135_, _41114_, _41134_);
  or (_43350_, _41135_, _41133_);
  and (_41136_, _41114_, _40966_);
  nor (_41137_, _41114_, _40850_);
  or (_43353_, _41137_, _41136_);
  and (_41138_, _40954_, _40638_);
  and (_41139_, _41138_, _40971_);
  and (_41140_, _41139_, _41056_);
  not (_41141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_41142_, _41139_, _41141_);
  or (_43361_, _41142_, _41140_);
  and (_41143_, _41139_, _41062_);
  not (_41144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_41145_, _41139_, _41144_);
  or (_43365_, _41145_, _41143_);
  and (_41146_, _41139_, _41066_);
  not (_41147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_41148_, _41139_, _41147_);
  or (_43369_, _41148_, _41146_);
  and (_41149_, _41139_, _41070_);
  not (_41150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_41151_, _41139_, _41150_);
  or (_43373_, _41151_, _41149_);
  and (_41152_, _41139_, _41074_);
  not (_41153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_41154_, _41139_, _41153_);
  or (_43389_, _41154_, _41152_);
  and (_41155_, _41139_, _41078_);
  not (_41156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_41157_, _41139_, _41156_);
  or (_43409_, _41157_, _41155_);
  and (_41158_, _41139_, _41082_);
  not (_41159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_41160_, _41139_, _41159_);
  or (_43427_, _41160_, _41158_);
  and (_41161_, _41139_, _40966_);
  not (_41162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_41163_, _41139_, _41162_);
  or (_43438_, _41163_, _41161_);
  and (_41164_, _41138_, _41057_);
  and (_41165_, _41164_, _41056_);
  not (_41166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_41167_, _41164_, _41166_);
  or (_43463_, _41167_, _41165_);
  and (_41168_, _41164_, _41062_);
  not (_41169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_41170_, _41164_, _41169_);
  or (_43482_, _41170_, _41168_);
  and (_41171_, _41164_, _41066_);
  not (_41172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_41173_, _41164_, _41172_);
  or (_43502_, _41173_, _41171_);
  and (_41174_, _41164_, _41070_);
  not (_41175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_41176_, _41164_, _41175_);
  or (_43521_, _41176_, _41174_);
  and (_41177_, _41164_, _41074_);
  not (_41178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_41179_, _41164_, _41178_);
  or (_43541_, _41179_, _41177_);
  and (_41180_, _41164_, _41078_);
  not (_41181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_41182_, _41164_, _41181_);
  or (_43561_, _41182_, _41180_);
  and (_41183_, _41164_, _41082_);
  not (_41184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_41185_, _41164_, _41184_);
  or (_43579_, _41185_, _41183_);
  and (_41186_, _41164_, _40966_);
  nor (_41187_, _41164_, _40878_);
  or (_43590_, _41187_, _41186_);
  and (_41188_, _41138_, _41088_);
  and (_41189_, _41188_, _41056_);
  not (_41190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_41191_, _41188_, _41190_);
  or (_43615_, _41191_, _41189_);
  and (_41192_, _41188_, _41062_);
  not (_41193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_41194_, _41188_, _41193_);
  or (_43619_, _41194_, _41192_);
  and (_41195_, _41188_, _41066_);
  not (_41196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_41197_, _41188_, _41196_);
  or (_43623_, _41197_, _41195_);
  and (_41198_, _41188_, _41070_);
  not (_41199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_41200_, _41188_, _41199_);
  or (_43627_, _41200_, _41198_);
  and (_41201_, _41188_, _41074_);
  not (_41202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_41203_, _41188_, _41202_);
  or (_43631_, _41203_, _41201_);
  and (_41204_, _41188_, _41078_);
  not (_41205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_41206_, _41188_, _41205_);
  or (_43635_, _41206_, _41204_);
  and (_41207_, _41188_, _41082_);
  not (_41208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_41209_, _41188_, _41208_);
  or (_43639_, _41209_, _41207_);
  and (_41210_, _41188_, _40966_);
  not (_41211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_41212_, _41188_, _41211_);
  or (_43642_, _41212_, _41210_);
  and (_41213_, _41138_, _40952_);
  and (_41214_, _41213_, _41056_);
  not (_41215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_41216_, _41213_, _41215_);
  or (_43647_, _41216_, _41214_);
  and (_41217_, _41213_, _41062_);
  not (_41218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_41219_, _41213_, _41218_);
  or (_43651_, _41219_, _41217_);
  and (_41220_, _41213_, _41066_);
  not (_41221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_41222_, _41213_, _41221_);
  or (_43655_, _41222_, _41220_);
  and (_41223_, _41213_, _41070_);
  not (_41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_41225_, _41213_, _41224_);
  or (_43659_, _41225_, _41223_);
  and (_41226_, _41213_, _41074_);
  not (_41227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_41228_, _41213_, _41227_);
  or (_43663_, _41228_, _41226_);
  and (_41229_, _41213_, _41078_);
  not (_41230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_41231_, _41213_, _41230_);
  or (_43667_, _41231_, _41229_);
  and (_41232_, _41213_, _41082_);
  not (_41233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_41234_, _41213_, _41233_);
  or (_43671_, _41234_, _41232_);
  and (_41235_, _41213_, _40966_);
  nor (_41236_, _41213_, _40889_);
  or (_43674_, _41236_, _41235_);
  and (_41237_, _40953_, _40512_);
  and (_41238_, _41237_, _40971_);
  and (_41239_, _41238_, _41056_);
  not (_41240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_41241_, _41238_, _41240_);
  or (_43682_, _41241_, _41239_);
  and (_41242_, _41238_, _41062_);
  not (_41243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_41244_, _41238_, _41243_);
  or (_43686_, _41244_, _41242_);
  and (_41245_, _41238_, _41066_);
  not (_41246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_41247_, _41238_, _41246_);
  or (_43689_, _41247_, _41245_);
  and (_41248_, _41238_, _41070_);
  not (_41249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_41250_, _41238_, _41249_);
  or (_43693_, _41250_, _41248_);
  and (_41251_, _41238_, _41074_);
  not (_41252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_41253_, _41238_, _41252_);
  or (_43697_, _41253_, _41251_);
  and (_41254_, _41238_, _41078_);
  not (_41255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_41256_, _41238_, _41255_);
  or (_43701_, _41256_, _41254_);
  and (_41257_, _41238_, _41082_);
  not (_41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_41259_, _41238_, _41258_);
  or (_43705_, _41259_, _41257_);
  and (_41260_, _41238_, _40966_);
  nor (_41261_, _41238_, _40919_);
  or (_43708_, _41261_, _41260_);
  and (_41262_, _41237_, _41057_);
  and (_41263_, _41262_, _41056_);
  not (_41264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_41265_, _41262_, _41264_);
  or (_43713_, _41265_, _41263_);
  and (_41266_, _41262_, _41062_);
  not (_41267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_41268_, _41262_, _41267_);
  or (_43717_, _41268_, _41266_);
  and (_41269_, _41262_, _41066_);
  not (_41270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_41271_, _41262_, _41270_);
  or (_43721_, _41271_, _41269_);
  and (_41272_, _41262_, _41070_);
  not (_41273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_41274_, _41262_, _41273_);
  or (_43725_, _41274_, _41272_);
  and (_41275_, _41262_, _41074_);
  not (_41276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_41277_, _41262_, _41276_);
  or (_43729_, _41277_, _41275_);
  and (_41278_, _41262_, _41078_);
  not (_41279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_41280_, _41262_, _41279_);
  or (_43733_, _41280_, _41278_);
  and (_41281_, _41262_, _41082_);
  not (_41282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_41283_, _41262_, _41282_);
  or (_43737_, _41283_, _41281_);
  and (_41284_, _41262_, _40966_);
  not (_41285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_41286_, _41262_, _41285_);
  or (_43740_, _41286_, _41284_);
  and (_41287_, _41237_, _41088_);
  and (_41288_, _41287_, _41056_);
  not (_41289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_41290_, _41287_, _41289_);
  or (_43745_, _41290_, _41288_);
  and (_41291_, _41287_, _41062_);
  not (_41292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_41293_, _41287_, _41292_);
  or (_43749_, _41293_, _41291_);
  and (_41294_, _41287_, _41066_);
  not (_41295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_41296_, _41287_, _41295_);
  or (_43753_, _41296_, _41294_);
  and (_41297_, _41287_, _41070_);
  not (_41299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_41301_, _41287_, _41299_);
  or (_43757_, _41301_, _41297_);
  and (_41304_, _41287_, _41074_);
  not (_41306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_41308_, _41287_, _41306_);
  or (_43761_, _41308_, _41304_);
  and (_41311_, _41287_, _41078_);
  not (_41313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_41315_, _41287_, _41313_);
  or (_43765_, _41315_, _41311_);
  and (_41318_, _41287_, _41082_);
  not (_41320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_41322_, _41287_, _41320_);
  or (_43769_, _41322_, _41318_);
  and (_41325_, _41287_, _40966_);
  nor (_41327_, _41287_, _40925_);
  or (_43772_, _41327_, _41325_);
  and (_41330_, _41237_, _40952_);
  and (_41332_, _41330_, _41056_);
  not (_41334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_41336_, _41330_, _41334_);
  or (_43777_, _41336_, _41332_);
  and (_41339_, _41330_, _41062_);
  not (_41341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_41343_, _41330_, _41341_);
  or (_43781_, _41343_, _41339_);
  and (_41346_, _41330_, _41066_);
  not (_41347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_41348_, _41330_, _41347_);
  or (_43785_, _41348_, _41346_);
  and (_41349_, _41330_, _41070_);
  not (_41350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_41351_, _41330_, _41350_);
  or (_43789_, _41351_, _41349_);
  and (_41352_, _41330_, _41074_);
  not (_41353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_41354_, _41330_, _41353_);
  or (_43793_, _41354_, _41352_);
  and (_41355_, _41330_, _41078_);
  not (_41356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_41357_, _41330_, _41356_);
  or (_43797_, _41357_, _41355_);
  and (_41358_, _41330_, _41082_);
  not (_41359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_41360_, _41330_, _41359_);
  or (_43801_, _41360_, _41358_);
  and (_41361_, _41330_, _40966_);
  not (_41362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_41363_, _41330_, _41362_);
  or (_43804_, _41363_, _41361_);
  and (_41364_, _40971_, _40955_);
  and (_41365_, _41364_, _41056_);
  not (_41366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_41367_, _41364_, _41366_);
  or (_43810_, _41367_, _41365_);
  and (_41368_, _41364_, _41062_);
  not (_41369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_41370_, _41364_, _41369_);
  or (_43814_, _41370_, _41368_);
  and (_41371_, _41364_, _41066_);
  not (_41372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_41373_, _41364_, _41372_);
  or (_43818_, _41373_, _41371_);
  and (_41374_, _41364_, _41070_);
  not (_41375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_41376_, _41364_, _41375_);
  or (_43822_, _41376_, _41374_);
  and (_41377_, _41364_, _41074_);
  not (_41378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_41379_, _41364_, _41378_);
  or (_43826_, _41379_, _41377_);
  and (_41380_, _41364_, _41078_);
  not (_41381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_41382_, _41364_, _41381_);
  or (_43830_, _41382_, _41380_);
  and (_41383_, _41364_, _41082_);
  not (_41384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_41385_, _41364_, _41384_);
  or (_43834_, _41385_, _41383_);
  and (_41386_, _41364_, _40966_);
  nor (_41387_, _41364_, _40931_);
  or (_43837_, _41387_, _41386_);
  and (_41388_, _41057_, _40955_);
  and (_41389_, _41388_, _41056_);
  not (_41390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_41391_, _41388_, _41390_);
  or (_43842_, _41391_, _41389_);
  and (_41392_, _41388_, _41062_);
  not (_41393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_41394_, _41388_, _41393_);
  or (_43846_, _41394_, _41392_);
  and (_41395_, _41388_, _41066_);
  not (_41396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_41397_, _41388_, _41396_);
  or (_43850_, _41397_, _41395_);
  and (_41398_, _41388_, _41070_);
  not (_41399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_41400_, _41388_, _41399_);
  or (_43854_, _41400_, _41398_);
  and (_41401_, _41388_, _41074_);
  not (_41402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_41403_, _41388_, _41402_);
  or (_43858_, _41403_, _41401_);
  and (_41404_, _41388_, _41078_);
  not (_41405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_41406_, _41388_, _41405_);
  or (_43862_, _41406_, _41404_);
  and (_41407_, _41388_, _41082_);
  not (_41408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_41409_, _41388_, _41408_);
  or (_43866_, _41409_, _41407_);
  and (_41410_, _41388_, _40966_);
  not (_41411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_41412_, _41388_, _41411_);
  or (_43869_, _41412_, _41410_);
  and (_41413_, _41088_, _40955_);
  and (_41414_, _41413_, _41056_);
  not (_41415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_41416_, _41413_, _41415_);
  or (_43874_, _41416_, _41414_);
  and (_41417_, _41413_, _41062_);
  not (_41418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_41419_, _41413_, _41418_);
  or (_43878_, _41419_, _41417_);
  and (_41420_, _41413_, _41066_);
  not (_41421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_41422_, _41413_, _41421_);
  or (_43882_, _41422_, _41420_);
  and (_41423_, _41413_, _41070_);
  not (_41424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_41425_, _41413_, _41424_);
  or (_43886_, _41425_, _41423_);
  and (_41426_, _41413_, _41074_);
  not (_41427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_41428_, _41413_, _41427_);
  or (_43890_, _41428_, _41426_);
  and (_41429_, _41413_, _41078_);
  not (_41430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_41431_, _41413_, _41430_);
  or (_43894_, _41431_, _41429_);
  and (_41432_, _41413_, _41082_);
  not (_41433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_41434_, _41413_, _41433_);
  or (_43898_, _41434_, _41432_);
  and (_41435_, _41413_, _40966_);
  nor (_41436_, _41413_, _40937_);
  or (_43901_, _41436_, _41435_);
  and (_41437_, _41056_, _40956_);
  not (_41438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_41439_, _40956_, _41438_);
  or (_43906_, _41439_, _41437_);
  and (_41440_, _41062_, _40956_);
  not (_41441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_41442_, _40956_, _41441_);
  or (_43910_, _41442_, _41440_);
  and (_41443_, _41066_, _40956_);
  not (_41444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_41445_, _40956_, _41444_);
  or (_43914_, _41445_, _41443_);
  and (_41446_, _41070_, _40956_);
  not (_41447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_41448_, _40956_, _41447_);
  or (_43918_, _41448_, _41446_);
  and (_41449_, _41074_, _40956_);
  not (_41450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_41451_, _40956_, _41450_);
  or (_43922_, _41451_, _41449_);
  and (_41452_, _41078_, _40956_);
  not (_41453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_41454_, _40956_, _41453_);
  or (_43926_, _41454_, _41452_);
  and (_41455_, _41082_, _40956_);
  not (_41456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_41457_, _40956_, _41456_);
  or (_43930_, _41457_, _41455_);
  and (_41458_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_41459_, _40588_, _41060_);
  or (_41460_, _41459_, _41458_);
  and (_41461_, _41460_, _40787_);
  nor (_41462_, _40588_, _41116_);
  and (_41463_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_41464_, _41463_, _41462_);
  and (_41465_, _41464_, _40849_);
  or (_41466_, _41465_, _41461_);
  or (_41467_, _41466_, _40833_);
  and (_41468_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_41469_, _40588_, _41166_);
  or (_41470_, _41469_, _41468_);
  and (_41471_, _41470_, _40787_);
  nor (_41472_, _40588_, _41215_);
  and (_41473_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_41474_, _41473_, _41472_);
  and (_41475_, _41474_, _40849_);
  or (_41476_, _41475_, _41471_);
  or (_41477_, _41476_, _40508_);
  and (_41478_, _41477_, _40873_);
  and (_41479_, _41478_, _41467_);
  nand (_41480_, _40588_, _41240_);
  or (_41481_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_41482_, _41481_, _41480_);
  and (_41483_, _41482_, _40787_);
  or (_41484_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand (_41485_, _40588_, _41289_);
  and (_41486_, _41485_, _41484_);
  and (_41487_, _41486_, _40849_);
  or (_41488_, _41487_, _41483_);
  or (_41489_, _41488_, _40833_);
  nand (_41490_, _40588_, _41366_);
  or (_41491_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_41492_, _41491_, _41490_);
  and (_41493_, _41492_, _40787_);
  or (_41494_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand (_41495_, _40588_, _41415_);
  and (_41496_, _41495_, _41494_);
  and (_41497_, _41496_, _40849_);
  or (_41498_, _41497_, _41493_);
  or (_41499_, _41498_, _40508_);
  and (_41500_, _41499_, _40634_);
  and (_41501_, _41500_, _41489_);
  or (_41502_, _41501_, _41479_);
  or (_41503_, _41502_, _40827_);
  or (_41504_, _40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_41505_, _41504_, _41894_);
  and (_01362_, _41505_, _41503_);
  and (_41506_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_41507_, _40588_, _41064_);
  or (_41508_, _41507_, _41506_);
  and (_41509_, _41508_, _40787_);
  nor (_41510_, _40588_, _41119_);
  and (_41511_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_41512_, _41511_, _41510_);
  and (_41513_, _41512_, _40849_);
  or (_41514_, _41513_, _41509_);
  or (_41515_, _41514_, _40833_);
  and (_41516_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_41517_, _40588_, _41169_);
  or (_41518_, _41517_, _41516_);
  and (_41519_, _41518_, _40787_);
  nor (_41520_, _40588_, _41218_);
  and (_41521_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_41522_, _41521_, _41520_);
  and (_41523_, _41522_, _40849_);
  or (_41524_, _41523_, _41519_);
  or (_41525_, _41524_, _40508_);
  and (_41526_, _41525_, _40873_);
  and (_41527_, _41526_, _41515_);
  nand (_41528_, _40588_, _41243_);
  or (_41529_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_41530_, _41529_, _41528_);
  and (_41531_, _41530_, _40787_);
  or (_41532_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand (_41533_, _40588_, _41292_);
  and (_41534_, _41533_, _41532_);
  and (_41535_, _41534_, _40849_);
  or (_41536_, _41535_, _41531_);
  or (_41537_, _41536_, _40833_);
  nand (_41538_, _40588_, _41369_);
  or (_41539_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_41540_, _41539_, _41538_);
  and (_41541_, _41540_, _40787_);
  or (_41542_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand (_41543_, _40588_, _41418_);
  and (_41544_, _41543_, _41542_);
  and (_41545_, _41544_, _40849_);
  or (_41546_, _41545_, _41541_);
  or (_41547_, _41546_, _40508_);
  and (_41548_, _41547_, _40634_);
  and (_41549_, _41548_, _41537_);
  or (_41550_, _41549_, _41527_);
  or (_41551_, _41550_, _40827_);
  or (_41552_, _40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_41553_, _41552_, _41894_);
  and (_01364_, _41553_, _41551_);
  and (_41554_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_41555_, _40588_, _41068_);
  or (_41556_, _41555_, _41554_);
  and (_41557_, _41556_, _40787_);
  nor (_41558_, _40588_, _41122_);
  and (_41559_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_41560_, _41559_, _41558_);
  and (_41561_, _41560_, _40849_);
  or (_41562_, _41561_, _41557_);
  or (_41563_, _41562_, _40833_);
  and (_41564_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_41565_, _40588_, _41172_);
  or (_41566_, _41565_, _41564_);
  and (_41567_, _41566_, _40787_);
  nor (_41568_, _40588_, _41221_);
  and (_41569_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_41570_, _41569_, _41568_);
  and (_41571_, _41570_, _40849_);
  or (_41572_, _41571_, _41567_);
  or (_41573_, _41572_, _40508_);
  and (_41574_, _41573_, _40873_);
  and (_41575_, _41574_, _41563_);
  nand (_41576_, _40588_, _41246_);
  or (_41577_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_41578_, _41577_, _41576_);
  and (_41579_, _41578_, _40787_);
  or (_41580_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_41581_, _40588_, _41295_);
  and (_41582_, _41581_, _41580_);
  and (_41583_, _41582_, _40849_);
  or (_41584_, _41583_, _41579_);
  or (_41585_, _41584_, _40833_);
  nand (_41586_, _40588_, _41372_);
  or (_41587_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_41588_, _41587_, _41586_);
  and (_41589_, _41588_, _40787_);
  or (_41590_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_41591_, _40588_, _41421_);
  and (_41592_, _41591_, _41590_);
  and (_41593_, _41592_, _40849_);
  or (_41594_, _41593_, _41589_);
  or (_41595_, _41594_, _40508_);
  and (_41596_, _41595_, _40634_);
  and (_41597_, _41596_, _41585_);
  or (_41598_, _41597_, _41575_);
  or (_41599_, _41598_, _40827_);
  or (_41600_, _40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_41601_, _41600_, _41894_);
  and (_01366_, _41601_, _41599_);
  and (_41602_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_41603_, _40588_, _41072_);
  or (_41604_, _41603_, _41602_);
  and (_41605_, _41604_, _40787_);
  nor (_41606_, _40588_, _41125_);
  and (_41607_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_41608_, _41607_, _41606_);
  and (_41609_, _41608_, _40849_);
  or (_41610_, _41609_, _41605_);
  or (_41611_, _41610_, _40833_);
  and (_41612_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_41613_, _40588_, _41175_);
  or (_41614_, _41613_, _41612_);
  and (_41615_, _41614_, _40787_);
  nor (_41616_, _40588_, _41224_);
  and (_41617_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_41618_, _41617_, _41616_);
  and (_41619_, _41618_, _40849_);
  or (_41620_, _41619_, _41615_);
  or (_41621_, _41620_, _40508_);
  and (_41622_, _41621_, _40873_);
  and (_41623_, _41622_, _41611_);
  nand (_41624_, _40588_, _41249_);
  or (_41625_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_41626_, _41625_, _41624_);
  and (_41627_, _41626_, _40787_);
  or (_41628_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_41629_, _40588_, _41299_);
  and (_41630_, _41629_, _41628_);
  and (_41631_, _41630_, _40849_);
  or (_41632_, _41631_, _41627_);
  or (_41633_, _41632_, _40833_);
  nand (_41634_, _40588_, _41375_);
  or (_41635_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_41636_, _41635_, _41634_);
  and (_41637_, _41636_, _40787_);
  or (_41638_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_41639_, _40588_, _41424_);
  and (_41640_, _41639_, _41638_);
  and (_41641_, _41640_, _40849_);
  or (_41642_, _41641_, _41637_);
  or (_41643_, _41642_, _40508_);
  and (_41644_, _41643_, _40634_);
  and (_41645_, _41644_, _41633_);
  or (_41646_, _41645_, _41623_);
  or (_41647_, _41646_, _40827_);
  or (_41648_, _40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_41649_, _41648_, _41894_);
  and (_01368_, _41649_, _41647_);
  and (_41650_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_41651_, _40588_, _41076_);
  or (_41652_, _41651_, _41650_);
  and (_41653_, _41652_, _40787_);
  nor (_41654_, _40588_, _41128_);
  and (_41655_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_41656_, _41655_, _41654_);
  and (_41657_, _41656_, _40849_);
  or (_41658_, _41657_, _41653_);
  or (_41659_, _41658_, _40833_);
  and (_41660_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_41661_, _40588_, _41178_);
  or (_41662_, _41661_, _41660_);
  and (_41663_, _41662_, _40787_);
  nor (_41664_, _40588_, _41227_);
  and (_41665_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_41666_, _41665_, _41664_);
  and (_41667_, _41666_, _40849_);
  or (_41668_, _41667_, _41663_);
  or (_41669_, _41668_, _40508_);
  and (_41670_, _41669_, _40873_);
  and (_41671_, _41670_, _41659_);
  nand (_41672_, _40588_, _41252_);
  or (_41673_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_41674_, _41673_, _41672_);
  and (_41675_, _41674_, _40787_);
  or (_41676_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_41677_, _40588_, _41306_);
  and (_41678_, _41677_, _41676_);
  and (_41679_, _41678_, _40849_);
  or (_41680_, _41679_, _41675_);
  or (_41681_, _41680_, _40833_);
  nand (_41682_, _40588_, _41378_);
  or (_41683_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_41684_, _41683_, _41682_);
  and (_41685_, _41684_, _40787_);
  or (_41686_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_41687_, _40588_, _41427_);
  and (_41688_, _41687_, _41686_);
  and (_41689_, _41688_, _40849_);
  or (_41690_, _41689_, _41685_);
  or (_41691_, _41690_, _40508_);
  and (_41692_, _41691_, _40634_);
  and (_41693_, _41692_, _41681_);
  or (_41694_, _41693_, _41671_);
  or (_41695_, _41694_, _40827_);
  or (_41696_, _40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_41697_, _41696_, _41894_);
  and (_01370_, _41697_, _41695_);
  and (_41698_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_41699_, _40588_, _41080_);
  or (_41700_, _41699_, _41698_);
  and (_41701_, _41700_, _40787_);
  nor (_41702_, _40588_, _41131_);
  and (_41703_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_41704_, _41703_, _41702_);
  and (_41705_, _41704_, _40849_);
  or (_41706_, _41705_, _41701_);
  or (_41707_, _41706_, _40833_);
  and (_41708_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_41709_, _40588_, _41181_);
  or (_41710_, _41709_, _41708_);
  and (_41711_, _41710_, _40787_);
  nor (_41712_, _40588_, _41230_);
  and (_41713_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_41714_, _41713_, _41712_);
  and (_41715_, _41714_, _40849_);
  or (_41716_, _41715_, _41711_);
  or (_41717_, _41716_, _40508_);
  and (_41718_, _41717_, _40873_);
  and (_41719_, _41718_, _41707_);
  nand (_41720_, _40588_, _41255_);
  or (_41721_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_41722_, _41721_, _41720_);
  and (_41723_, _41722_, _40787_);
  or (_41724_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_41725_, _40588_, _41313_);
  and (_41726_, _41725_, _41724_);
  and (_41727_, _41726_, _40849_);
  or (_41728_, _41727_, _41723_);
  or (_41729_, _41728_, _40833_);
  nand (_41730_, _40588_, _41381_);
  or (_41731_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_41732_, _41731_, _41730_);
  and (_41733_, _41732_, _40787_);
  or (_41734_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_41735_, _40588_, _41430_);
  and (_41736_, _41735_, _41734_);
  and (_41737_, _41736_, _40849_);
  or (_41738_, _41737_, _41733_);
  or (_41739_, _41738_, _40508_);
  and (_41740_, _41739_, _40634_);
  and (_41741_, _41740_, _41729_);
  or (_41742_, _41741_, _41719_);
  or (_41743_, _41742_, _40827_);
  or (_41744_, _40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_41745_, _41744_, _41894_);
  and (_01372_, _41745_, _41743_);
  and (_41746_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_41747_, _40588_, _41084_);
  or (_41748_, _41747_, _41746_);
  and (_41749_, _41748_, _40787_);
  nor (_41750_, _40588_, _41134_);
  and (_41751_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_41752_, _41751_, _41750_);
  and (_41753_, _41752_, _40849_);
  or (_41754_, _41753_, _41749_);
  or (_41755_, _41754_, _40833_);
  and (_41756_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_41757_, _40588_, _41184_);
  or (_41758_, _41757_, _41756_);
  and (_41759_, _41758_, _40787_);
  nor (_41760_, _40588_, _41233_);
  and (_41761_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_41762_, _41761_, _41760_);
  and (_41763_, _41762_, _40849_);
  or (_41764_, _41763_, _41759_);
  or (_41765_, _41764_, _40508_);
  and (_41766_, _41765_, _40873_);
  and (_41767_, _41766_, _41755_);
  nand (_41768_, _40588_, _41258_);
  or (_41769_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_41770_, _41769_, _41768_);
  and (_41771_, _41770_, _40787_);
  or (_41772_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_41773_, _40588_, _41320_);
  and (_41774_, _41773_, _41772_);
  and (_41775_, _41774_, _40849_);
  or (_41776_, _41775_, _41771_);
  or (_41777_, _41776_, _40833_);
  nand (_41778_, _40588_, _41384_);
  or (_41779_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_41780_, _41779_, _41778_);
  and (_41781_, _41780_, _40787_);
  or (_41782_, _40588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_41783_, _40588_, _41433_);
  and (_41784_, _41783_, _41782_);
  and (_41785_, _41784_, _40849_);
  or (_41786_, _41785_, _41781_);
  or (_41787_, _41786_, _40508_);
  and (_41788_, _41787_, _40634_);
  and (_41789_, _41788_, _41777_);
  or (_41790_, _41789_, _41767_);
  or (_41791_, _41790_, _40827_);
  or (_41792_, _40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_41793_, _41792_, _41894_);
  and (_01374_, _41793_, _41791_);
  or (_41794_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_41795_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_41796_, _41795_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_41797_, _41796_, _41794_);
  nand (_41798_, _41797_, _41894_);
  or (_41799_, \oc8051_gm_cxrom_1.cell0.data [7], _41894_);
  and (_01382_, _41799_, _41798_);
  or (_41800_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41801_, \oc8051_gm_cxrom_1.cell0.data [0], _41795_);
  nand (_41802_, _41801_, _41800_);
  nand (_41803_, _41802_, _41894_);
  or (_41804_, \oc8051_gm_cxrom_1.cell0.data [0], _41894_);
  and (_01389_, _41804_, _41803_);
  or (_41805_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41806_, \oc8051_gm_cxrom_1.cell0.data [1], _41795_);
  nand (_41807_, _41806_, _41805_);
  nand (_41808_, _41807_, _41894_);
  or (_41809_, \oc8051_gm_cxrom_1.cell0.data [1], _41894_);
  and (_01393_, _41809_, _41808_);
  or (_41810_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41811_, \oc8051_gm_cxrom_1.cell0.data [2], _41795_);
  nand (_41812_, _41811_, _41810_);
  nand (_41813_, _41812_, _41894_);
  or (_41814_, \oc8051_gm_cxrom_1.cell0.data [2], _41894_);
  and (_01397_, _41814_, _41813_);
  or (_41815_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41816_, \oc8051_gm_cxrom_1.cell0.data [3], _41795_);
  nand (_41817_, _41816_, _41815_);
  nand (_41818_, _41817_, _41894_);
  or (_41819_, \oc8051_gm_cxrom_1.cell0.data [3], _41894_);
  and (_01401_, _41819_, _41818_);
  or (_41820_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41821_, \oc8051_gm_cxrom_1.cell0.data [4], _41795_);
  nand (_41822_, _41821_, _41820_);
  nand (_41823_, _41822_, _41894_);
  or (_41824_, \oc8051_gm_cxrom_1.cell0.data [4], _41894_);
  and (_01405_, _41824_, _41823_);
  or (_41825_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41826_, \oc8051_gm_cxrom_1.cell0.data [5], _41795_);
  nand (_41827_, _41826_, _41825_);
  nand (_41828_, _41827_, _41894_);
  or (_41829_, \oc8051_gm_cxrom_1.cell0.data [5], _41894_);
  and (_01409_, _41829_, _41828_);
  or (_41830_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41831_, \oc8051_gm_cxrom_1.cell0.data [6], _41795_);
  nand (_41832_, _41831_, _41830_);
  nand (_41833_, _41832_, _41894_);
  or (_41834_, \oc8051_gm_cxrom_1.cell0.data [6], _41894_);
  and (_01413_, _41834_, _41833_);
  or (_41835_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_41837_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_41838_, _41837_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_41840_, _41838_, _41835_);
  nand (_41842_, _41840_, _41894_);
  or (_41843_, \oc8051_gm_cxrom_1.cell1.data [7], _41894_);
  and (_01435_, _41843_, _41842_);
  or (_41846_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41848_, \oc8051_gm_cxrom_1.cell1.data [0], _41837_);
  nand (_41850_, _41848_, _41846_);
  nand (_41851_, _41850_, _41894_);
  or (_41852_, \oc8051_gm_cxrom_1.cell1.data [0], _41894_);
  and (_01442_, _41852_, _41851_);
  or (_41853_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41854_, \oc8051_gm_cxrom_1.cell1.data [1], _41837_);
  nand (_41855_, _41854_, _41853_);
  nand (_41856_, _41855_, _41894_);
  or (_41857_, \oc8051_gm_cxrom_1.cell1.data [1], _41894_);
  and (_01446_, _41857_, _41856_);
  or (_41858_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41859_, \oc8051_gm_cxrom_1.cell1.data [2], _41837_);
  nand (_41860_, _41859_, _41858_);
  nand (_41861_, _41860_, _41894_);
  or (_41862_, \oc8051_gm_cxrom_1.cell1.data [2], _41894_);
  and (_01450_, _41862_, _41861_);
  or (_41863_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41864_, \oc8051_gm_cxrom_1.cell1.data [3], _41837_);
  nand (_41865_, _41864_, _41863_);
  nand (_41866_, _41865_, _41894_);
  or (_41867_, \oc8051_gm_cxrom_1.cell1.data [3], _41894_);
  and (_01454_, _41867_, _41866_);
  or (_41868_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41869_, \oc8051_gm_cxrom_1.cell1.data [4], _41837_);
  nand (_41870_, _41869_, _41868_);
  nand (_41871_, _41870_, _41894_);
  or (_41872_, \oc8051_gm_cxrom_1.cell1.data [4], _41894_);
  and (_01458_, _41872_, _41871_);
  or (_41873_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41874_, \oc8051_gm_cxrom_1.cell1.data [5], _41837_);
  nand (_41875_, _41874_, _41873_);
  nand (_41876_, _41875_, _41894_);
  or (_41877_, \oc8051_gm_cxrom_1.cell1.data [5], _41894_);
  and (_01462_, _41877_, _41876_);
  or (_41878_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41879_, \oc8051_gm_cxrom_1.cell1.data [6], _41837_);
  nand (_41880_, _41879_, _41878_);
  nand (_41882_, _41880_, _41894_);
  or (_41884_, \oc8051_gm_cxrom_1.cell1.data [6], _41894_);
  and (_01466_, _41884_, _41882_);
  or (_41887_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_41889_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_41891_, _41889_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_41893_, _41891_, _41887_);
  nand (_41895_, _41893_, _41894_);
  or (_41896_, \oc8051_gm_cxrom_1.cell2.data [7], _41894_);
  and (_01488_, _41896_, _41895_);
  or (_41897_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41898_, \oc8051_gm_cxrom_1.cell2.data [0], _41889_);
  nand (_41899_, _41898_, _41897_);
  nand (_41900_, _41899_, _41894_);
  or (_41901_, \oc8051_gm_cxrom_1.cell2.data [0], _41894_);
  and (_01495_, _41901_, _41900_);
  or (_41902_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41903_, \oc8051_gm_cxrom_1.cell2.data [1], _41889_);
  nand (_41904_, _41903_, _41902_);
  nand (_41905_, _41904_, _41894_);
  or (_41906_, \oc8051_gm_cxrom_1.cell2.data [1], _41894_);
  and (_01499_, _41906_, _41905_);
  or (_41907_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41908_, \oc8051_gm_cxrom_1.cell2.data [2], _41889_);
  nand (_41909_, _41908_, _41907_);
  nand (_41910_, _41909_, _41894_);
  or (_41911_, \oc8051_gm_cxrom_1.cell2.data [2], _41894_);
  and (_01503_, _41911_, _41910_);
  or (_41912_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41913_, \oc8051_gm_cxrom_1.cell2.data [3], _41889_);
  nand (_41914_, _41913_, _41912_);
  nand (_41915_, _41914_, _41894_);
  or (_41916_, \oc8051_gm_cxrom_1.cell2.data [3], _41894_);
  and (_01507_, _41916_, _41915_);
  or (_41917_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41918_, \oc8051_gm_cxrom_1.cell2.data [4], _41889_);
  nand (_41919_, _41918_, _41917_);
  nand (_41920_, _41919_, _41894_);
  or (_41921_, \oc8051_gm_cxrom_1.cell2.data [4], _41894_);
  and (_01511_, _41921_, _41920_);
  or (_41922_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41923_, \oc8051_gm_cxrom_1.cell2.data [5], _41889_);
  nand (_41924_, _41923_, _41922_);
  nand (_41925_, _41924_, _41894_);
  or (_41926_, \oc8051_gm_cxrom_1.cell2.data [5], _41894_);
  and (_01515_, _41926_, _41925_);
  or (_41927_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41928_, \oc8051_gm_cxrom_1.cell2.data [6], _41889_);
  nand (_41929_, _41928_, _41927_);
  nand (_41930_, _41929_, _41894_);
  or (_41931_, \oc8051_gm_cxrom_1.cell2.data [6], _41894_);
  and (_01519_, _41931_, _41930_);
  or (_41932_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_41933_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_41934_, _41933_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_41935_, _41934_, _41932_);
  nand (_41936_, _41935_, _41894_);
  or (_41937_, \oc8051_gm_cxrom_1.cell3.data [7], _41894_);
  and (_01540_, _41937_, _41936_);
  or (_41938_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41939_, \oc8051_gm_cxrom_1.cell3.data [0], _41933_);
  nand (_41940_, _41939_, _41938_);
  nand (_41941_, _41940_, _41894_);
  or (_41942_, \oc8051_gm_cxrom_1.cell3.data [0], _41894_);
  and (_01547_, _41942_, _41941_);
  or (_41943_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41944_, \oc8051_gm_cxrom_1.cell3.data [1], _41933_);
  nand (_41945_, _41944_, _41943_);
  nand (_41946_, _41945_, _41894_);
  or (_41947_, \oc8051_gm_cxrom_1.cell3.data [1], _41894_);
  and (_01551_, _41947_, _41946_);
  or (_41948_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41949_, \oc8051_gm_cxrom_1.cell3.data [2], _41933_);
  nand (_41950_, _41949_, _41948_);
  nand (_41951_, _41950_, _41894_);
  or (_41952_, \oc8051_gm_cxrom_1.cell3.data [2], _41894_);
  and (_01555_, _41952_, _41951_);
  or (_41953_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41954_, \oc8051_gm_cxrom_1.cell3.data [3], _41933_);
  nand (_41955_, _41954_, _41953_);
  nand (_41956_, _41955_, _41894_);
  or (_41957_, \oc8051_gm_cxrom_1.cell3.data [3], _41894_);
  and (_01559_, _41957_, _41956_);
  or (_41958_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41959_, \oc8051_gm_cxrom_1.cell3.data [4], _41933_);
  nand (_41960_, _41959_, _41958_);
  nand (_41961_, _41960_, _41894_);
  or (_41962_, \oc8051_gm_cxrom_1.cell3.data [4], _41894_);
  and (_01562_, _41962_, _41961_);
  or (_41963_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41964_, \oc8051_gm_cxrom_1.cell3.data [5], _41933_);
  nand (_41965_, _41964_, _41963_);
  nand (_41966_, _41965_, _41894_);
  or (_41967_, \oc8051_gm_cxrom_1.cell3.data [5], _41894_);
  and (_01566_, _41967_, _41966_);
  or (_41968_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41969_, \oc8051_gm_cxrom_1.cell3.data [6], _41933_);
  nand (_41970_, _41969_, _41968_);
  nand (_41971_, _41970_, _41894_);
  or (_41972_, \oc8051_gm_cxrom_1.cell3.data [6], _41894_);
  and (_01570_, _41972_, _41971_);
  or (_41973_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_41974_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_41975_, _41974_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_41976_, _41975_, _41973_);
  nand (_41977_, _41976_, _41894_);
  or (_41978_, \oc8051_gm_cxrom_1.cell4.data [7], _41894_);
  and (_01592_, _41978_, _41977_);
  or (_41979_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41980_, \oc8051_gm_cxrom_1.cell4.data [0], _41974_);
  nand (_41981_, _41980_, _41979_);
  nand (_41982_, _41981_, _41894_);
  or (_41983_, \oc8051_gm_cxrom_1.cell4.data [0], _41894_);
  and (_01599_, _41983_, _41982_);
  or (_41984_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41985_, \oc8051_gm_cxrom_1.cell4.data [1], _41974_);
  nand (_41986_, _41985_, _41984_);
  nand (_41987_, _41986_, _41894_);
  or (_41988_, \oc8051_gm_cxrom_1.cell4.data [1], _41894_);
  and (_01603_, _41988_, _41987_);
  or (_41989_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41990_, \oc8051_gm_cxrom_1.cell4.data [2], _41974_);
  nand (_41991_, _41990_, _41989_);
  nand (_41992_, _41991_, _41894_);
  or (_41993_, \oc8051_gm_cxrom_1.cell4.data [2], _41894_);
  and (_01607_, _41993_, _41992_);
  or (_41994_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41995_, \oc8051_gm_cxrom_1.cell4.data [3], _41974_);
  nand (_41996_, _41995_, _41994_);
  nand (_41997_, _41996_, _41894_);
  or (_41998_, \oc8051_gm_cxrom_1.cell4.data [3], _41894_);
  and (_01611_, _41998_, _41997_);
  or (_41999_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42000_, \oc8051_gm_cxrom_1.cell4.data [4], _41974_);
  nand (_42001_, _42000_, _41999_);
  nand (_42002_, _42001_, _41894_);
  or (_42003_, \oc8051_gm_cxrom_1.cell4.data [4], _41894_);
  and (_01615_, _42003_, _42002_);
  or (_42004_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42005_, \oc8051_gm_cxrom_1.cell4.data [5], _41974_);
  nand (_42006_, _42005_, _42004_);
  nand (_42007_, _42006_, _41894_);
  or (_42008_, \oc8051_gm_cxrom_1.cell4.data [5], _41894_);
  and (_01619_, _42008_, _42007_);
  or (_42009_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42010_, \oc8051_gm_cxrom_1.cell4.data [6], _41974_);
  nand (_42011_, _42010_, _42009_);
  nand (_42012_, _42011_, _41894_);
  or (_42013_, \oc8051_gm_cxrom_1.cell4.data [6], _41894_);
  and (_01622_, _42013_, _42012_);
  or (_42014_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_42015_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_42016_, _42015_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_42017_, _42016_, _42014_);
  nand (_42018_, _42017_, _41894_);
  or (_42019_, \oc8051_gm_cxrom_1.cell5.data [7], _41894_);
  and (_01644_, _42019_, _42018_);
  or (_42020_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42021_, \oc8051_gm_cxrom_1.cell5.data [0], _42015_);
  nand (_42022_, _42021_, _42020_);
  nand (_42023_, _42022_, _41894_);
  or (_42024_, \oc8051_gm_cxrom_1.cell5.data [0], _41894_);
  and (_01651_, _42024_, _42023_);
  or (_42025_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42026_, \oc8051_gm_cxrom_1.cell5.data [1], _42015_);
  nand (_42027_, _42026_, _42025_);
  nand (_42028_, _42027_, _41894_);
  or (_42029_, \oc8051_gm_cxrom_1.cell5.data [1], _41894_);
  and (_01655_, _42029_, _42028_);
  or (_42030_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42031_, \oc8051_gm_cxrom_1.cell5.data [2], _42015_);
  nand (_42032_, _42031_, _42030_);
  nand (_42033_, _42032_, _41894_);
  or (_42034_, \oc8051_gm_cxrom_1.cell5.data [2], _41894_);
  and (_01659_, _42034_, _42033_);
  or (_42035_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42036_, \oc8051_gm_cxrom_1.cell5.data [3], _42015_);
  nand (_42037_, _42036_, _42035_);
  nand (_42038_, _42037_, _41894_);
  or (_42039_, \oc8051_gm_cxrom_1.cell5.data [3], _41894_);
  and (_01662_, _42039_, _42038_);
  or (_42040_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42041_, \oc8051_gm_cxrom_1.cell5.data [4], _42015_);
  nand (_42042_, _42041_, _42040_);
  nand (_42043_, _42042_, _41894_);
  or (_42044_, \oc8051_gm_cxrom_1.cell5.data [4], _41894_);
  and (_01666_, _42044_, _42043_);
  or (_42045_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42046_, \oc8051_gm_cxrom_1.cell5.data [5], _42015_);
  nand (_42047_, _42046_, _42045_);
  nand (_42048_, _42047_, _41894_);
  or (_42049_, \oc8051_gm_cxrom_1.cell5.data [5], _41894_);
  and (_01670_, _42049_, _42048_);
  or (_42050_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42051_, \oc8051_gm_cxrom_1.cell5.data [6], _42015_);
  nand (_42052_, _42051_, _42050_);
  nand (_42053_, _42052_, _41894_);
  or (_42054_, \oc8051_gm_cxrom_1.cell5.data [6], _41894_);
  and (_01674_, _42054_, _42053_);
  or (_42055_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_42056_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_42057_, _42056_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_42058_, _42057_, _42055_);
  nand (_42059_, _42058_, _41894_);
  or (_42060_, \oc8051_gm_cxrom_1.cell6.data [7], _41894_);
  and (_01696_, _42060_, _42059_);
  or (_42061_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42062_, \oc8051_gm_cxrom_1.cell6.data [0], _42056_);
  nand (_42063_, _42062_, _42061_);
  nand (_42064_, _42063_, _41894_);
  or (_42065_, \oc8051_gm_cxrom_1.cell6.data [0], _41894_);
  and (_01702_, _42065_, _42064_);
  or (_42066_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42067_, \oc8051_gm_cxrom_1.cell6.data [1], _42056_);
  nand (_42068_, _42067_, _42066_);
  nand (_42069_, _42068_, _41894_);
  or (_42070_, \oc8051_gm_cxrom_1.cell6.data [1], _41894_);
  and (_01706_, _42070_, _42069_);
  or (_42071_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42072_, \oc8051_gm_cxrom_1.cell6.data [2], _42056_);
  nand (_42073_, _42072_, _42071_);
  nand (_42074_, _42073_, _41894_);
  or (_42075_, \oc8051_gm_cxrom_1.cell6.data [2], _41894_);
  and (_01710_, _42075_, _42074_);
  or (_42076_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42077_, \oc8051_gm_cxrom_1.cell6.data [3], _42056_);
  nand (_42078_, _42077_, _42076_);
  nand (_42079_, _42078_, _41894_);
  or (_42080_, \oc8051_gm_cxrom_1.cell6.data [3], _41894_);
  and (_01714_, _42080_, _42079_);
  or (_42081_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42082_, \oc8051_gm_cxrom_1.cell6.data [4], _42056_);
  nand (_42083_, _42082_, _42081_);
  nand (_42084_, _42083_, _41894_);
  or (_42085_, \oc8051_gm_cxrom_1.cell6.data [4], _41894_);
  and (_01718_, _42085_, _42084_);
  or (_42086_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42087_, \oc8051_gm_cxrom_1.cell6.data [5], _42056_);
  nand (_42088_, _42087_, _42086_);
  nand (_42089_, _42088_, _41894_);
  or (_42090_, \oc8051_gm_cxrom_1.cell6.data [5], _41894_);
  and (_01722_, _42090_, _42089_);
  or (_42091_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42092_, \oc8051_gm_cxrom_1.cell6.data [6], _42056_);
  nand (_42093_, _42092_, _42091_);
  nand (_42094_, _42093_, _41894_);
  or (_42095_, \oc8051_gm_cxrom_1.cell6.data [6], _41894_);
  and (_01726_, _42095_, _42094_);
  or (_42096_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_42097_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_42098_, _42097_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_42099_, _42098_, _42096_);
  nand (_42100_, _42099_, _41894_);
  or (_42101_, \oc8051_gm_cxrom_1.cell7.data [7], _41894_);
  and (_01747_, _42101_, _42100_);
  or (_42102_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42103_, \oc8051_gm_cxrom_1.cell7.data [0], _42097_);
  nand (_42104_, _42103_, _42102_);
  nand (_42105_, _42104_, _41894_);
  or (_42106_, \oc8051_gm_cxrom_1.cell7.data [0], _41894_);
  and (_01754_, _42106_, _42105_);
  or (_42107_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42108_, \oc8051_gm_cxrom_1.cell7.data [1], _42097_);
  nand (_42109_, _42108_, _42107_);
  nand (_42110_, _42109_, _41894_);
  or (_42111_, \oc8051_gm_cxrom_1.cell7.data [1], _41894_);
  and (_01758_, _42111_, _42110_);
  or (_42112_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42113_, \oc8051_gm_cxrom_1.cell7.data [2], _42097_);
  nand (_42114_, _42113_, _42112_);
  nand (_42115_, _42114_, _41894_);
  or (_42116_, \oc8051_gm_cxrom_1.cell7.data [2], _41894_);
  and (_01762_, _42116_, _42115_);
  or (_42117_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42118_, \oc8051_gm_cxrom_1.cell7.data [3], _42097_);
  nand (_42119_, _42118_, _42117_);
  nand (_42120_, _42119_, _41894_);
  or (_42121_, \oc8051_gm_cxrom_1.cell7.data [3], _41894_);
  and (_01766_, _42121_, _42120_);
  or (_42122_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42123_, \oc8051_gm_cxrom_1.cell7.data [4], _42097_);
  nand (_42124_, _42123_, _42122_);
  nand (_42125_, _42124_, _41894_);
  or (_42126_, \oc8051_gm_cxrom_1.cell7.data [4], _41894_);
  and (_01770_, _42126_, _42125_);
  or (_42127_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42128_, \oc8051_gm_cxrom_1.cell7.data [5], _42097_);
  nand (_42129_, _42128_, _42127_);
  nand (_42130_, _42129_, _41894_);
  or (_42131_, \oc8051_gm_cxrom_1.cell7.data [5], _41894_);
  and (_01774_, _42131_, _42130_);
  or (_42132_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42133_, \oc8051_gm_cxrom_1.cell7.data [6], _42097_);
  nand (_42134_, _42133_, _42132_);
  nand (_42135_, _42134_, _41894_);
  or (_42136_, \oc8051_gm_cxrom_1.cell7.data [6], _41894_);
  and (_01777_, _42136_, _42135_);
  or (_42137_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_42138_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_42139_, _42138_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_42140_, _42139_, _42137_);
  nand (_42141_, _42140_, _41894_);
  or (_42142_, \oc8051_gm_cxrom_1.cell8.data [7], _41894_);
  and (_01799_, _42142_, _42141_);
  or (_42143_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42144_, \oc8051_gm_cxrom_1.cell8.data [0], _42138_);
  nand (_42145_, _42144_, _42143_);
  nand (_42146_, _42145_, _41894_);
  or (_42147_, \oc8051_gm_cxrom_1.cell8.data [0], _41894_);
  and (_01806_, _42147_, _42146_);
  or (_42148_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42149_, \oc8051_gm_cxrom_1.cell8.data [1], _42138_);
  nand (_42150_, _42149_, _42148_);
  nand (_42151_, _42150_, _41894_);
  or (_42152_, \oc8051_gm_cxrom_1.cell8.data [1], _41894_);
  and (_01810_, _42152_, _42151_);
  or (_42153_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42154_, \oc8051_gm_cxrom_1.cell8.data [2], _42138_);
  nand (_42155_, _42154_, _42153_);
  nand (_42156_, _42155_, _41894_);
  or (_42157_, \oc8051_gm_cxrom_1.cell8.data [2], _41894_);
  and (_01813_, _42157_, _42156_);
  or (_42158_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42159_, \oc8051_gm_cxrom_1.cell8.data [3], _42138_);
  nand (_42160_, _42159_, _42158_);
  nand (_42161_, _42160_, _41894_);
  or (_42162_, \oc8051_gm_cxrom_1.cell8.data [3], _41894_);
  and (_01817_, _42162_, _42161_);
  or (_42163_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42164_, \oc8051_gm_cxrom_1.cell8.data [4], _42138_);
  nand (_42165_, _42164_, _42163_);
  nand (_42166_, _42165_, _41894_);
  or (_42167_, \oc8051_gm_cxrom_1.cell8.data [4], _41894_);
  and (_01821_, _42167_, _42166_);
  or (_42168_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42169_, \oc8051_gm_cxrom_1.cell8.data [5], _42138_);
  nand (_42170_, _42169_, _42168_);
  nand (_42171_, _42170_, _41894_);
  or (_42172_, \oc8051_gm_cxrom_1.cell8.data [5], _41894_);
  and (_01825_, _42172_, _42171_);
  or (_42173_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42174_, \oc8051_gm_cxrom_1.cell8.data [6], _42138_);
  nand (_42175_, _42174_, _42173_);
  nand (_42176_, _42175_, _41894_);
  or (_42177_, \oc8051_gm_cxrom_1.cell8.data [6], _41894_);
  and (_01829_, _42177_, _42176_);
  or (_42178_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_42179_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_42180_, _42179_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_42181_, _42180_, _42178_);
  nand (_42182_, _42181_, _41894_);
  or (_42183_, \oc8051_gm_cxrom_1.cell9.data [7], _41894_);
  and (_01850_, _42183_, _42182_);
  or (_42184_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42185_, \oc8051_gm_cxrom_1.cell9.data [0], _42179_);
  nand (_42186_, _42185_, _42184_);
  nand (_42187_, _42186_, _41894_);
  or (_42188_, \oc8051_gm_cxrom_1.cell9.data [0], _41894_);
  and (_01857_, _42188_, _42187_);
  or (_42189_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42190_, \oc8051_gm_cxrom_1.cell9.data [1], _42179_);
  nand (_42191_, _42190_, _42189_);
  nand (_42192_, _42191_, _41894_);
  or (_42193_, \oc8051_gm_cxrom_1.cell9.data [1], _41894_);
  and (_01861_, _42193_, _42192_);
  or (_42194_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42195_, \oc8051_gm_cxrom_1.cell9.data [2], _42179_);
  nand (_42196_, _42195_, _42194_);
  nand (_42197_, _42196_, _41894_);
  or (_42198_, \oc8051_gm_cxrom_1.cell9.data [2], _41894_);
  and (_01865_, _42198_, _42197_);
  or (_42199_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42200_, \oc8051_gm_cxrom_1.cell9.data [3], _42179_);
  nand (_42201_, _42200_, _42199_);
  nand (_42202_, _42201_, _41894_);
  or (_42203_, \oc8051_gm_cxrom_1.cell9.data [3], _41894_);
  and (_01869_, _42203_, _42202_);
  or (_42204_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42205_, \oc8051_gm_cxrom_1.cell9.data [4], _42179_);
  nand (_42206_, _42205_, _42204_);
  nand (_42207_, _42206_, _41894_);
  or (_42208_, \oc8051_gm_cxrom_1.cell9.data [4], _41894_);
  and (_01873_, _42208_, _42207_);
  or (_42209_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42210_, \oc8051_gm_cxrom_1.cell9.data [5], _42179_);
  nand (_42211_, _42210_, _42209_);
  nand (_42212_, _42211_, _41894_);
  or (_42213_, \oc8051_gm_cxrom_1.cell9.data [5], _41894_);
  and (_01877_, _42213_, _42212_);
  or (_42214_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42215_, \oc8051_gm_cxrom_1.cell9.data [6], _42179_);
  nand (_42216_, _42215_, _42214_);
  nand (_42217_, _42216_, _41894_);
  or (_42218_, \oc8051_gm_cxrom_1.cell9.data [6], _41894_);
  and (_01881_, _42218_, _42217_);
  or (_42219_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_42220_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_42221_, _42220_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_42222_, _42221_, _42219_);
  nand (_42223_, _42222_, _41894_);
  or (_42224_, \oc8051_gm_cxrom_1.cell10.data [7], _41894_);
  and (_01889_, _42224_, _42223_);
  or (_42225_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42226_, \oc8051_gm_cxrom_1.cell10.data [0], _42220_);
  nand (_42227_, _42226_, _42225_);
  nand (_42228_, _42227_, _41894_);
  or (_42229_, \oc8051_gm_cxrom_1.cell10.data [0], _41894_);
  and (_01896_, _42229_, _42228_);
  or (_42230_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42231_, \oc8051_gm_cxrom_1.cell10.data [1], _42220_);
  nand (_42232_, _42231_, _42230_);
  nand (_42233_, _42232_, _41894_);
  or (_42234_, \oc8051_gm_cxrom_1.cell10.data [1], _41894_);
  and (_01900_, _42234_, _42233_);
  or (_42235_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42236_, \oc8051_gm_cxrom_1.cell10.data [2], _42220_);
  nand (_42237_, _42236_, _42235_);
  nand (_42238_, _42237_, _41894_);
  or (_42239_, \oc8051_gm_cxrom_1.cell10.data [2], _41894_);
  and (_01904_, _42239_, _42238_);
  or (_42240_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42241_, \oc8051_gm_cxrom_1.cell10.data [3], _42220_);
  nand (_42242_, _42241_, _42240_);
  nand (_42243_, _42242_, _41894_);
  or (_42244_, \oc8051_gm_cxrom_1.cell10.data [3], _41894_);
  and (_01908_, _42244_, _42243_);
  or (_42245_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42246_, \oc8051_gm_cxrom_1.cell10.data [4], _42220_);
  nand (_42247_, _42246_, _42245_);
  nand (_42248_, _42247_, _41894_);
  or (_42249_, \oc8051_gm_cxrom_1.cell10.data [4], _41894_);
  and (_01912_, _42249_, _42248_);
  or (_42250_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42251_, \oc8051_gm_cxrom_1.cell10.data [5], _42220_);
  nand (_42252_, _42251_, _42250_);
  nand (_42253_, _42252_, _41894_);
  or (_42254_, \oc8051_gm_cxrom_1.cell10.data [5], _41894_);
  and (_01916_, _42254_, _42253_);
  or (_42255_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42256_, \oc8051_gm_cxrom_1.cell10.data [6], _42220_);
  nand (_42257_, _42256_, _42255_);
  nand (_42258_, _42257_, _41894_);
  or (_42259_, \oc8051_gm_cxrom_1.cell10.data [6], _41894_);
  and (_01920_, _42259_, _42258_);
  or (_42260_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_42261_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_42262_, _42261_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_42263_, _42262_, _42260_);
  nand (_42264_, _42263_, _41894_);
  or (_42265_, \oc8051_gm_cxrom_1.cell11.data [7], _41894_);
  and (_01942_, _42265_, _42264_);
  or (_42266_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42267_, \oc8051_gm_cxrom_1.cell11.data [0], _42261_);
  nand (_42268_, _42267_, _42266_);
  nand (_42269_, _42268_, _41894_);
  or (_42270_, \oc8051_gm_cxrom_1.cell11.data [0], _41894_);
  and (_01949_, _42270_, _42269_);
  or (_42271_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42272_, \oc8051_gm_cxrom_1.cell11.data [1], _42261_);
  nand (_42273_, _42272_, _42271_);
  nand (_42274_, _42273_, _41894_);
  or (_42275_, \oc8051_gm_cxrom_1.cell11.data [1], _41894_);
  and (_01953_, _42275_, _42274_);
  or (_42276_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42277_, \oc8051_gm_cxrom_1.cell11.data [2], _42261_);
  nand (_42278_, _42277_, _42276_);
  nand (_42279_, _42278_, _41894_);
  or (_42280_, \oc8051_gm_cxrom_1.cell11.data [2], _41894_);
  and (_01957_, _42280_, _42279_);
  or (_42281_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42282_, \oc8051_gm_cxrom_1.cell11.data [3], _42261_);
  nand (_42283_, _42282_, _42281_);
  nand (_42284_, _42283_, _41894_);
  or (_42285_, \oc8051_gm_cxrom_1.cell11.data [3], _41894_);
  and (_01961_, _42285_, _42284_);
  or (_42286_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42287_, \oc8051_gm_cxrom_1.cell11.data [4], _42261_);
  nand (_42288_, _42287_, _42286_);
  nand (_42289_, _42288_, _41894_);
  or (_42290_, \oc8051_gm_cxrom_1.cell11.data [4], _41894_);
  and (_01965_, _42290_, _42289_);
  or (_42291_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42292_, \oc8051_gm_cxrom_1.cell11.data [5], _42261_);
  nand (_42293_, _42292_, _42291_);
  nand (_42294_, _42293_, _41894_);
  or (_42295_, \oc8051_gm_cxrom_1.cell11.data [5], _41894_);
  and (_01969_, _42295_, _42294_);
  or (_42296_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42297_, \oc8051_gm_cxrom_1.cell11.data [6], _42261_);
  nand (_42298_, _42297_, _42296_);
  nand (_42299_, _42298_, _41894_);
  or (_42300_, \oc8051_gm_cxrom_1.cell11.data [6], _41894_);
  and (_01973_, _42300_, _42299_);
  or (_42301_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_42302_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_42303_, _42302_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_42304_, _42303_, _42301_);
  nand (_42305_, _42304_, _41894_);
  or (_42306_, \oc8051_gm_cxrom_1.cell12.data [7], _41894_);
  and (_01995_, _42306_, _42305_);
  or (_42307_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42308_, \oc8051_gm_cxrom_1.cell12.data [0], _42302_);
  nand (_42309_, _42308_, _42307_);
  nand (_42310_, _42309_, _41894_);
  or (_42311_, \oc8051_gm_cxrom_1.cell12.data [0], _41894_);
  and (_02001_, _42311_, _42310_);
  or (_42312_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42313_, \oc8051_gm_cxrom_1.cell12.data [1], _42302_);
  nand (_42314_, _42313_, _42312_);
  nand (_42315_, _42314_, _41894_);
  or (_42316_, \oc8051_gm_cxrom_1.cell12.data [1], _41894_);
  and (_02005_, _42316_, _42315_);
  or (_42317_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42318_, \oc8051_gm_cxrom_1.cell12.data [2], _42302_);
  nand (_42319_, _42318_, _42317_);
  nand (_42320_, _42319_, _41894_);
  or (_42321_, \oc8051_gm_cxrom_1.cell12.data [2], _41894_);
  and (_02009_, _42321_, _42320_);
  or (_42322_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42323_, \oc8051_gm_cxrom_1.cell12.data [3], _42302_);
  nand (_42324_, _42323_, _42322_);
  nand (_42325_, _42324_, _41894_);
  or (_42326_, \oc8051_gm_cxrom_1.cell12.data [3], _41894_);
  and (_02013_, _42326_, _42325_);
  or (_42327_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42328_, \oc8051_gm_cxrom_1.cell12.data [4], _42302_);
  nand (_42329_, _42328_, _42327_);
  nand (_42330_, _42329_, _41894_);
  or (_42331_, \oc8051_gm_cxrom_1.cell12.data [4], _41894_);
  and (_02017_, _42331_, _42330_);
  or (_42332_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42333_, \oc8051_gm_cxrom_1.cell12.data [5], _42302_);
  nand (_42334_, _42333_, _42332_);
  nand (_42335_, _42334_, _41894_);
  or (_42336_, \oc8051_gm_cxrom_1.cell12.data [5], _41894_);
  and (_02021_, _42336_, _42335_);
  or (_42337_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42338_, \oc8051_gm_cxrom_1.cell12.data [6], _42302_);
  nand (_42339_, _42338_, _42337_);
  nand (_42340_, _42339_, _41894_);
  or (_42341_, \oc8051_gm_cxrom_1.cell12.data [6], _41894_);
  and (_02025_, _42341_, _42340_);
  or (_42342_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_42343_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_42344_, _42343_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_42345_, _42344_, _42342_);
  nand (_42346_, _42345_, _41894_);
  or (_42347_, \oc8051_gm_cxrom_1.cell13.data [7], _41894_);
  and (_02046_, _42347_, _42346_);
  or (_42348_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42349_, \oc8051_gm_cxrom_1.cell13.data [0], _42343_);
  nand (_42350_, _42349_, _42348_);
  nand (_42351_, _42350_, _41894_);
  or (_42352_, \oc8051_gm_cxrom_1.cell13.data [0], _41894_);
  and (_02053_, _42352_, _42351_);
  or (_42353_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42354_, \oc8051_gm_cxrom_1.cell13.data [1], _42343_);
  nand (_42355_, _42354_, _42353_);
  nand (_42356_, _42355_, _41894_);
  or (_42357_, \oc8051_gm_cxrom_1.cell13.data [1], _41894_);
  and (_02057_, _42357_, _42356_);
  or (_42358_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42359_, \oc8051_gm_cxrom_1.cell13.data [2], _42343_);
  nand (_42360_, _42359_, _42358_);
  nand (_42361_, _42360_, _41894_);
  or (_42362_, \oc8051_gm_cxrom_1.cell13.data [2], _41894_);
  and (_02061_, _42362_, _42361_);
  or (_42363_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42364_, \oc8051_gm_cxrom_1.cell13.data [3], _42343_);
  nand (_42365_, _42364_, _42363_);
  nand (_42366_, _42365_, _41894_);
  or (_42367_, \oc8051_gm_cxrom_1.cell13.data [3], _41894_);
  and (_02065_, _42367_, _42366_);
  or (_42368_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42369_, \oc8051_gm_cxrom_1.cell13.data [4], _42343_);
  nand (_42370_, _42369_, _42368_);
  nand (_42371_, _42370_, _41894_);
  or (_42372_, \oc8051_gm_cxrom_1.cell13.data [4], _41894_);
  and (_02069_, _42372_, _42371_);
  or (_42373_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42374_, \oc8051_gm_cxrom_1.cell13.data [5], _42343_);
  nand (_42375_, _42374_, _42373_);
  nand (_42376_, _42375_, _41894_);
  or (_42377_, \oc8051_gm_cxrom_1.cell13.data [5], _41894_);
  and (_02073_, _42377_, _42376_);
  or (_42378_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42379_, \oc8051_gm_cxrom_1.cell13.data [6], _42343_);
  nand (_42380_, _42379_, _42378_);
  nand (_42381_, _42380_, _41894_);
  or (_42382_, \oc8051_gm_cxrom_1.cell13.data [6], _41894_);
  and (_02076_, _42382_, _42381_);
  or (_42383_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_42384_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_42385_, _42384_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_42386_, _42385_, _42383_);
  nand (_42387_, _42386_, _41894_);
  or (_42388_, \oc8051_gm_cxrom_1.cell14.data [7], _41894_);
  and (_02098_, _42388_, _42387_);
  or (_42389_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42390_, \oc8051_gm_cxrom_1.cell14.data [0], _42384_);
  nand (_42391_, _42390_, _42389_);
  nand (_42392_, _42391_, _41894_);
  or (_42393_, \oc8051_gm_cxrom_1.cell14.data [0], _41894_);
  and (_02105_, _42393_, _42392_);
  or (_42394_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42395_, \oc8051_gm_cxrom_1.cell14.data [1], _42384_);
  nand (_42396_, _42395_, _42394_);
  nand (_42397_, _42396_, _41894_);
  or (_42398_, \oc8051_gm_cxrom_1.cell14.data [1], _41894_);
  and (_02109_, _42398_, _42397_);
  or (_42399_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42400_, \oc8051_gm_cxrom_1.cell14.data [2], _42384_);
  nand (_42401_, _42400_, _42399_);
  nand (_42402_, _42401_, _41894_);
  or (_42403_, \oc8051_gm_cxrom_1.cell14.data [2], _41894_);
  and (_02112_, _42403_, _42402_);
  or (_42404_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42405_, \oc8051_gm_cxrom_1.cell14.data [3], _42384_);
  nand (_42406_, _42405_, _42404_);
  nand (_42407_, _42406_, _41894_);
  or (_42408_, \oc8051_gm_cxrom_1.cell14.data [3], _41894_);
  and (_02116_, _42408_, _42407_);
  or (_42409_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42410_, \oc8051_gm_cxrom_1.cell14.data [4], _42384_);
  nand (_42411_, _42410_, _42409_);
  nand (_42412_, _42411_, _41894_);
  or (_42413_, \oc8051_gm_cxrom_1.cell14.data [4], _41894_);
  and (_02120_, _42413_, _42412_);
  or (_42414_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42415_, \oc8051_gm_cxrom_1.cell14.data [5], _42384_);
  nand (_42416_, _42415_, _42414_);
  nand (_42417_, _42416_, _41894_);
  or (_42418_, \oc8051_gm_cxrom_1.cell14.data [5], _41894_);
  and (_02124_, _42418_, _42417_);
  or (_42419_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42420_, \oc8051_gm_cxrom_1.cell14.data [6], _42384_);
  nand (_42421_, _42420_, _42419_);
  nand (_42422_, _42421_, _41894_);
  or (_42423_, \oc8051_gm_cxrom_1.cell14.data [6], _41894_);
  and (_02128_, _42423_, _42422_);
  or (_42424_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_42425_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_42426_, _42425_, \oc8051_gm_cxrom_1.cell15.data [7]);
  and (_42427_, _42426_, _42424_);
  or (_42428_, _42427_, rst);
  or (_42429_, \oc8051_gm_cxrom_1.cell15.data [7], _41894_);
  and (_02150_, _42429_, _42428_);
  or (_42430_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42431_, \oc8051_gm_cxrom_1.cell15.data [0], _42425_);
  and (_42432_, _42431_, _42430_);
  or (_42433_, _42432_, rst);
  or (_42434_, \oc8051_gm_cxrom_1.cell15.data [0], _41894_);
  and (_02157_, _42434_, _42433_);
  or (_42435_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42436_, \oc8051_gm_cxrom_1.cell15.data [1], _42425_);
  and (_42437_, _42436_, _42435_);
  or (_42438_, _42437_, rst);
  or (_42439_, \oc8051_gm_cxrom_1.cell15.data [1], _41894_);
  and (_02161_, _42439_, _42438_);
  or (_42440_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42441_, \oc8051_gm_cxrom_1.cell15.data [2], _42425_);
  and (_42442_, _42441_, _42440_);
  or (_42443_, _42442_, rst);
  or (_42444_, \oc8051_gm_cxrom_1.cell15.data [2], _41894_);
  and (_02164_, _42444_, _42443_);
  or (_42445_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42446_, \oc8051_gm_cxrom_1.cell15.data [3], _42425_);
  and (_42447_, _42446_, _42445_);
  or (_42448_, _42447_, rst);
  or (_42449_, \oc8051_gm_cxrom_1.cell15.data [3], _41894_);
  and (_02168_, _42449_, _42448_);
  or (_42450_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42451_, \oc8051_gm_cxrom_1.cell15.data [4], _42425_);
  and (_42452_, _42451_, _42450_);
  or (_42453_, _42452_, rst);
  or (_42454_, \oc8051_gm_cxrom_1.cell15.data [4], _41894_);
  and (_02172_, _42454_, _42453_);
  or (_42455_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42456_, \oc8051_gm_cxrom_1.cell15.data [5], _42425_);
  and (_42457_, _42456_, _42455_);
  or (_42458_, _42457_, rst);
  or (_42459_, \oc8051_gm_cxrom_1.cell15.data [5], _41894_);
  and (_02176_, _42459_, _42458_);
  or (_42460_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42461_, \oc8051_gm_cxrom_1.cell15.data [6], _42425_);
  and (_42462_, _42461_, _42460_);
  or (_42463_, _42462_, rst);
  or (_42464_, \oc8051_gm_cxrom_1.cell15.data [6], _41894_);
  and (_02180_, _42464_, _42463_);
  nor (_05948_, _36938_, rst);
  and (_42465_, _34358_, _41894_);
  nand (_42466_, _42465_, _37102_);
  nor (_42467_, _36807_, _36599_);
  or (_05951_, _42467_, _42466_);
  not (_42468_, _35243_);
  and (_42469_, _35489_, _42468_);
  not (_42470_, _34740_);
  and (_42471_, _42470_, _34991_);
  and (_42472_, _42471_, _42469_);
  not (_42473_, _35764_);
  nor (_42474_, _36039_, _42473_);
  and (_42475_, _36523_, _36281_);
  and (_42476_, _42475_, _42474_);
  and (_42477_, _42476_, _42472_);
  not (_42478_, _35489_);
  and (_42479_, _42478_, _35243_);
  and (_42480_, _42479_, _34740_);
  and (_42481_, _42480_, _42476_);
  not (_42482_, _36039_);
  not (_42483_, _36281_);
  nor (_42484_, _36523_, _42483_);
  and (_42485_, _42484_, _42482_);
  nor (_42486_, _42470_, _34991_);
  and (_42487_, _42486_, _42469_);
  and (_42488_, _42487_, _42485_);
  or (_42489_, _42488_, _42481_);
  or (_42490_, _42489_, _42477_);
  not (_42491_, _34991_);
  nor (_42492_, _35489_, _35243_);
  and (_42493_, _42492_, _42491_);
  and (_42494_, _42493_, _42476_);
  and (_42495_, _42475_, _36039_);
  and (_42496_, _42492_, _42486_);
  and (_42497_, _42496_, _42495_);
  or (_42498_, _42497_, _42494_);
  nor (_42499_, _34740_, _34991_);
  and (_42500_, _42499_, _42492_);
  and (_42501_, _42500_, _42495_);
  and (_42502_, _34740_, _34991_);
  and (_42503_, _42492_, _42502_);
  and (_42504_, _42503_, _42483_);
  or (_42505_, _42504_, _42501_);
  or (_42506_, _42505_, _42498_);
  or (_42507_, _42506_, _42490_);
  and (_42508_, _42484_, _42474_);
  and (_42509_, _42508_, _42470_);
  and (_42510_, _42509_, _42469_);
  and (_42511_, _42499_, _42479_);
  nor (_42512_, _42511_, _42473_);
  not (_42513_, _42512_);
  and (_42514_, _42475_, _42482_);
  and (_42515_, _42514_, _42513_);
  not (_42516_, _42515_);
  and (_42517_, _35489_, _35243_);
  and (_42518_, _42517_, _42486_);
  and (_42519_, _42518_, _42476_);
  and (_42520_, _42479_, _42471_);
  and (_42521_, _42520_, _42476_);
  nor (_42522_, _42521_, _42519_);
  and (_42523_, _42522_, _42516_);
  not (_42524_, _42523_);
  or (_42525_, _42524_, _42510_);
  or (_42526_, _42525_, _42507_);
  nor (_42527_, _42499_, _42502_);
  not (_42528_, _42527_);
  and (_42529_, _42517_, _42476_);
  and (_42530_, _42529_, _42528_);
  and (_42531_, _42485_, _42473_);
  and (_42532_, _42531_, _42503_);
  and (_42533_, _42517_, _42491_);
  and (_42534_, _42495_, _35764_);
  and (_42535_, _42534_, _42533_);
  or (_42536_, _42535_, _42532_);
  or (_42537_, _42536_, _42530_);
  and (_42538_, _42486_, _42479_);
  and (_42539_, _42495_, _42473_);
  nand (_42540_, _42539_, _42538_);
  and (_42541_, _42469_, _42491_);
  and (_42542_, _34740_, _36039_);
  and (_42543_, _42542_, _42484_);
  and (_42544_, _42543_, _42541_);
  and (_42545_, _42487_, _42483_);
  nor (_42546_, _42545_, _42544_);
  nand (_42547_, _42546_, _42540_);
  and (_42548_, _42469_, _34991_);
  and (_42549_, _42539_, _42548_);
  and (_42550_, _42517_, _34991_);
  and (_42551_, _42550_, _42534_);
  or (_42552_, _42551_, _42549_);
  or (_42553_, _42552_, _42547_);
  or (_42554_, _42553_, _42537_);
  or (_42555_, _42554_, _42526_);
  and (_42556_, _42555_, _34369_);
  not (_42557_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_42558_, _34347_, _16097_);
  and (_42559_, _42558_, _36752_);
  nor (_42560_, _42559_, _42557_);
  or (_42561_, _42560_, rst);
  or (_05954_, _42561_, _42556_);
  nand (_42562_, _35243_, _34303_);
  or (_42563_, _34303_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_42564_, _42563_, _41894_);
  and (_05957_, _42564_, _42562_);
  and (_42565_, \oc8051_top_1.oc8051_sfr1.wait_data , _41894_);
  and (_42566_, _42565_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_42567_, _36610_, _36851_);
  and (_42568_, _36884_, _37113_);
  or (_42569_, _42568_, _42567_);
  and (_42570_, _36851_, _36807_);
  or (_42571_, _42570_, _36818_);
  or (_42572_, _42571_, _37593_);
  and (_42573_, _36610_, _37244_);
  and (_42574_, _37494_, _36599_);
  or (_42575_, _42574_, _42573_);
  nor (_42576_, _42575_, _42572_);
  nand (_42577_, _42576_, _37731_);
  or (_42578_, _42577_, _42569_);
  and (_42579_, _42578_, _42465_);
  or (_05960_, _42579_, _42566_);
  and (_42580_, _36884_, _37244_);
  or (_42581_, _42580_, _37254_);
  and (_42582_, _36807_, _36654_);
  or (_42583_, _42582_, _36621_);
  and (_42584_, _37309_, _37167_);
  or (_42585_, _42584_, _38138_);
  or (_42586_, _42585_, _42583_);
  or (_42587_, _42586_, _42581_);
  and (_42588_, _42587_, _34358_);
  and (_42589_, \oc8051_top_1.oc8051_decoder1.state [0], _16097_);
  and (_42590_, _42589_, _42557_);
  not (_42591_, _36916_);
  and (_42592_, _42591_, _42590_);
  and (_42593_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42594_, _42593_, _42592_);
  or (_42595_, _42594_, _42588_);
  and (_05963_, _42595_, _41894_);
  and (_42596_, _42565_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_42597_, _38270_);
  and (_42598_, _36884_, _37342_);
  or (_42599_, _37505_, _37353_);
  or (_42600_, _42599_, _42598_);
  and (_42601_, _37331_, _37309_);
  nor (_42602_, _34794_, _36325_);
  and (_42603_, _42602_, _37156_);
  and (_42604_, _42603_, _35298_);
  or (_42605_, _42604_, _42601_);
  and (_42606_, _42602_, _37331_);
  or (_42607_, _42606_, _42605_);
  and (_42608_, _36873_, _36083_);
  and (_42609_, _42608_, _37488_);
  or (_42610_, _42609_, _42607_);
  or (_42611_, _42610_, _42600_);
  or (_42612_, _42611_, _42597_);
  and (_42613_, _42602_, _35555_);
  and (_42614_, _36884_, _37069_);
  or (_42615_, _42614_, _42613_);
  or (_42616_, _42615_, _42583_);
  or (_42617_, _42616_, _42612_);
  and (_42618_, _42617_, _42465_);
  or (_05966_, _42618_, _42596_);
  and (_42619_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42620_, _37458_, _34358_);
  or (_42621_, _42620_, _42619_);
  or (_42622_, _42621_, _42592_);
  and (_05969_, _42622_, _41894_);
  and (_42623_, _36610_, _36643_);
  not (_42624_, _37113_);
  nor (_42625_, _42467_, _42624_);
  nor (_42626_, _42625_, _42623_);
  not (_42627_, _42626_);
  and (_42628_, _42627_, _42590_);
  or (_42629_, _42628_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42630_, _37488_, _36982_);
  and (_42631_, _37036_, _36577_);
  and (_42632_, _42631_, _36632_);
  or (_42633_, _42632_, _42630_);
  not (_42634_, _34314_);
  and (_42635_, _42567_, _42634_);
  or (_42636_, _42635_, _42633_);
  and (_42637_, _42636_, _36752_);
  or (_42638_, _42637_, _42629_);
  or (_42639_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _16097_);
  and (_42640_, _42639_, _41894_);
  and (_05972_, _42640_, _42638_);
  and (_42641_, _42565_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_42642_, _36325_);
  and (_42643_, _37488_, _42642_);
  and (_42644_, _37494_, _42642_);
  or (_42645_, _42644_, _42643_);
  or (_42646_, _36621_, _37505_);
  or (_42647_, _42646_, _42645_);
  and (_42648_, _38138_, _34794_);
  or (_42649_, _42574_, _37775_);
  or (_42650_, _42649_, _42648_);
  or (_42651_, _42584_, _37254_);
  and (_42652_, _37331_, _38072_);
  or (_42653_, _42609_, _42652_);
  or (_42654_, _42653_, _37582_);
  or (_42655_, _42654_, _42651_);
  or (_42656_, _42655_, _42650_);
  or (_42657_, _42656_, _42647_);
  and (_42658_, _42657_, _42465_);
  or (_05975_, _42658_, _42641_);
  and (_42659_, _42565_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  not (_42660_, _37637_);
  and (_42661_, _36884_, _37538_);
  or (_42662_, _42661_, _42660_);
  and (_42663_, _42608_, _37244_);
  and (_42664_, _37309_, _37156_);
  and (_42665_, _37309_, _36675_);
  or (_42666_, _42665_, _42664_);
  or (_42667_, _42666_, _42663_);
  and (_42668_, _36610_, _36993_);
  nor (_42669_, _38248_, _37145_);
  not (_42670_, _42669_);
  or (_42671_, _42670_, _42668_);
  or (_42672_, _42671_, _42667_);
  and (_42673_, _38072_, _37167_);
  and (_42674_, _38017_, _37156_);
  or (_42675_, _38171_, _42674_);
  or (_42676_, _42675_, _42673_);
  not (_42677_, _37560_);
  and (_42678_, _42608_, _37135_);
  or (_42679_, _42678_, _42677_);
  or (_42680_, _42679_, _42676_);
  or (_42681_, _42680_, _42672_);
  or (_42682_, _42681_, _42662_);
  or (_42683_, _42682_, _42611_);
  and (_42684_, _42683_, _42465_);
  or (_05978_, _42684_, _42659_);
  and (_42685_, _42602_, _36643_);
  and (_42686_, _36873_, _37004_);
  or (_42687_, _42686_, _42685_);
  and (_42688_, _37004_, _42642_);
  or (_42689_, _42688_, _38127_);
  or (_42690_, _42689_, _42687_);
  and (_42691_, _42608_, _36654_);
  or (_42692_, _42691_, _42591_);
  or (_42693_, _42692_, _42690_);
  and (_42694_, _42693_, _42465_);
  nor (_42695_, _36916_, _42634_);
  and (_42696_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_42697_, _42696_, _42695_);
  and (_42698_, _42697_, _41894_);
  or (_05981_, _42698_, _42694_);
  nand (_42699_, _37604_, _37466_);
  or (_42700_, _37786_, _37254_);
  or (_42701_, _42700_, _42599_);
  or (_42702_, _42701_, _42699_);
  and (_42703_, _36632_, _37047_);
  and (_42704_, _42703_, _36665_);
  or (_42705_, _42630_, _37200_);
  or (_42706_, _42705_, _42704_);
  or (_42707_, _37626_, _37489_);
  or (_42708_, _42707_, _42632_);
  and (_42709_, _37309_, _36643_);
  or (_42710_, _42709_, _38160_);
  or (_42711_, _42710_, _37753_);
  or (_42712_, _42711_, _42708_);
  or (_42713_, _42712_, _42706_);
  or (_42714_, _42713_, _42702_);
  and (_42715_, _38072_, _36665_);
  not (_42716_, _38248_);
  nand (_42717_, _42716_, _37298_);
  or (_42718_, _42717_, _42715_);
  and (_42719_, _42602_, _36665_);
  or (_42720_, _42719_, _37320_);
  or (_42721_, _42720_, _42585_);
  or (_42722_, _42721_, _42718_);
  or (_42723_, _42722_, _42607_);
  or (_42724_, _42723_, _42714_);
  and (_42725_, _42724_, _34358_);
  and (_42726_, _42633_, _36774_);
  or (_42727_, _42726_, _42592_);
  and (_42728_, _36774_, _37863_);
  or (_42729_, _42728_, _42727_);
  and (_42730_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42731_, _42730_, _42729_);
  or (_42732_, _42731_, _42725_);
  and (_05984_, _42732_, _41894_);
  nor (_06043_, _38368_, rst);
  nor (_06045_, _37962_, rst);
  nand (_06048_, _42627_, _42465_);
  and (_42733_, _36807_, _37102_);
  or (_42734_, _42733_, _42623_);
  nand (_06051_, _42734_, _42465_);
  or (_42735_, _42549_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_42736_, _42735_, _42535_);
  or (_42737_, _42736_, _42510_);
  and (_42738_, _42737_, _42559_);
  nor (_42739_, _42558_, _36752_);
  or (_42740_, _42739_, rst);
  or (_06054_, _42740_, _42738_);
  nand (_42741_, _35764_, _34303_);
  or (_42742_, _34303_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_42743_, _42742_, _41894_);
  and (_06057_, _42743_, _42741_);
  not (_42744_, _34303_);
  or (_42745_, _36039_, _42744_);
  or (_42746_, _34303_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_42747_, _42746_, _41894_);
  and (_06060_, _42747_, _42745_);
  nand (_42748_, _36523_, _34303_);
  or (_42749_, _34303_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_42750_, _42749_, _41894_);
  and (_06063_, _42750_, _42748_);
  nand (_42751_, _36281_, _34303_);
  or (_42752_, _34303_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_42753_, _42752_, _41894_);
  and (_06066_, _42753_, _42751_);
  or (_42754_, _34740_, _42744_);
  or (_42755_, _34303_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_42756_, _42755_, _41894_);
  and (_06069_, _42756_, _42754_);
  nand (_42757_, _34991_, _34303_);
  or (_42758_, _34303_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_42759_, _42758_, _41894_);
  and (_06072_, _42759_, _42757_);
  nand (_42760_, _35489_, _34303_);
  or (_42761_, _34303_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_42762_, _42761_, _41894_);
  and (_06075_, _42762_, _42760_);
  or (_42763_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _16097_);
  and (_42764_, _42763_, _42629_);
  nor (_42765_, _37427_, _36325_);
  or (_42766_, _37494_, _37331_);
  and (_42767_, _42766_, _36884_);
  or (_42768_, _42767_, _42687_);
  or (_42769_, _42768_, _42765_);
  or (_42770_, _38171_, _38127_);
  or (_42771_, _42678_, _42665_);
  or (_42772_, _42771_, _42770_);
  or (_42773_, _36621_, _37124_);
  or (_42774_, _42773_, _42772_);
  and (_42775_, _37309_, _37102_);
  and (_42776_, _42664_, _35287_);
  or (_42777_, _42691_, _42776_);
  nor (_42778_, _42777_, _42775_);
  nand (_42779_, _42778_, _38050_);
  or (_42780_, _42779_, _42774_);
  and (_42781_, _42608_, _37419_);
  and (_42782_, _36884_, _36686_);
  or (_42783_, _42782_, _38083_);
  or (_42784_, _42783_, _42781_);
  or (_42785_, _42668_, _42568_);
  and (_42786_, _37102_, _36632_);
  and (_42787_, _42786_, _36884_);
  and (_42788_, _42608_, _37538_);
  or (_42789_, _42788_, _42582_);
  or (_42790_, _42789_, _42787_);
  or (_42791_, _42790_, _42785_);
  or (_42792_, _42791_, _42784_);
  or (_42793_, _42792_, _42780_);
  or (_42794_, _42793_, _42769_);
  and (_42795_, _42794_, _34358_);
  or (_42796_, _42795_, _42764_);
  and (_30379_, _42796_, _41894_);
  and (_42797_, _42565_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not (_42798_, _37427_);
  and (_42799_, _36884_, _42798_);
  or (_42800_, _42799_, _42676_);
  and (_42801_, _36884_, _37135_);
  nor (_42802_, _42801_, _42614_);
  nand (_42803_, _42802_, _37265_);
  or (_42804_, _42803_, _42800_);
  or (_42805_, _42789_, _42666_);
  nor (_42806_, _42613_, _38259_);
  and (_42807_, _36785_, _34794_);
  nand (_42808_, _42807_, _36982_);
  nand (_42809_, _42808_, _42806_);
  or (_42810_, _42809_, _42805_);
  or (_42812_, _42810_, _42569_);
  or (_42814_, _42812_, _42804_);
  and (_42816_, _42814_, _42465_);
  or (_30382_, _42816_, _42797_);
  and (_42819_, _42714_, _34358_);
  and (_42821_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42823_, _42821_, _42729_);
  or (_42825_, _42823_, _42819_);
  and (_30384_, _42825_, _41894_);
  and (_42828_, _37178_, _34794_);
  or (_42830_, _42828_, _38138_);
  or (_42832_, _42830_, _42718_);
  or (_42834_, _42832_, _42633_);
  and (_42836_, _42834_, _34358_);
  and (_42838_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42840_, _42838_, _42727_);
  or (_42842_, _42840_, _42836_);
  and (_30386_, _42842_, _41894_);
  and (_42845_, _37419_, _36982_);
  and (_42847_, _36610_, _36686_);
  and (_42849_, _42703_, _37102_);
  or (_42851_, _42849_, _42847_);
  or (_42853_, _42851_, _42845_);
  or (_42855_, _42715_, _42661_);
  and (_42857_, _42608_, _37670_);
  or (_42859_, _42857_, _42801_);
  or (_42861_, _42859_, _42855_);
  or (_42863_, _42719_, _38127_);
  or (_42865_, _42863_, _42782_);
  or (_42867_, _42865_, _42861_);
  or (_42869_, _42867_, _42853_);
  and (_42870_, _42608_, _37698_);
  or (_42871_, _42870_, _42623_);
  or (_42872_, _42781_, _36906_);
  or (_42873_, _42872_, _42871_);
  or (_42874_, _42873_, _42633_);
  or (_42875_, _42874_, _42869_);
  or (_42876_, _42691_, _36895_);
  or (_42877_, _42876_, _42787_);
  or (_42878_, _42877_, _42580_);
  and (_42879_, _42608_, _37058_);
  or (_42880_, _42879_, _42568_);
  or (_42881_, _42880_, _42767_);
  or (_42882_, _42881_, _42878_);
  or (_42883_, _42685_, _42668_);
  or (_42884_, _42883_, _38105_);
  or (_42885_, _42884_, _42765_);
  or (_42886_, _42885_, _42882_);
  or (_42887_, _42886_, _42875_);
  and (_42888_, _42887_, _34358_);
  and (_42889_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42890_, _42628_, _42695_);
  or (_42891_, _42890_, _42889_);
  or (_42892_, _42891_, _42888_);
  and (_30388_, _42892_, _41894_);
  or (_42893_, _36697_, _37135_);
  and (_42894_, _42893_, _36610_);
  or (_42895_, _36906_, _38127_);
  or (_42896_, _42895_, _37753_);
  and (_42897_, _37626_, _35819_);
  or (_42898_, _42897_, _42704_);
  or (_42899_, _42898_, _42896_);
  and (_42900_, _42602_, _37102_);
  and (_42901_, _38072_, _37102_);
  or (_42902_, _42901_, _42582_);
  or (_42903_, _42902_, _42900_);
  or (_42904_, _42903_, _37435_);
  or (_42905_, _42904_, _42899_);
  or (_42906_, _42905_, _42894_);
  or (_42907_, _42906_, _42886_);
  and (_42908_, _42907_, _34358_);
  and (_42909_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42910_, _42909_, _42890_);
  or (_42911_, _42910_, _42908_);
  and (_30390_, _42911_, _41894_);
  and (_42912_, _42565_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_42913_, _40416_);
  or (_42914_, _42691_, _42913_);
  and (_42915_, _36610_, _37331_);
  and (_42916_, _42915_, _36632_);
  and (_42917_, _42574_, _35819_);
  or (_42918_, _42917_, _42916_);
  or (_42919_, _42918_, _42647_);
  or (_42920_, _42919_, _42914_);
  and (_42921_, _36884_, _37494_);
  or (_42922_, _42921_, _42609_);
  not (_42923_, _40414_);
  or (_42924_, _42700_, _42923_);
  or (_42925_, _42924_, _42922_);
  or (_42926_, _42685_, _42584_);
  and (_42927_, _36610_, _37698_);
  and (_42928_, _36610_, _37058_);
  or (_42929_, _42928_, _42927_);
  or (_42930_, _42929_, _42926_);
  and (_42931_, _42602_, _37004_);
  or (_42932_, _42931_, _38127_);
  and (_42933_, _38072_, _36993_);
  or (_42934_, _42933_, _42870_);
  or (_42935_, _42934_, _42932_);
  or (_42936_, _42648_, _37450_);
  or (_42937_, _42936_, _42935_);
  or (_42938_, _42937_, _42930_);
  or (_42939_, _42938_, _42925_);
  or (_42940_, _42939_, _42920_);
  and (_42941_, _42940_, _42465_);
  or (_30392_, _42941_, _42912_);
  or (_42942_, _42921_, _42927_);
  or (_42943_, _42942_, _42916_);
  not (_42944_, _37764_);
  or (_42945_, _42765_, _42944_);
  or (_42946_, _42945_, _42943_);
  or (_42948_, _42873_, _42662_);
  or (_42949_, _42857_, _42674_);
  or (_42950_, _42949_, _42581_);
  or (_42951_, _42664_, _42673_);
  or (_42952_, _42951_, _36621_);
  or (_42953_, _42847_, _37549_);
  or (_42954_, _42953_, _42952_);
  or (_42955_, _42954_, _38105_);
  or (_42956_, _42955_, _42950_);
  or (_42957_, _42956_, _42948_);
  or (_42958_, _42957_, _42946_);
  and (_42960_, _42958_, _42465_);
  and (_42961_, _34314_, _41894_);
  and (_42962_, _42961_, _36906_);
  and (_42963_, _42565_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_42964_, _42963_, _42962_);
  or (_30394_, _42964_, _42960_);
  and (_42965_, _42602_, _37408_);
  or (_42966_, _42965_, _38083_);
  and (_42967_, _36610_, _37004_);
  and (_42968_, _37058_, _36599_);
  or (_42969_, _42968_, _42787_);
  or (_42970_, _42969_, _42967_);
  or (_42971_, _42970_, _42966_);
  not (_42972_, _42781_);
  and (_42973_, _42972_, _37764_);
  and (_42974_, _37527_, _34794_);
  or (_42975_, _42663_, _42974_);
  or (_42976_, _42975_, _42926_);
  nor (_42977_, _42691_, _42613_);
  nand (_42978_, _42977_, _38149_);
  or (_42979_, _42978_, _42880_);
  nor (_42980_, _42979_, _42976_);
  nand (_42981_, _42980_, _42973_);
  or (_42982_, _42981_, _42971_);
  or (_42983_, _42982_, _42612_);
  and (_42984_, _42983_, _34358_);
  and (_42985_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42986_, _36906_, _16097_);
  or (_42987_, _42986_, _42985_);
  or (_42988_, _42987_, _42984_);
  and (_30396_, _42988_, _41894_);
  or (_42989_, _42969_, _42922_);
  or (_42990_, _42989_, _42966_);
  or (_42991_, _38248_, _38138_);
  or (_42992_, _42991_, _37753_);
  or (_42993_, _42915_, _42781_);
  or (_42994_, _42993_, _42992_);
  or (_42995_, _42651_, _42913_);
  or (_42996_, _42995_, _42994_);
  or (_42997_, _42607_, _42600_);
  or (_42998_, _42997_, _42996_);
  or (_42999_, _42998_, _42990_);
  and (_43000_, _42999_, _34358_);
  and (_43001_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_43002_, _36895_, _16097_);
  or (_43003_, _43002_, _43001_);
  or (_43004_, _43003_, _43000_);
  and (_30398_, _43004_, _41894_);
  and (_43005_, _42565_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_43006_, _42573_, _37775_);
  nand (_43007_, _43006_, _40414_);
  or (_43008_, _36610_, _36588_);
  and (_43009_, _43008_, _37058_);
  or (_43010_, _43009_, _42942_);
  or (_43011_, _43010_, _43007_);
  or (_43012_, _42918_, _42690_);
  or (_43013_, _43012_, _42914_);
  or (_43014_, _43013_, _43011_);
  and (_43015_, _43014_, _42465_);
  or (_30400_, _43015_, _43005_);
  nor (_38864_, _35243_, rst);
  nor (_38866_, _40405_, rst);
  and (_43016_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_43017_, _34478_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_43018_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_43019_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_43020_, _43019_, _43018_);
  and (_43021_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_43022_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_43023_, _43022_, _43021_);
  and (_43024_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_43025_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_43026_, _43025_, _43024_);
  and (_43027_, _43026_, _43023_);
  and (_43028_, _43027_, _43020_);
  nor (_43029_, _43028_, _34478_);
  nor (_43030_, _43029_, _43017_);
  nor (_43031_, _43030_, _40389_);
  nor (_43032_, _43031_, _43016_);
  nor (_38867_, _43032_, rst);
  nor (_38879_, _35764_, rst);
  and (_38880_, _36039_, _41894_);
  nor (_38881_, _36523_, rst);
  nor (_38882_, _36281_, rst);
  and (_38883_, _34740_, _41894_);
  nor (_38884_, _34991_, rst);
  nor (_38885_, _35489_, rst);
  nor (_38886_, _40568_, rst);
  nor (_38888_, _40736_, rst);
  nor (_38889_, _40485_, rst);
  nor (_38890_, _40530_, rst);
  nor (_38891_, _40663_, rst);
  nor (_38892_, _40442_, rst);
  nor (_38894_, _40624_, rst);
  and (_43033_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_43034_, _34478_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_43035_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_43036_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_43037_, _43036_, _43035_);
  and (_43038_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_43039_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_43040_, _43039_, _43038_);
  and (_43041_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_43042_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_43043_, _43042_, _43041_);
  and (_43044_, _43043_, _43040_);
  and (_43045_, _43044_, _43037_);
  nor (_43046_, _43045_, _34478_);
  nor (_43047_, _43046_, _43034_);
  nor (_43048_, _43047_, _40389_);
  nor (_43049_, _43048_, _43033_);
  nor (_38895_, _43049_, rst);
  and (_43050_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_43051_, _34478_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_43052_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_43053_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_43054_, _43053_, _43052_);
  and (_43055_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_43056_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_43057_, _43056_, _43055_);
  and (_43058_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_43059_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_43060_, _43059_, _43058_);
  and (_43061_, _43060_, _43057_);
  and (_43062_, _43061_, _43054_);
  nor (_43063_, _43062_, _34478_);
  nor (_43064_, _43063_, _43051_);
  nor (_43065_, _43064_, _40389_);
  nor (_43066_, _43065_, _43050_);
  nor (_38896_, _43066_, rst);
  and (_43067_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_43068_, _34478_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_43069_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_43070_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_43071_, _43070_, _43069_);
  and (_43072_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_43073_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_43074_, _43073_, _43072_);
  and (_43075_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_43076_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_43077_, _43076_, _43075_);
  and (_43078_, _43077_, _43074_);
  and (_43079_, _43078_, _43071_);
  nor (_43080_, _43079_, _34478_);
  nor (_43081_, _43080_, _43068_);
  nor (_43082_, _43081_, _40389_);
  nor (_43083_, _43082_, _43067_);
  nor (_38897_, _43083_, rst);
  and (_43084_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_43085_, _34478_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_43086_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_43087_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_43088_, _43087_, _43086_);
  and (_43089_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_43090_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_43091_, _43090_, _43089_);
  and (_43092_, _43091_, _43088_);
  and (_43093_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_43094_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_43095_, _43094_, _43093_);
  and (_43096_, _43095_, _43092_);
  nor (_43097_, _43096_, _34478_);
  nor (_43098_, _43097_, _43085_);
  nor (_43099_, _43098_, _40389_);
  nor (_43100_, _43099_, _43084_);
  nor (_38898_, _43100_, rst);
  and (_43101_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_43102_, _34478_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_43103_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_43104_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_43105_, _43104_, _43103_);
  and (_43106_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_43107_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_43108_, _43107_, _43106_);
  and (_43109_, _43108_, _43105_);
  and (_43110_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_43111_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_43112_, _43111_, _43110_);
  and (_43113_, _43112_, _43109_);
  nor (_43114_, _43113_, _34478_);
  nor (_43115_, _43114_, _43102_);
  nor (_43116_, _43115_, _40389_);
  nor (_43117_, _43116_, _43101_);
  nor (_38900_, _43117_, rst);
  and (_43118_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_43119_, _34478_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_43120_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_43121_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_43122_, _43121_, _43120_);
  and (_43123_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_43124_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_43125_, _43124_, _43123_);
  and (_43126_, _43125_, _43122_);
  and (_43127_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_43128_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_43129_, _43128_, _43127_);
  and (_43130_, _43129_, _43126_);
  nor (_43131_, _43130_, _34478_);
  nor (_43132_, _43131_, _43119_);
  nor (_43133_, _43132_, _40389_);
  nor (_43134_, _43133_, _43118_);
  nor (_38901_, _43134_, rst);
  and (_43135_, _40389_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_43136_, _34478_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_43137_, _34413_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_43138_, _34576_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_43139_, _43138_, _43137_);
  and (_43140_, _34445_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_43141_, _34511_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_43142_, _43141_, _43140_);
  and (_43143_, _43142_, _43139_);
  and (_43144_, _34631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_43145_, _34609_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_43146_, _43145_, _43144_);
  and (_43147_, _43146_, _43143_);
  nor (_43148_, _43147_, _34478_);
  nor (_43149_, _43148_, _43136_);
  nor (_43150_, _43149_, _40389_);
  nor (_43151_, _43150_, _43135_);
  nor (_38902_, _43151_, rst);
  and (_43152_, _34369_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_43153_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_43154_, _43152_, _38667_);
  and (_43155_, _43154_, _41894_);
  and (_38923_, _43155_, _43153_);
  not (_43156_, _43152_);
  or (_43157_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _43152_, _41894_);
  and (_43158_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _41894_);
  or (_43159_, _43158_, _00000_);
  and (_38924_, _43159_, _43157_);
  nor (_38959_, _40410_, rst);
  nor (_38961_, _40647_, rst);
  nor (_38962_, _40383_, rst);
  nor (_43160_, _40410_, _25406_);
  and (_43161_, _40410_, _25406_);
  nor (_43162_, _43161_, _43160_);
  nor (_43163_, _40550_, _25558_);
  and (_43164_, _40550_, _25558_);
  nor (_43165_, _43164_, _43163_);
  and (_43166_, _40682_, _38443_);
  nor (_43167_, _40682_, _38443_);
  nor (_43168_, _43167_, _43166_);
  and (_43169_, _43168_, _43165_);
  nor (_43170_, _40467_, _39112_);
  and (_43171_, _40467_, _39112_);
  or (_43172_, _43171_, _43170_);
  and (_43173_, _40632_, _38955_);
  nor (_43174_, _40632_, _38955_);
  or (_43175_, _43174_, _43173_);
  nor (_43176_, _43175_, _43172_);
  and (_43177_, _43176_, _43169_);
  and (_43178_, _43177_, _43162_);
  nor (_43179_, _37731_, _42589_);
  and (_43180_, _38938_, _28573_);
  and (_43181_, _43180_, _43179_);
  and (_43182_, _43181_, _43178_);
  nor (_43183_, _42570_, _42847_);
  and (_43184_, _30752_, _26478_);
  nand (_43185_, _43184_, _31374_);
  nor (_43186_, _43185_, _32105_);
  and (_43187_, _43186_, _32921_);
  and (_43188_, _43187_, _33607_);
  and (_43189_, _43188_, _27092_);
  not (_43190_, _37681_);
  and (_43191_, _40423_, _43190_);
  nor (_43192_, _43191_, _42589_);
  nor (_43193_, _43192_, _36829_);
  and (_43194_, _43193_, _29559_);
  and (_43195_, _43194_, _43189_);
  and (_43196_, _43179_, _26840_);
  nor (_43197_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_43198_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_43199_, _43198_, _43197_);
  nor (_43200_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_43201_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_43202_, _43201_, _43200_);
  and (_43203_, _43202_, _43199_);
  and (_43204_, _43203_, _38346_);
  nor (_43205_, _43179_, _35034_);
  nor (_43206_, _43205_, _36840_);
  and (_43207_, _43206_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_43208_, _43207_, _43204_);
  or (_43209_, _43208_, _43196_);
  nor (_43210_, _43209_, _43195_);
  and (_43211_, _36818_, _34794_);
  not (_43212_, _43211_);
  and (_43213_, _43212_, _37874_);
  nor (_43215_, _43213_, _43210_);
  or (_43216_, _37698_, _36686_);
  nor (_43217_, _43216_, _37419_);
  nor (_43218_, _43217_, _37692_);
  not (_43219_, _43218_);
  not (_43221_, _42644_);
  nor (_43222_, _42879_, _37505_);
  and (_43223_, _43222_, _43221_);
  and (_43224_, _43223_, _42806_);
  and (_43225_, _43224_, _43219_);
  not (_43227_, _43225_);
  and (_43228_, _43227_, _43210_);
  nor (_43229_, _43228_, _43215_);
  and (_43230_, _43229_, _43183_);
  nor (_43231_, _43230_, _37885_);
  and (_43233_, _37331_, _36982_);
  nor (_43234_, _43233_, _42631_);
  nor (_43235_, _43234_, _34314_);
  nor (_43236_, _43235_, _37918_);
  not (_43237_, _43236_);
  nor (_43239_, _43237_, _43231_);
  not (_43240_, _39174_);
  and (_43241_, _43240_, _38346_);
  nor (_43242_, _38958_, _38945_);
  and (_43243_, _43242_, _38953_);
  not (_43245_, _43243_);
  and (_43246_, _43245_, _43206_);
  nor (_43247_, _43246_, _43241_);
  not (_43248_, _43247_);
  nor (_43249_, _43248_, _43239_);
  not (_43251_, _43249_);
  nor (_43252_, _43251_, _43182_);
  and (_43254_, _40778_, _31178_);
  nor (_43255_, _40778_, _31178_);
  or (_43256_, _43255_, _43254_);
  not (_43257_, _43256_);
  nor (_43258_, _40586_, _24884_);
  and (_43259_, _40586_, _24884_);
  nor (_43260_, _43259_, _43258_);
  not (_43262_, _43260_);
  nor (_43263_, _40506_, _24644_);
  and (_43264_, _40506_, _24644_);
  nor (_43266_, _43264_, _43263_);
  nor (_43267_, _43266_, _39234_);
  and (_43268_, _43267_, _43262_);
  and (_43270_, _43268_, _43257_);
  and (_43271_, _43270_, _43178_);
  nor (_43272_, _25395_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_43274_, _43272_, _43271_);
  not (_43275_, _43274_);
  and (_43276_, _43275_, _43252_);
  nor (_43278_, _37929_, rst);
  and (_38966_, _43278_, _43276_);
  and (_38967_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _41894_);
  and (_38968_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _41894_);
  nor (_43280_, _37940_, _28496_);
  and (_43281_, _42847_, _36774_);
  not (_43283_, _43281_);
  nor (_43284_, _43283_, _38678_);
  and (_43286_, _42806_, _37731_);
  and (_43287_, _43286_, _43222_);
  nor (_43288_, _43287_, _37885_);
  and (_43289_, _36763_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_43290_, _43289_, _37015_);
  and (_43291_, _43233_, _42634_);
  nor (_43292_, _43291_, _43290_);
  not (_43294_, _43292_);
  nor (_43295_, _43294_, _43288_);
  and (_43296_, _43295_, _43235_);
  and (_43298_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43299_, _43298_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_43300_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43302_, _43300_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_43303_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43304_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_43306_, _43304_, _43303_);
  and (_43307_, _43306_, _43302_);
  and (_43308_, _43307_, _43299_);
  and (_43310_, _43308_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43311_, _43310_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43312_, _43311_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_43314_, _43312_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43315_, _43314_, _38667_);
  or (_43316_, _43314_, _38667_);
  and (_43318_, _43316_, _43315_);
  and (_43319_, _43318_, _43296_);
  nor (_43321_, _43281_, _43235_);
  and (_43322_, _43295_, _43321_);
  not (_43323_, _36818_);
  and (_43324_, _43183_, _43323_);
  and (_43325_, _43324_, _43223_);
  and (_43327_, _43325_, _43286_);
  nor (_43328_, _43327_, _37885_);
  and (_43329_, _36807_, _42634_);
  and (_43331_, _43329_, _37004_);
  nor (_43332_, _43331_, _43328_);
  and (_43333_, _43332_, _43322_);
  and (_43335_, _43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43336_, _43291_, _40406_);
  or (_43337_, _43336_, _43335_);
  or (_43339_, _43337_, _43319_);
  nor (_43340_, _43339_, _43284_);
  nand (_43341_, _43340_, _43276_);
  or (_43343_, _43341_, _43280_);
  not (_43344_, _43331_);
  and (_43345_, _43295_, _43344_);
  and (_43347_, _43345_, _40405_);
  not (_43348_, _43345_);
  and (_43349_, _43348_, _43032_);
  nor (_43351_, _43349_, _43347_);
  and (_43352_, _43351_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_43354_, _43351_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_43355_, _43345_, _40624_);
  not (_43356_, _43151_);
  nor (_43357_, _43345_, _43356_);
  nor (_43358_, _43357_, _43355_);
  and (_43359_, _43358_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_43360_, _43358_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_43362_, _43360_, _43359_);
  and (_43363_, _43345_, _40442_);
  not (_43364_, _43134_);
  nor (_43366_, _43345_, _43364_);
  nor (_43367_, _43366_, _43363_);
  and (_43368_, _43367_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_43370_, _43367_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_43371_, _43345_, _40663_);
  not (_43372_, _43117_);
  nor (_43374_, _43345_, _43372_);
  nor (_43375_, _43374_, _43371_);
  nand (_43388_, _43375_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43393_, _43345_, _40530_);
  not (_43394_, _43100_);
  nor (_43408_, _43345_, _43394_);
  nor (_43413_, _43408_, _43393_);
  and (_43414_, _43413_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_43426_, _43413_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_43433_, _43345_, _40485_);
  not (_43434_, _43083_);
  nor (_43445_, _43345_, _43434_);
  nor (_43446_, _43445_, _43433_);
  and (_43454_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43462_, _43345_, _40736_);
  not (_43471_, _43066_);
  nor (_43472_, _43345_, _43471_);
  nor (_43481_, _43472_, _43462_);
  and (_43489_, _43481_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_43490_, _43345_, _40568_);
  not (_43501_, _43049_);
  nor (_43507_, _43345_, _43501_);
  nor (_43508_, _43507_, _43490_);
  and (_43520_, _43508_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_43526_, _43481_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_43527_, _43526_, _43489_);
  and (_43540_, _43527_, _43520_);
  nor (_43545_, _43540_, _43489_);
  not (_43546_, _43545_);
  nor (_43560_, _43446_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_43565_, _43560_, _43454_);
  and (_43566_, _43565_, _43546_);
  nor (_43578_, _43566_, _43454_);
  nor (_43585_, _43578_, _43426_);
  or (_43586_, _43585_, _43414_);
  or (_43597_, _43375_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43598_, _43597_, _43388_);
  nand (_43606_, _43598_, _43586_);
  and (_43614_, _43606_, _43388_);
  nor (_43616_, _43614_, _43370_);
  or (_43617_, _43616_, _43368_);
  and (_43618_, _43617_, _43362_);
  nor (_43620_, _43618_, _43359_);
  nor (_43621_, _43620_, _43354_);
  or (_43622_, _43621_, _43352_);
  and (_43624_, _43622_, _43299_);
  and (_43625_, _43624_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43626_, _43625_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43628_, _43626_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_43629_, _43628_, _43351_);
  not (_43630_, _43351_);
  nor (_43632_, _43622_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43633_, _43632_, _38645_);
  and (_43634_, _43633_, _38650_);
  and (_43636_, _43634_, _38635_);
  nor (_43637_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43638_, _43637_, _43636_);
  nor (_43640_, _43638_, _43630_);
  nor (_43641_, _43640_, _43629_);
  or (_43643_, _43351_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43644_, _43351_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_43645_, _43644_, _43643_);
  and (_43646_, _43645_, _43641_);
  or (_43648_, _43646_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_43649_, _43646_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_43650_, _43649_, _43648_);
  nor (_43652_, _43348_, _43321_);
  nor (_43653_, _43332_, _43652_);
  and (_43654_, _43653_, _43650_);
  or (_43656_, _43654_, _43343_);
  not (_43657_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_43660_, _43658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_43661_, _43660_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_43662_, _43661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_43664_, _43662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_43665_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_43666_, _43665_, _43664_);
  and (_43668_, _43666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_43669_, _43668_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_43670_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_43672_, _34402_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43673_, _43672_, _40389_);
  nor (_43675_, _43673_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_43676_, _43675_);
  and (_43677_, _43676_, _43670_);
  and (_43678_, _43677_, _43669_);
  nand (_43679_, _43678_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_43680_, _43679_, _43657_);
  or (_43681_, _43679_, _43657_);
  and (_43683_, _43681_, _43680_);
  or (_43684_, _43683_, _43276_);
  and (_43685_, _43684_, _41894_);
  and (_38970_, _43685_, _43656_);
  and (_43687_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _41894_);
  and (_43688_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_43690_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_43691_, _34358_, _43690_);
  not (_43692_, _43691_);
  not (_43694_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_43695_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_43696_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_43698_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_43699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_43700_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_43702_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_43703_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43704_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_43706_, _43704_, _43702_);
  and (_43707_, _43706_, _43703_);
  nor (_43709_, _43707_, _43702_);
  nor (_43710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43711_, _43710_, _43700_);
  not (_43712_, _43711_);
  nor (_43714_, _43712_, _43709_);
  nor (_43715_, _43714_, _43700_);
  not (_43716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_43718_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_43719_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_43720_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_43722_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_43723_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43724_, _43723_, _43722_);
  and (_43726_, _43724_, _43720_);
  and (_43727_, _43726_, _43719_);
  and (_43728_, _43727_, _43718_);
  and (_43730_, _43728_, _43716_);
  and (_43731_, _43730_, _43715_);
  and (_43732_, _43731_, _43699_);
  and (_43734_, _43732_, _43698_);
  and (_43735_, _43734_, _43696_);
  and (_43736_, _43735_, _43695_);
  and (_43738_, _43736_, _43694_);
  nor (_43739_, _43738_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43741_, _43738_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_43742_, _43741_, _43739_);
  nor (_43743_, _43736_, _43694_);
  nor (_43744_, _43743_, _43738_);
  not (_43746_, _43744_);
  nor (_43747_, _43735_, _43695_);
  nor (_43748_, _43747_, _43736_);
  not (_43750_, _43748_);
  nor (_43751_, _43734_, _43696_);
  nor (_43752_, _43751_, _43735_);
  not (_43754_, _43752_);
  nor (_43755_, _43732_, _43698_);
  nor (_43756_, _43755_, _43734_);
  not (_43758_, _43756_);
  nor (_43759_, _43731_, _43699_);
  nor (_43760_, _43759_, _43732_);
  not (_43762_, _43760_);
  and (_43763_, _43728_, _43715_);
  nor (_43764_, _43763_, _43716_);
  nor (_43766_, _43764_, _43731_);
  not (_43767_, _43766_);
  and (_43768_, _43715_, _43726_);
  nor (_43770_, _43768_, _43719_);
  and (_43771_, _43727_, _43715_);
  nor (_43773_, _43771_, _43770_);
  not (_43774_, _43773_);
  and (_43775_, _43715_, _43724_);
  nor (_43776_, _43775_, _43720_);
  nor (_43778_, _43776_, _43768_);
  not (_43779_, _43778_);
  and (_43780_, _43715_, _43723_);
  nor (_43782_, _43780_, _43722_);
  nor (_43783_, _43782_, _43775_);
  not (_43784_, _43783_);
  not (_43786_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43787_, _43715_, _43786_);
  nor (_43788_, _43715_, _43786_);
  nor (_43790_, _43788_, _43787_);
  not (_43791_, _43790_);
  or (_43792_, _42495_, _42485_);
  nand (_43794_, _43792_, _42511_);
  and (_43795_, _42520_, _42508_);
  nor (_43796_, _43795_, _42534_);
  and (_43798_, _42527_, _42479_);
  nor (_43799_, _43798_, _42503_);
  nor (_43800_, _43799_, _43796_);
  and (_43802_, _42502_, _42469_);
  and (_43803_, _43802_, _42485_);
  nor (_43805_, _43803_, _43800_);
  and (_43806_, _43805_, _43794_);
  not (_43807_, _42531_);
  nor (_43808_, _42538_, _42472_);
  nor (_43809_, _43808_, _43807_);
  and (_43811_, _42499_, _42469_);
  or (_43812_, _43802_, _43811_);
  and (_43813_, _43812_, _42534_);
  nor (_43815_, _43813_, _43809_);
  and (_43816_, _43815_, _43806_);
  not (_43817_, _43811_);
  and (_43819_, _43808_, _43817_);
  nor (_43820_, _43819_, _36281_);
  and (_43821_, _42508_, _42538_);
  and (_43823_, _42531_, _42500_);
  or (_43824_, _43823_, _43821_);
  and (_43825_, _43802_, _42476_);
  and (_43827_, _42487_, _42476_);
  or (_43828_, _43827_, _43825_);
  or (_43829_, _43828_, _43824_);
  and (_43831_, _42539_, _42520_);
  and (_43832_, _42492_, _42471_);
  and (_43833_, _43832_, _42531_);
  nor (_43835_, _43833_, _43831_);
  nand (_43836_, _43835_, _42546_);
  or (_43838_, _43836_, _43829_);
  nor (_43839_, _43838_, _43820_);
  and (_43840_, _42508_, _42487_);
  not (_43841_, _43840_);
  nor (_43843_, _42532_, _42530_);
  and (_43844_, _43843_, _43841_);
  not (_43845_, _42476_);
  and (_43847_, _42492_, _34991_);
  nor (_43848_, _43811_, _43847_);
  nor (_43849_, _43848_, _43845_);
  and (_43851_, _42502_, _42479_);
  not (_43852_, _43851_);
  nor (_43853_, _42534_, _42485_);
  nor (_43855_, _43853_, _43852_);
  nor (_43856_, _43855_, _43849_);
  and (_43857_, _43856_, _43844_);
  and (_43859_, _42479_, _42491_);
  and (_43860_, _42543_, _43859_);
  not (_43861_, _43860_);
  and (_43863_, _42518_, _42508_);
  and (_43864_, _42534_, _42472_);
  nor (_43865_, _43864_, _43863_);
  and (_43867_, _43865_, _43861_);
  and (_43868_, _42470_, _36039_);
  and (_43870_, _43868_, _42469_);
  and (_43871_, _43870_, _42484_);
  and (_43872_, _42533_, _42509_);
  nor (_43873_, _43872_, _43871_);
  and (_43875_, _43873_, _43867_);
  and (_43876_, _43875_, _43857_);
  and (_43877_, _43876_, _43839_);
  nor (_43879_, _42504_, _42477_);
  nor (_43880_, _42524_, _42481_);
  and (_43881_, _43880_, _43879_);
  not (_43883_, _42534_);
  nor (_43884_, _43832_, _42487_);
  nor (_43885_, _43884_, _43883_);
  and (_43887_, _42531_, _42533_);
  nor (_43888_, _43887_, _43885_);
  and (_43889_, _42531_, _42487_);
  and (_43891_, _42539_, _43851_);
  nor (_43892_, _43891_, _43889_);
  nand (_43893_, _42550_, _42531_);
  and (_43895_, _43893_, _43892_);
  and (_43896_, _43895_, _43888_);
  nor (_43897_, _42520_, _42496_);
  nor (_43899_, _43897_, _43807_);
  nor (_43900_, _43899_, _42551_);
  and (_43902_, _43900_, _43896_);
  and (_43903_, _43902_, _43881_);
  and (_43904_, _43903_, _43877_);
  and (_43905_, _43904_, _43816_);
  nor (_43907_, _43706_, _43703_);
  nor (_43908_, _43907_, _43707_);
  not (_43909_, _43908_);
  nor (_43911_, _43909_, _43905_);
  not (_43912_, _43911_);
  nand (_43913_, _43892_, _43844_);
  not (_43915_, _42551_);
  nand (_43916_, _43915_, _42546_);
  or (_43917_, _43916_, _43809_);
  or (_43919_, _43831_, _42519_);
  and (_43920_, _42539_, _42511_);
  or (_43921_, _43825_, _43920_);
  or (_43923_, _43921_, _43919_);
  or (_43924_, _43923_, _43917_);
  or (_43925_, _43924_, _43913_);
  nor (_43927_, _43925_, _43905_);
  not (_43928_, _43927_);
  nor (_43929_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43931_, _43929_, _43703_);
  and (_43932_, _43931_, _43928_);
  and (_43933_, _43909_, _43905_);
  nor (_43934_, _43933_, _43911_);
  nand (_43935_, _43934_, _43932_);
  and (_43936_, _43935_, _43912_);
  not (_43937_, _43936_);
  and (_43938_, _43712_, _43709_);
  nor (_43939_, _43938_, _43714_);
  and (_43940_, _43939_, _43937_);
  and (_43941_, _43940_, _43791_);
  not (_43942_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_43943_, _43787_, _43942_);
  or (_43944_, _43943_, _43780_);
  and (_43945_, _43944_, _43941_);
  and (_43946_, _43945_, _43784_);
  and (_43947_, _43946_, _43779_);
  and (_43948_, _43947_, _43774_);
  nor (_43949_, _43771_, _43718_);
  or (_43950_, _43949_, _43763_);
  and (_43951_, _43950_, _43948_);
  and (_43952_, _43951_, _43767_);
  and (_43953_, _43952_, _43762_);
  and (_43954_, _43953_, _43758_);
  and (_43955_, _43954_, _43754_);
  and (_43956_, _43955_, _43750_);
  and (_43957_, _43956_, _43746_);
  or (_43958_, _43957_, _43742_);
  nand (_43959_, _43957_, _43742_);
  and (_43960_, _43959_, _43958_);
  or (_43961_, _43960_, _43692_);
  or (_43962_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_43963_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_43964_, _43963_, _43962_);
  and (_43965_, _43964_, _43961_);
  or (_38971_, _43965_, _43688_);
  nor (_43966_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_38972_, _43966_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_38973_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _41894_);
  nor (_43967_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_43968_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_43969_, _43968_, _43967_);
  nor (_43970_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_43971_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_43972_, _43971_, _43970_);
  and (_43973_, _43972_, _43969_);
  nor (_43974_, _43973_, rst);
  and (_43975_, \oc8051_top_1.oc8051_rom1.ea_int , _34325_);
  nand (_43976_, _43975_, _34358_);
  and (_43977_, _43976_, _38973_);
  or (_38975_, _43977_, _43974_);
  and (_43978_, _43973_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_43979_, _43978_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_38976_, _43979_, _41894_);
  nor (_43980_, _43675_, _40389_);
  or (_43981_, _43905_, _34554_);
  nor (_43982_, _43927_, _34489_);
  nand (_43983_, _43905_, _34554_);
  and (_43984_, _43983_, _43981_);
  nand (_43985_, _43984_, _43982_);
  and (_43986_, _43985_, _43981_);
  nor (_43987_, _43986_, _40389_);
  and (_43988_, _43987_, _34391_);
  nor (_43989_, _43987_, _34391_);
  nor (_43990_, _43989_, _43988_);
  nor (_43991_, _43990_, _43980_);
  and (_43992_, _34565_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_43993_, _43992_, _43980_);
  and (_43994_, _43993_, _43925_);
  or (_43995_, _43994_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_43996_, _43995_, _43991_);
  and (_38977_, _43996_, _41894_);
  not (_43997_, _34684_);
  and (_43998_, _43997_, _35199_);
  not (_43999_, _36468_);
  nor (_44000_, _43999_, _35962_);
  and (_44001_, _44000_, _43998_);
  and (_44002_, _34369_, _41894_);
  and (_44003_, _44002_, _35444_);
  and (_44004_, _44003_, _34947_);
  nor (_44005_, _36237_, _35720_);
  and (_44006_, _44005_, _44004_);
  and (_38980_, _44006_, _44001_);
  nor (_44007_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_44008_, _44007_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_44009_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_38983_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _41894_);
  and (_44010_, _38983_, _44009_);
  or (_38982_, _44010_, _44008_);
  not (_44011_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_44012_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44013_, _44012_, _44011_);
  and (_44014_, _44012_, _44011_);
  nor (_44015_, _44014_, _44013_);
  not (_44016_, _44015_);
  and (_44017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_44018_, _44017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44019_, _44017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44020_, _44019_, _44018_);
  or (_44021_, _44020_, _44012_);
  and (_44022_, _44021_, _44016_);
  nor (_44023_, _44013_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_44024_, _44013_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_44025_, _44024_, _44023_);
  or (_44026_, _44018_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_38985_, _44026_, _41894_);
  and (_44027_, _38985_, _44025_);
  and (_38984_, _44027_, _44022_);
  not (_44028_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_44029_, _43675_, _44028_);
  and (_44030_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_44031_, _44029_);
  and (_44032_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_44033_, _44032_, _44030_);
  and (_38986_, _44033_, _41894_);
  and (_44034_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_44035_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_44036_, _44035_, _44034_);
  and (_38987_, _44036_, _41894_);
  and (_44037_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_44038_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_44039_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _44038_);
  and (_44040_, _44039_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_44041_, _44040_, _44037_);
  and (_38989_, _44041_, _41894_);
  and (_44042_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_44043_, _44042_, _44039_);
  and (_38990_, _44043_, _41894_);
  or (_44044_, _44038_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_38991_, _44044_, _41894_);
  not (_44045_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_44046_, _44045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_44047_, _44046_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_44048_, _44038_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_44049_, _44048_, _41894_);
  and (_38992_, _44049_, _44047_);
  or (_44050_, _44038_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_38993_, _44050_, _41894_);
  nor (_44051_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_44052_, _44051_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_44053_, _44052_, _41894_);
  and (_44054_, _38983_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_38994_, _44054_, _44053_);
  and (_44055_, _44028_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_44056_, _44055_, _44052_);
  and (_38995_, _44056_, _41894_);
  nand (_44057_, _44052_, _38678_);
  or (_44058_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_44059_, _44058_, _41894_);
  and (_38996_, _44059_, _44057_);
  nand (_44060_, _36960_, _41894_);
  nor (_38997_, _44060_, _38389_);
  or (_44061_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_44062_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_44063_, _43152_, _44062_);
  and (_44064_, _44063_, _41894_);
  and (_39034_, _44064_, _44061_);
  or (_44065_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_44066_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_44067_, _43152_, _44066_);
  and (_44068_, _44067_, _41894_);
  and (_39035_, _44068_, _44065_);
  or (_44069_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_44070_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_44071_, _43152_, _44070_);
  and (_44072_, _44071_, _41894_);
  and (_39036_, _44072_, _44069_);
  or (_44073_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_44074_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_44075_, _43152_, _44074_);
  and (_44076_, _44075_, _41894_);
  and (_39038_, _44076_, _44073_);
  or (_44077_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_44078_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_44079_, _43152_, _44078_);
  and (_44080_, _44079_, _41894_);
  and (_39039_, _44080_, _44077_);
  or (_44081_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_44082_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_44083_, _43152_, _44082_);
  and (_44084_, _44083_, _41894_);
  and (_39040_, _44084_, _44081_);
  or (_44085_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_44086_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_44087_, _43152_, _44086_);
  and (_44088_, _44087_, _41894_);
  and (_39041_, _44088_, _44085_);
  or (_44089_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_44090_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_44091_, _43152_, _44090_);
  and (_44092_, _44091_, _41894_);
  and (_39042_, _44092_, _44089_);
  or (_44093_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_44094_, _43152_, _38639_);
  and (_44095_, _44094_, _41894_);
  and (_39043_, _44095_, _44093_);
  or (_44096_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_44097_, _43152_, _38645_);
  and (_44098_, _44097_, _41894_);
  and (_39044_, _44098_, _44096_);
  or (_44099_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_44100_, _43152_, _38650_);
  and (_44101_, _44100_, _41894_);
  and (_39045_, _44101_, _44099_);
  or (_44102_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_44103_, _43152_, _38635_);
  and (_44104_, _44103_, _41894_);
  and (_39046_, _44104_, _44102_);
  or (_44105_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_44106_, _43152_, _38656_);
  and (_44107_, _44106_, _41894_);
  and (_39047_, _44107_, _44105_);
  or (_44108_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_44109_, _43152_, _38631_);
  and (_44110_, _44109_, _41894_);
  and (_39049_, _44110_, _44108_);
  or (_44111_, _43152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_44112_, _43152_, _38662_);
  and (_44113_, _44112_, _41894_);
  and (_39050_, _44113_, _44111_);
  or (_44114_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_44115_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _41894_);
  or (_44116_, _44115_, _00000_);
  and (_39054_, _44116_, _44114_);
  or (_44117_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_44118_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _41894_);
  or (_44119_, _44118_, _00000_);
  and (_39055_, _44119_, _44117_);
  or (_44120_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_44121_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _41894_);
  or (_44122_, _44121_, _00000_);
  and (_39056_, _44122_, _44120_);
  or (_44123_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_44124_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _41894_);
  or (_44125_, _44124_, _00000_);
  and (_39057_, _44125_, _44123_);
  or (_44126_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_44127_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _41894_);
  or (_44128_, _44127_, _00000_);
  and (_39058_, _44128_, _44126_);
  or (_44129_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_44130_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _41894_);
  or (_44131_, _44130_, _00000_);
  and (_39059_, _44131_, _44129_);
  or (_44132_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_44133_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _41894_);
  or (_44134_, _44133_, _00000_);
  and (_39060_, _44134_, _44132_);
  or (_44135_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_44136_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _41894_);
  or (_44137_, _44136_, _00000_);
  and (_39061_, _44137_, _44135_);
  or (_44138_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_44139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _41894_);
  or (_44140_, _44139_, _00000_);
  and (_39063_, _44140_, _44138_);
  or (_44141_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_44142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _41894_);
  or (_44143_, _44142_, _00000_);
  and (_39064_, _44143_, _44141_);
  or (_44144_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_44145_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _41894_);
  or (_44146_, _44145_, _00000_);
  and (_39065_, _44146_, _44144_);
  or (_44147_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_44148_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _41894_);
  or (_44149_, _44148_, _00000_);
  and (_39066_, _44149_, _44147_);
  or (_44150_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_44151_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _41894_);
  or (_44152_, _44151_, _00000_);
  and (_39067_, _44152_, _44150_);
  or (_00006_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_00007_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _41894_);
  or (_00008_, _00007_, _00000_);
  and (_39068_, _00008_, _00006_);
  or (_00009_, _43156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_00010_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _41894_);
  or (_00011_, _00010_, _00000_);
  and (_39069_, _00011_, _00009_);
  nor (_39245_, _35808_, rst);
  nor (_39246_, _36083_, rst);
  nor (_39247_, _36566_, rst);
  nor (_39248_, _40365_, rst);
  and (_00012_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00013_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_00014_, _00013_, _00012_);
  and (_39249_, _00014_, _41894_);
  and (_00015_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00016_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00017_, _00016_, _44029_);
  or (_00018_, _00017_, _00015_);
  and (_39250_, _00018_, _41894_);
  and (_00019_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00020_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_00021_, _00020_, _00019_);
  and (_39252_, _00021_, _41894_);
  and (_00022_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00023_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_00024_, _00023_, _00022_);
  and (_39253_, _00024_, _41894_);
  and (_00025_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00026_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_00027_, _00026_, _00025_);
  and (_39254_, _00027_, _41894_);
  and (_00028_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00029_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_00030_, _00029_, _44029_);
  or (_00031_, _00030_, _00028_);
  and (_39255_, _00031_, _41894_);
  and (_00032_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00033_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_00034_, _00033_, _00032_);
  and (_39256_, _00034_, _41894_);
  and (_00035_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00036_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_00037_, _00036_, _00035_);
  and (_39257_, _00037_, _41894_);
  and (_00038_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_00039_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_00040_, _00039_, _00038_);
  and (_39258_, _00040_, _41894_);
  and (_00041_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_00042_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_00043_, _00042_, _00041_);
  and (_39259_, _00043_, _41894_);
  and (_00044_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_00045_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_00046_, _00045_, _00044_);
  and (_39260_, _00046_, _41894_);
  and (_00047_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_00048_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_00049_, _00048_, _00047_);
  and (_39261_, _00049_, _41894_);
  and (_00050_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_00051_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_00052_, _00051_, _00050_);
  and (_39263_, _00052_, _41894_);
  and (_00053_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_00054_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_00055_, _00054_, _00053_);
  and (_39264_, _00055_, _41894_);
  and (_00056_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_00057_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_00058_, _00057_, _00056_);
  and (_39265_, _00058_, _41894_);
  and (_00059_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_00060_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_00061_, _00060_, _00059_);
  and (_39266_, _00061_, _41894_);
  and (_00062_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_00063_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_00064_, _00063_, _00062_);
  and (_39267_, _00064_, _41894_);
  and (_00065_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_00066_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_00067_, _00066_, _00065_);
  and (_39268_, _00067_, _41894_);
  and (_00068_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_00069_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_00070_, _00069_, _00068_);
  and (_39269_, _00070_, _41894_);
  and (_00071_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_00072_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_00073_, _00072_, _00071_);
  and (_39270_, _00073_, _41894_);
  and (_00074_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_00075_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_00076_, _00075_, _00074_);
  and (_39271_, _00076_, _41894_);
  and (_00077_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_00078_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_00079_, _00078_, _00077_);
  and (_39272_, _00079_, _41894_);
  and (_00080_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_00081_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_00082_, _00081_, _00080_);
  and (_39274_, _00082_, _41894_);
  and (_00083_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_00084_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_00085_, _00084_, _00083_);
  and (_39275_, _00085_, _41894_);
  and (_00086_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_00087_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_00088_, _00087_, _00086_);
  and (_39276_, _00088_, _41894_);
  and (_00089_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_00090_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_00091_, _00090_, _00089_);
  and (_39277_, _00091_, _41894_);
  and (_00092_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_00093_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_00094_, _00093_, _00092_);
  and (_39278_, _00094_, _41894_);
  and (_00095_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_00096_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_00097_, _00096_, _00095_);
  and (_39279_, _00097_, _41894_);
  and (_00098_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_00099_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_00100_, _00099_, _00098_);
  and (_39280_, _00100_, _41894_);
  and (_00101_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_00102_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_00103_, _00102_, _00101_);
  and (_39281_, _00103_, _41894_);
  and (_00104_, _44029_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_00105_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_00106_, _00105_, _00104_);
  and (_39282_, _00106_, _41894_);
  nor (_39284_, _40582_, rst);
  nor (_39285_, _40764_, rst);
  nor (_39286_, _40502_, rst);
  nor (_39287_, _40546_, rst);
  and (_39288_, _40675_, _41894_);
  nor (_39290_, _40463_, rst);
  nor (_39291_, _40608_, rst);
  and (_39307_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _41894_);
  and (_39308_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _41894_);
  and (_39309_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _41894_);
  and (_39311_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _41894_);
  and (_39312_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _41894_);
  and (_39313_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _41894_);
  and (_39314_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _41894_);
  nor (_00107_, _43333_, _43281_);
  nor (_00108_, _00107_, _29679_);
  and (_00109_, _43290_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00110_, _43296_, _40569_);
  and (_00111_, _43291_, _43501_);
  or (_00112_, _00111_, _00110_);
  or (_00113_, _00112_, _00109_);
  nor (_00114_, _43508_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00115_, _00114_, _43520_);
  and (_00116_, _00115_, _43653_);
  nor (_00117_, _00116_, _00113_);
  nand (_00118_, _00117_, _43276_);
  or (_00119_, _00118_, _00108_);
  or (_00120_, _43276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00121_, _00120_, _41894_);
  and (_39315_, _00121_, _00119_);
  nor (_00122_, _00107_, _30358_);
  and (_00123_, _43296_, _40737_);
  and (_00124_, _43291_, _43471_);
  and (_00125_, _37929_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00126_, _00125_, _00124_);
  or (_00127_, _00126_, _00123_);
  or (_00128_, _00127_, _00122_);
  nor (_00129_, _43527_, _43520_);
  nor (_00130_, _00129_, _43540_);
  nand (_00131_, _00130_, _43653_);
  nand (_00132_, _00131_, _43276_);
  or (_00133_, _00132_, _00128_);
  or (_00134_, _43276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00135_, _00134_, _41894_);
  and (_39316_, _00135_, _00133_);
  nor (_00136_, _00107_, _31069_);
  and (_00137_, _43290_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_00138_, _43296_, _40486_);
  and (_00139_, _43291_, _43434_);
  or (_00140_, _00139_, _00138_);
  or (_00141_, _00140_, _00137_);
  or (_00142_, _43565_, _43546_);
  not (_00143_, _43653_);
  nor (_00144_, _00143_, _43566_);
  and (_00145_, _00144_, _00142_);
  nor (_00146_, _00145_, _00141_);
  nand (_00147_, _00146_, _43276_);
  or (_00148_, _00147_, _00136_);
  not (_00149_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00150_, _43675_, _00149_);
  and (_00151_, _43675_, _00149_);
  nor (_00152_, _00151_, _00150_);
  or (_00153_, _00152_, _43276_);
  and (_00154_, _00153_, _41894_);
  and (_39317_, _00154_, _00148_);
  nor (_00155_, _00107_, _31822_);
  and (_00156_, _43290_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_00157_, _43296_, _40531_);
  and (_00158_, _43291_, _43394_);
  or (_00159_, _00158_, _00157_);
  or (_00160_, _00159_, _00156_);
  or (_00161_, _00160_, _00155_);
  not (_00162_, _43578_);
  or (_00163_, _43426_, _43414_);
  nor (_00164_, _00163_, _00162_);
  and (_00165_, _00163_, _00162_);
  or (_00166_, _00165_, _00164_);
  nand (_00167_, _00166_, _43653_);
  nand (_00168_, _00167_, _43276_);
  or (_00169_, _00168_, _00161_);
  and (_00170_, _00150_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00171_, _00150_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00172_, _00171_, _00170_);
  or (_00173_, _00172_, _43276_);
  and (_00174_, _00173_, _41894_);
  and (_39318_, _00174_, _00169_);
  nor (_00175_, _00107_, _32585_);
  and (_00176_, _43296_, _40664_);
  and (_00177_, _43291_, _43372_);
  or (_00178_, _00177_, _00176_);
  or (_00179_, _43598_, _43586_);
  and (_00180_, _43653_, _43606_);
  and (_00181_, _00180_, _00179_);
  or (_00182_, _00181_, _00178_);
  or (_00183_, _00182_, _00175_);
  nand (_00184_, _43290_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nand (_00185_, _00184_, _43276_);
  or (_00186_, _00185_, _00183_);
  and (_00187_, _43660_, _43676_);
  nor (_00188_, _00170_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00189_, _00188_, _00187_);
  or (_00190_, _00189_, _43276_);
  and (_00191_, _00190_, _41894_);
  and (_39319_, _00191_, _00186_);
  nor (_00192_, _00107_, _33379_);
  and (_00193_, _43296_, _40443_);
  and (_00194_, _43291_, _43364_);
  and (_00195_, _37929_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00196_, _00195_, _00194_);
  or (_00197_, _00196_, _00193_);
  or (_00198_, _00197_, _00192_);
  or (_00199_, _43370_, _43368_);
  nand (_00200_, _00199_, _43614_);
  or (_00201_, _00199_, _43614_);
  and (_00202_, _00201_, _00200_);
  nand (_00203_, _00202_, _43653_);
  nand (_00204_, _00203_, _43276_);
  or (_00205_, _00204_, _00198_);
  and (_00206_, _43661_, _43676_);
  nor (_00207_, _00187_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00208_, _00207_, _00206_);
  or (_00209_, _00208_, _43276_);
  and (_00210_, _00209_, _41894_);
  and (_39320_, _00210_, _00205_);
  not (_00211_, _43276_);
  nor (_00212_, _43617_, _43362_);
  nor (_00213_, _00212_, _43618_);
  and (_00214_, _00213_, _43653_);
  nor (_00215_, _00107_, _34098_);
  and (_00216_, _43296_, _40625_);
  and (_00217_, _43291_, _43356_);
  and (_00218_, _37929_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00219_, _00218_, _00217_);
  or (_00220_, _00219_, _00216_);
  or (_00221_, _00220_, _00215_);
  or (_00222_, _00221_, _00214_);
  or (_00223_, _00222_, _00211_);
  and (_00224_, _00206_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00225_, _00206_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00226_, _00225_, _00224_);
  or (_00227_, _00226_, _43276_);
  and (_00228_, _00227_, _41894_);
  and (_39322_, _00228_, _00223_);
  or (_00229_, _43352_, _43354_);
  nor (_00230_, _00229_, _43620_);
  and (_00231_, _00229_, _43620_);
  or (_00232_, _00231_, _00230_);
  or (_00233_, _00232_, _00143_);
  or (_00234_, _00107_, _28496_);
  nand (_00235_, _43290_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nand (_00236_, _43296_, _40406_);
  not (_00237_, _43032_);
  nand (_00238_, _43291_, _00237_);
  and (_00239_, _00238_, _00236_);
  and (_00240_, _00239_, _00235_);
  and (_00241_, _00240_, _00234_);
  and (_00242_, _00241_, _00233_);
  nand (_00243_, _00242_, _43276_);
  and (_00244_, _00224_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00245_, _00224_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00246_, _00245_, _00244_);
  or (_00247_, _00246_, _43276_);
  and (_00248_, _00247_, _41894_);
  and (_39323_, _00248_, _00243_);
  and (_00249_, _43622_, _38639_);
  nor (_00250_, _43622_, _38639_);
  nor (_00251_, _00250_, _00249_);
  nor (_00252_, _00251_, _43351_);
  and (_00253_, _00251_, _43351_);
  or (_00254_, _00253_, _00252_);
  and (_00255_, _00254_, _43653_);
  not (_00256_, _43290_);
  nor (_00257_, _00256_, _29679_);
  nor (_00258_, _43283_, _38712_);
  and (_00259_, _43296_, _42491_);
  and (_00260_, _43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_00261_, _43291_, _40569_);
  or (_00262_, _00261_, _00260_);
  or (_00263_, _00262_, _00259_);
  or (_00264_, _00263_, _00258_);
  or (_00265_, _00264_, _00257_);
  or (_00266_, _00265_, _00255_);
  or (_00267_, _00266_, _00211_);
  and (_00268_, _00244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00269_, _00244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00270_, _00269_, _00268_);
  or (_00271_, _00270_, _43276_);
  and (_00272_, _00271_, _41894_);
  and (_39324_, _00272_, _00267_);
  nor (_00273_, _43283_, _38740_);
  and (_00274_, _43296_, _42478_);
  and (_00275_, _43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_00276_, _43291_, _40737_);
  or (_00277_, _00276_, _00275_);
  or (_00278_, _00277_, _00274_);
  or (_00279_, _00278_, _00273_);
  nor (_00280_, _00256_, _30358_);
  or (_00281_, _00280_, _00279_);
  and (_00282_, _43622_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00283_, _00282_, _43630_);
  and (_00284_, _43632_, _43351_);
  nor (_00285_, _00284_, _00283_);
  nor (_00286_, _00285_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00287_, _00285_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_00288_, _00287_, _00286_);
  and (_00289_, _00288_, _43653_);
  or (_00290_, _00289_, _00211_);
  or (_00291_, _00290_, _00281_);
  and (_00292_, _43666_, _43676_);
  nor (_00293_, _00268_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00294_, _00293_, _00292_);
  or (_00295_, _00294_, _43276_);
  and (_00296_, _00295_, _41894_);
  and (_39325_, _00296_, _00291_);
  nor (_00297_, _00256_, _31069_);
  nor (_00298_, _43283_, _38768_);
  and (_00299_, _43296_, _42468_);
  and (_00300_, _43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00301_, _43291_, _40486_);
  or (_00302_, _00301_, _00300_);
  or (_00303_, _00302_, _00299_);
  or (_00304_, _00303_, _00298_);
  and (_00305_, _43633_, _43351_);
  and (_00306_, _00283_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_00307_, _00306_, _00305_);
  nand (_00308_, _00307_, _38650_);
  or (_00309_, _00307_, _38650_);
  and (_00310_, _00309_, _00308_);
  and (_00311_, _00310_, _43653_);
  or (_00312_, _00311_, _00304_);
  or (_00313_, _00312_, _00297_);
  or (_00314_, _00313_, _00211_);
  and (_00315_, _00292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00316_, _00292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00317_, _00316_, _00315_);
  or (_00318_, _00317_, _43276_);
  and (_00319_, _00318_, _41894_);
  and (_39326_, _00319_, _00314_);
  and (_00320_, _43624_, _43630_);
  and (_00321_, _43634_, _43351_);
  nor (_00322_, _00321_, _00320_);
  nand (_00323_, _00322_, _38635_);
  or (_00324_, _00322_, _38635_);
  and (_00325_, _00324_, _00323_);
  and (_00326_, _00325_, _43653_);
  nor (_00327_, _43283_, _38796_);
  nor (_00328_, _43308_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00329_, _00328_, _43310_);
  and (_00330_, _00329_, _43296_);
  and (_00331_, _43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_00332_, _43291_, _40531_);
  or (_00333_, _00332_, _00331_);
  or (_00334_, _00333_, _00330_);
  or (_00335_, _00334_, _00327_);
  nor (_00336_, _00256_, _31822_);
  or (_00337_, _00336_, _00335_);
  or (_00338_, _00337_, _00326_);
  or (_00339_, _00338_, _00211_);
  and (_00340_, _00315_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00341_, _00315_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00342_, _00341_, _00340_);
  or (_00343_, _00342_, _43276_);
  and (_00344_, _00343_, _41894_);
  and (_39327_, _00344_, _00339_);
  and (_00345_, _43625_, _43630_);
  and (_00346_, _43636_, _43351_);
  nor (_00347_, _00346_, _00345_);
  or (_00348_, _00347_, _38656_);
  nand (_00349_, _00347_, _38656_);
  and (_00350_, _00349_, _43653_);
  and (_00351_, _00350_, _00348_);
  nor (_00352_, _43310_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00353_, _00352_, _43311_);
  and (_00354_, _00353_, _43296_);
  nor (_00355_, _00256_, _32585_);
  nor (_00356_, _43283_, _38824_);
  and (_00357_, _43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_00358_, _43291_, _40664_);
  or (_00359_, _00358_, _00357_);
  or (_00360_, _00359_, _00356_);
  or (_00361_, _00360_, _00355_);
  or (_00362_, _00361_, _00354_);
  or (_00363_, _00362_, _00351_);
  or (_00364_, _00363_, _00211_);
  and (_00365_, _00340_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00366_, _00340_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00367_, _00366_, _00365_);
  or (_00368_, _00367_, _43276_);
  and (_00369_, _00368_, _41894_);
  and (_39328_, _00369_, _00364_);
  nor (_00370_, _00256_, _33379_);
  nor (_00371_, _43283_, _38854_);
  and (_00372_, _43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_00373_, _43291_, _40443_);
  or (_00374_, _00373_, _00372_);
  or (_00375_, _00374_, _00371_);
  or (_00376_, _00375_, _00370_);
  and (_00377_, _43626_, _43630_);
  and (_00378_, _00346_, _38656_);
  nor (_00379_, _00378_, _00377_);
  nand (_00380_, _00379_, _38631_);
  or (_00381_, _00379_, _38631_);
  and (_00382_, _00381_, _00380_);
  and (_00383_, _00382_, _43653_);
  or (_00384_, _00383_, _00376_);
  nor (_00385_, _43311_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00386_, _00385_, _43312_);
  nand (_00387_, _00386_, _43296_);
  nand (_00388_, _00387_, _43276_);
  or (_00389_, _00388_, _00384_);
  or (_00390_, _00365_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_00391_, _00365_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_00392_, _00391_, _00390_);
  or (_00393_, _00392_, _43276_);
  and (_00394_, _00393_, _41894_);
  and (_39329_, _00394_, _00389_);
  or (_00395_, _43312_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00396_, _00395_, _43314_);
  nand (_00397_, _00396_, _43296_);
  or (_00398_, _00256_, _34098_);
  or (_00399_, _43283_, _38905_);
  nand (_00400_, _43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_00401_, _43291_, _40625_);
  and (_00402_, _00401_, _00400_);
  and (_00403_, _00402_, _00399_);
  and (_00404_, _00403_, _00398_);
  and (_00405_, _00404_, _00397_);
  and (_00406_, _43641_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_00407_, _43641_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_00408_, _00407_, _00406_);
  or (_00409_, _00408_, _00143_);
  and (_00410_, _00409_, _00405_);
  nand (_00411_, _00410_, _43276_);
  or (_00412_, _43678_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00413_, _00412_, _43679_);
  or (_00414_, _00413_, _43276_);
  and (_00415_, _00414_, _41894_);
  and (_39330_, _00415_, _00411_);
  and (_00416_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_00417_, _43931_, _43928_);
  nor (_00418_, _00417_, _43932_);
  or (_00419_, _00418_, _43692_);
  or (_00420_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00421_, _00420_, _43963_);
  and (_00422_, _00421_, _00419_);
  or (_39331_, _00422_, _00416_);
  or (_00423_, _43934_, _43932_);
  and (_00424_, _00423_, _43935_);
  or (_00425_, _00424_, _43692_);
  or (_00426_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00427_, _00426_, _43963_);
  and (_00428_, _00427_, _00425_);
  and (_00429_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39333_, _00429_, _00428_);
  and (_00430_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00431_, _43939_, _43937_);
  nor (_00432_, _00431_, _43940_);
  or (_00433_, _00432_, _43692_);
  or (_00434_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00435_, _00434_, _43963_);
  and (_00436_, _00435_, _00433_);
  or (_39334_, _00436_, _00430_);
  nor (_00437_, _43940_, _43791_);
  nor (_00438_, _00437_, _43941_);
  or (_00439_, _00438_, _43692_);
  or (_00440_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00441_, _00440_, _43963_);
  and (_00442_, _00441_, _00439_);
  and (_00443_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_39335_, _00443_, _00442_);
  and (_00444_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00445_, _43944_, _43941_);
  nor (_00446_, _00445_, _43945_);
  or (_00447_, _00446_, _43692_);
  or (_00448_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00449_, _00448_, _43963_);
  and (_00450_, _00449_, _00447_);
  or (_39336_, _00450_, _00444_);
  and (_00451_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00452_, _43945_, _43784_);
  nor (_00453_, _00452_, _43946_);
  or (_00454_, _00453_, _43692_);
  or (_00455_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_00456_, _00455_, _43963_);
  and (_00457_, _00456_, _00454_);
  or (_39337_, _00457_, _00451_);
  nor (_00458_, _43946_, _43779_);
  nor (_00459_, _00458_, _43947_);
  or (_00460_, _00459_, _43692_);
  or (_00461_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00462_, _00461_, _43963_);
  and (_00463_, _00462_, _00460_);
  and (_00464_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39338_, _00464_, _00463_);
  and (_00465_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00466_, _43947_, _43774_);
  nor (_00467_, _00466_, _43948_);
  or (_00468_, _00467_, _43692_);
  or (_00469_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_00470_, _00469_, _43963_);
  and (_00471_, _00470_, _00468_);
  or (_39339_, _00471_, _00465_);
  nor (_00472_, _43950_, _43948_);
  nor (_00473_, _00472_, _43951_);
  or (_00474_, _00473_, _43692_);
  or (_00475_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00476_, _00475_, _43963_);
  and (_00477_, _00476_, _00474_);
  and (_00478_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_39340_, _00478_, _00477_);
  nor (_00479_, _43951_, _43767_);
  nor (_00480_, _00479_, _43952_);
  or (_00481_, _00480_, _43692_);
  or (_00482_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00483_, _00482_, _43963_);
  and (_00484_, _00483_, _00481_);
  and (_00485_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39341_, _00485_, _00484_);
  nor (_00486_, _43952_, _43762_);
  nor (_00487_, _00486_, _43953_);
  or (_00488_, _00487_, _43692_);
  or (_00489_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00490_, _00489_, _43963_);
  and (_00491_, _00490_, _00488_);
  and (_00492_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_39342_, _00492_, _00491_);
  nor (_00493_, _43953_, _43758_);
  nor (_00494_, _00493_, _43954_);
  or (_00495_, _00494_, _43692_);
  or (_00496_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00497_, _00496_, _43963_);
  and (_00498_, _00497_, _00495_);
  and (_00499_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39343_, _00499_, _00498_);
  nor (_00500_, _43954_, _43754_);
  nor (_00501_, _00500_, _43955_);
  or (_00502_, _00501_, _43692_);
  or (_00503_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00504_, _00503_, _43963_);
  and (_00505_, _00504_, _00502_);
  and (_00506_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_39344_, _00506_, _00505_);
  nor (_00507_, _43955_, _43750_);
  nor (_00508_, _00507_, _43956_);
  or (_00509_, _00508_, _43692_);
  or (_00510_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00511_, _00510_, _43963_);
  and (_00512_, _00511_, _00509_);
  and (_00513_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_39345_, _00513_, _00512_);
  and (_00514_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_00515_, _43956_, _43746_);
  nor (_00516_, _00515_, _43957_);
  or (_00517_, _00516_, _43692_);
  or (_00518_, _43691_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00519_, _00518_, _43963_);
  and (_00520_, _00519_, _00517_);
  or (_39346_, _00520_, _00514_);
  and (_00521_, _43973_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_00522_, _00521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39347_, _00522_, _41894_);
  and (_00523_, _43973_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_00524_, _00523_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39348_, _00524_, _41894_);
  and (_00525_, _43973_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_00526_, _00525_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39349_, _00526_, _41894_);
  and (_00527_, _43973_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_00528_, _00527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39350_, _00528_, _41894_);
  and (_00529_, _43973_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_00530_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39351_, _00530_, _41894_);
  and (_00531_, _43973_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_00532_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39352_, _00532_, _41894_);
  and (_00533_, _43973_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_00534_, _00533_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39354_, _00534_, _41894_);
  nor (_00535_, _43927_, _40389_);
  nand (_00536_, _00535_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00537_, _00535_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00538_, _00537_, _43963_);
  and (_39355_, _00538_, _00536_);
  or (_00539_, _43984_, _43982_);
  and (_00540_, _00539_, _43985_);
  or (_00541_, _00540_, _40389_);
  or (_00542_, _34358_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00543_, _00542_, _43963_);
  and (_39356_, _00543_, _00541_);
  and (_00544_, _44007_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_00545_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_00546_, _00545_, _38983_);
  or (_39372_, _00546_, _00544_);
  and (_00547_, _44007_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00548_, _00016_, _38983_);
  or (_39373_, _00548_, _00547_);
  and (_00549_, _44007_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00550_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00551_, _00550_, _38983_);
  or (_39374_, _00551_, _00549_);
  and (_00552_, _44007_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00553_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_00554_, _00553_, _38983_);
  or (_39376_, _00554_, _00552_);
  and (_00555_, _44007_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00556_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_00557_, _00556_, _38983_);
  or (_39377_, _00557_, _00555_);
  and (_00558_, _44007_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00559_, _00029_, _38983_);
  or (_39378_, _00559_, _00558_);
  and (_00560_, _44007_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00561_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_00562_, _00561_, _38983_);
  or (_39379_, _00562_, _00560_);
  and (_39380_, _44015_, _41894_);
  nor (_39381_, _44025_, rst);
  and (_39382_, _44021_, _41894_);
  and (_00563_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00564_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00565_, _00564_, _00563_);
  and (_39383_, _00565_, _41894_);
  and (_00566_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00567_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00568_, _00567_, _00566_);
  and (_39384_, _00568_, _41894_);
  and (_00569_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00570_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00571_, _00570_, _00569_);
  and (_39385_, _00571_, _41894_);
  and (_00572_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00573_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00574_, _00573_, _00572_);
  and (_39387_, _00574_, _41894_);
  and (_00575_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00576_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00577_, _00576_, _00575_);
  and (_39388_, _00577_, _41894_);
  and (_00578_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00579_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00580_, _00579_, _00578_);
  and (_39389_, _00580_, _41894_);
  and (_00581_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00582_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00583_, _00582_, _00581_);
  and (_39390_, _00583_, _41894_);
  and (_00584_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00585_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00586_, _00585_, _00584_);
  and (_39391_, _00586_, _41894_);
  and (_00587_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00588_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00589_, _00588_, _00587_);
  and (_39392_, _00589_, _41894_);
  and (_00590_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00591_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00592_, _00591_, _00590_);
  and (_39393_, _00592_, _41894_);
  and (_00593_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00594_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00595_, _00594_, _00593_);
  and (_39394_, _00595_, _41894_);
  and (_00596_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00597_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00598_, _00597_, _00596_);
  and (_39395_, _00598_, _41894_);
  and (_00599_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00600_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00601_, _00600_, _00599_);
  and (_39396_, _00601_, _41894_);
  and (_00602_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00603_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00604_, _00603_, _00602_);
  and (_39398_, _00604_, _41894_);
  and (_00605_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00606_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00607_, _00606_, _00605_);
  and (_39399_, _00607_, _41894_);
  and (_00608_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00609_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00610_, _00609_, _00608_);
  and (_39400_, _00610_, _41894_);
  and (_00611_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00612_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00613_, _00612_, _00611_);
  and (_39401_, _00613_, _41894_);
  and (_00614_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00615_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00616_, _00615_, _00614_);
  and (_39402_, _00616_, _41894_);
  and (_00617_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00618_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00619_, _00618_, _00617_);
  and (_39403_, _00619_, _41894_);
  and (_00620_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00621_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00622_, _00621_, _00620_);
  and (_39404_, _00622_, _41894_);
  and (_00623_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00624_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00625_, _00624_, _00623_);
  and (_39405_, _00625_, _41894_);
  and (_00626_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00627_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00628_, _00627_, _00626_);
  and (_39406_, _00628_, _41894_);
  and (_00629_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00630_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00631_, _00630_, _00629_);
  and (_39407_, _00631_, _41894_);
  and (_00632_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00633_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00634_, _00633_, _00632_);
  and (_39409_, _00634_, _41894_);
  and (_00635_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00636_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00637_, _00636_, _00635_);
  and (_39410_, _00637_, _41894_);
  and (_00638_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00639_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00640_, _00639_, _00638_);
  and (_39411_, _00640_, _41894_);
  and (_00641_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00642_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00643_, _00642_, _00641_);
  and (_39412_, _00643_, _41894_);
  and (_00644_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00645_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00646_, _00645_, _00644_);
  and (_39413_, _00646_, _41894_);
  and (_00647_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00648_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00649_, _00648_, _00647_);
  and (_39414_, _00649_, _41894_);
  and (_00650_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00651_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00652_, _00651_, _00650_);
  and (_39415_, _00652_, _41894_);
  and (_00653_, _44029_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00654_, _44031_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00655_, _00654_, _00653_);
  and (_39416_, _00655_, _41894_);
  and (_00656_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00657_, _44039_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00658_, _00657_, _00656_);
  and (_39417_, _00658_, _41894_);
  and (_00659_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00660_, _44039_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00661_, _00660_, _00659_);
  and (_39418_, _00661_, _41894_);
  and (_00662_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00663_, _44039_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00664_, _00663_, _00662_);
  and (_39420_, _00664_, _41894_);
  and (_00665_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00666_, _44039_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00667_, _00666_, _00665_);
  and (_39421_, _00667_, _41894_);
  and (_00668_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00669_, _44039_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00670_, _00669_, _00668_);
  and (_39422_, _00670_, _41894_);
  and (_00671_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00672_, _44039_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00673_, _00672_, _00671_);
  and (_39423_, _00673_, _41894_);
  and (_00674_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00675_, _44039_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00676_, _00675_, _00674_);
  and (_39424_, _00676_, _41894_);
  and (_00677_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00678_, _40582_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00679_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00680_, _00679_, _44038_);
  and (_00681_, _00680_, _00678_);
  or (_00682_, _00681_, _00677_);
  and (_39425_, _00682_, _41894_);
  and (_00683_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00684_, _40764_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00685_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00686_, _00685_, _44038_);
  and (_00687_, _00686_, _00684_);
  or (_00688_, _00687_, _00683_);
  and (_39426_, _00688_, _41894_);
  and (_00689_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00690_, _40502_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00691_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00692_, _00691_, _44038_);
  and (_00693_, _00692_, _00690_);
  or (_00694_, _00693_, _00689_);
  and (_39427_, _00694_, _41894_);
  and (_00695_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00696_, _40546_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00697_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00698_, _00697_, _44038_);
  and (_00699_, _00698_, _00696_);
  or (_00700_, _00699_, _00695_);
  and (_39428_, _00700_, _41894_);
  and (_00701_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00702_, _40675_, _44045_);
  or (_00703_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00704_, _00703_, _44038_);
  and (_00705_, _00704_, _00702_);
  or (_00706_, _00705_, _00701_);
  and (_39429_, _00706_, _41894_);
  and (_00707_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00708_, _40463_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00709_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00710_, _00709_, _44038_);
  and (_00711_, _00710_, _00708_);
  or (_00712_, _00711_, _00707_);
  and (_39431_, _00712_, _41894_);
  and (_00713_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00714_, _40608_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00715_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00716_, _00715_, _44038_);
  and (_00717_, _00716_, _00714_);
  or (_00718_, _00717_, _00713_);
  and (_39432_, _00718_, _41894_);
  and (_00719_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00720_, _40383_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00721_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00722_, _00721_, _44038_);
  and (_00723_, _00722_, _00720_);
  or (_00724_, _00723_, _00719_);
  and (_39433_, _00724_, _41894_);
  and (_00725_, _44045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00726_, _00725_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00727_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _44038_);
  and (_00728_, _00727_, _41894_);
  and (_39434_, _00728_, _00726_);
  and (_00729_, _44045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00730_, _00729_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00731_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _44038_);
  and (_00732_, _00731_, _41894_);
  and (_39435_, _00732_, _00730_);
  and (_00733_, _44045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00734_, _00733_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00735_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _44038_);
  and (_00736_, _00735_, _41894_);
  and (_39436_, _00736_, _00734_);
  and (_00737_, _44045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00738_, _00737_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00739_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _44038_);
  and (_00740_, _00739_, _41894_);
  and (_39437_, _00740_, _00738_);
  and (_00741_, _44045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00742_, _00741_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00743_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _44038_);
  and (_00744_, _00743_, _41894_);
  and (_39438_, _00744_, _00742_);
  and (_00745_, _44045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_00746_, _00745_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00747_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _44038_);
  and (_00748_, _00747_, _41894_);
  and (_39439_, _00748_, _00746_);
  and (_00749_, _44045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_00750_, _00749_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00751_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _44038_);
  and (_00752_, _00751_, _41894_);
  and (_39440_, _00752_, _00750_);
  nand (_00753_, _44052_, _29679_);
  or (_00754_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00755_, _00754_, _41894_);
  and (_39442_, _00755_, _00753_);
  nand (_00756_, _44052_, _30358_);
  or (_00757_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00758_, _00757_, _41894_);
  and (_39443_, _00758_, _00756_);
  nand (_00759_, _44052_, _31069_);
  or (_00760_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00761_, _00760_, _41894_);
  and (_39444_, _00761_, _00759_);
  nand (_00762_, _44052_, _31822_);
  or (_00763_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00764_, _00763_, _41894_);
  and (_39445_, _00764_, _00762_);
  nand (_00765_, _44052_, _32585_);
  or (_00766_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00767_, _00766_, _41894_);
  and (_39446_, _00767_, _00765_);
  nand (_00768_, _44052_, _33379_);
  or (_00769_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00770_, _00769_, _41894_);
  and (_39447_, _00770_, _00768_);
  nand (_00771_, _44052_, _34098_);
  or (_00772_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00773_, _00772_, _41894_);
  and (_39448_, _00773_, _00771_);
  nand (_00774_, _44052_, _28496_);
  or (_00775_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00776_, _00775_, _41894_);
  and (_39449_, _00776_, _00774_);
  nand (_00777_, _44052_, _38712_);
  or (_00778_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00779_, _00778_, _41894_);
  and (_39450_, _00779_, _00777_);
  nand (_00780_, _44052_, _38740_);
  or (_00781_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00782_, _00781_, _41894_);
  and (_39451_, _00782_, _00780_);
  nand (_00783_, _44052_, _38768_);
  or (_00784_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00785_, _00784_, _41894_);
  and (_39453_, _00785_, _00783_);
  nand (_00786_, _44052_, _38796_);
  or (_00787_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00788_, _00787_, _41894_);
  and (_39454_, _00788_, _00786_);
  nand (_00789_, _44052_, _38824_);
  or (_00790_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00791_, _00790_, _41894_);
  and (_39455_, _00791_, _00789_);
  nand (_00792_, _44052_, _38854_);
  or (_00793_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00794_, _00793_, _41894_);
  and (_39456_, _00794_, _00792_);
  nand (_00795_, _44052_, _38905_);
  or (_00796_, _44052_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00797_, _00796_, _41894_);
  and (_39457_, _00797_, _00795_);
  nor (_39668_, _40425_, rst);
  and (_00798_, _39111_, _25395_);
  and (_00799_, _00798_, _40359_);
  nand (_00800_, _00799_, _38540_);
  or (_00801_, _00799_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_00802_, _00801_, _41894_);
  and (_39669_, _00802_, _00800_);
  and (_00803_, _38452_, _25395_);
  not (_00804_, _00803_);
  nor (_00805_, _00804_, _38540_);
  not (_00806_, _40359_);
  and (_00807_, _00804_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_00808_, _00807_, _00806_);
  or (_00809_, _00808_, _00805_);
  or (_00810_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_00811_, _00810_, _41894_);
  and (_39670_, _00811_, _00809_);
  not (_00812_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_00813_, _39959_, _24895_);
  and (_00814_, _00813_, _25395_);
  and (_00815_, _00814_, _40359_);
  nor (_00816_, _00815_, _00812_);
  and (_00817_, _00815_, _40355_);
  or (_00818_, _00817_, _00816_);
  and (_39672_, _00818_, _41894_);
  and (_00819_, _39959_, _30479_);
  and (_00820_, _00819_, _25395_);
  not (_00821_, _00820_);
  nor (_00822_, _00821_, _38540_);
  and (_00823_, _00821_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_00824_, _00823_, _00806_);
  or (_00825_, _00824_, _00822_);
  or (_00826_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_00827_, _00826_, _41894_);
  and (_39673_, _00827_, _00825_);
  nand (_00828_, _00799_, _38518_);
  or (_00829_, _00799_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_00830_, _00829_, _41894_);
  and (_39701_, _00830_, _00828_);
  nand (_00831_, _00799_, _38509_);
  or (_00832_, _00799_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_00833_, _00832_, _41894_);
  and (_39702_, _00833_, _00831_);
  nand (_00834_, _00799_, _38502_);
  or (_00835_, _00799_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_00836_, _00835_, _41894_);
  and (_39703_, _00836_, _00834_);
  nand (_00837_, _00799_, _38494_);
  or (_00838_, _00799_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_00840_, _00838_, _41894_);
  and (_39704_, _00840_, _00837_);
  nand (_00841_, _00799_, _38486_);
  or (_00842_, _00799_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_00843_, _00842_, _41894_);
  and (_39705_, _00843_, _00841_);
  nand (_00844_, _00799_, _38479_);
  or (_00845_, _00799_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_00846_, _00845_, _41894_);
  and (_39707_, _00846_, _00844_);
  nand (_00847_, _00799_, _38472_);
  or (_00848_, _00799_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_00849_, _00848_, _41894_);
  and (_39708_, _00849_, _00847_);
  nor (_00850_, _00804_, _38518_);
  and (_00851_, _00804_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_00852_, _00851_, _00806_);
  or (_00853_, _00852_, _00850_);
  or (_00854_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_00855_, _00854_, _41894_);
  and (_39709_, _00855_, _00853_);
  not (_00856_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_00857_, _00803_, _40359_);
  nor (_00858_, _00857_, _00856_);
  and (_00859_, _00857_, _38510_);
  or (_00860_, _00859_, _00858_);
  and (_39710_, _00860_, _41894_);
  nor (_00861_, _00804_, _38502_);
  and (_00862_, _00804_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_00863_, _00862_, _00806_);
  or (_00865_, _00863_, _00861_);
  or (_00866_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_00867_, _00866_, _41894_);
  and (_39711_, _00867_, _00865_);
  nor (_00868_, _00804_, _38494_);
  and (_00869_, _00804_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_00870_, _00869_, _00806_);
  or (_00871_, _00870_, _00868_);
  or (_00872_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_00873_, _00872_, _41894_);
  and (_39712_, _00873_, _00871_);
  nor (_00874_, _00804_, _38486_);
  and (_00875_, _00804_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_00876_, _00875_, _00806_);
  or (_00877_, _00876_, _00874_);
  or (_00878_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_00879_, _00878_, _41894_);
  and (_39713_, _00879_, _00877_);
  nor (_00880_, _00804_, _38479_);
  and (_00881_, _00804_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_00883_, _00881_, _00806_);
  or (_00884_, _00883_, _00880_);
  or (_00885_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_00886_, _00885_, _41894_);
  and (_39714_, _00886_, _00884_);
  nor (_00887_, _00804_, _38472_);
  and (_00888_, _00804_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_00889_, _00888_, _00806_);
  or (_00890_, _00889_, _00887_);
  or (_00891_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_00892_, _00891_, _41894_);
  and (_39715_, _00892_, _00890_);
  or (_00893_, _00814_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand (_00894_, _00814_, _38518_);
  and (_00895_, _00894_, _00893_);
  or (_00896_, _00895_, _00806_);
  or (_00897_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_00898_, _00897_, _41894_);
  and (_39716_, _00898_, _00896_);
  not (_00899_, _00814_);
  nor (_00900_, _00899_, _38509_);
  and (_00901_, _00899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_00902_, _00901_, _00806_);
  or (_00903_, _00902_, _00900_);
  or (_00904_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_00905_, _00904_, _41894_);
  and (_39718_, _00905_, _00903_);
  nor (_00906_, _00899_, _38502_);
  and (_00907_, _00899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_00908_, _00907_, _00806_);
  or (_00909_, _00908_, _00906_);
  or (_00910_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_00911_, _00910_, _41894_);
  and (_39719_, _00911_, _00909_);
  nor (_00912_, _00899_, _38494_);
  and (_00913_, _00899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_00914_, _00913_, _00806_);
  or (_00915_, _00914_, _00912_);
  or (_00916_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_00917_, _00916_, _41894_);
  and (_39720_, _00917_, _00915_);
  nor (_00918_, _00899_, _38486_);
  and (_00919_, _00899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_00920_, _00919_, _00806_);
  or (_00921_, _00920_, _00918_);
  or (_00922_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_00923_, _00922_, _41894_);
  and (_39721_, _00923_, _00921_);
  nor (_00924_, _00899_, _38479_);
  and (_00925_, _00899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_00926_, _00925_, _00806_);
  or (_00927_, _00926_, _00924_);
  or (_00928_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_00929_, _00928_, _41894_);
  and (_39722_, _00929_, _00927_);
  nor (_00930_, _00899_, _38472_);
  and (_00931_, _00899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_00932_, _00931_, _00806_);
  or (_00933_, _00932_, _00930_);
  or (_00934_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_00935_, _00934_, _41894_);
  and (_39723_, _00935_, _00933_);
  and (_00936_, _00821_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_00937_, _00821_, _38518_);
  or (_00938_, _00937_, _00806_);
  or (_00939_, _00938_, _00936_);
  or (_00940_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_00941_, _00940_, _41894_);
  and (_39724_, _00941_, _00939_);
  nor (_00942_, _00821_, _38509_);
  and (_00943_, _00821_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_00944_, _00943_, _00806_);
  or (_00945_, _00944_, _00942_);
  or (_00946_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_00947_, _00946_, _41894_);
  and (_39725_, _00947_, _00945_);
  nor (_00948_, _00821_, _38502_);
  and (_00949_, _00821_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_00950_, _00949_, _00806_);
  or (_00951_, _00950_, _00948_);
  or (_00952_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_00953_, _00952_, _41894_);
  and (_39726_, _00953_, _00951_);
  nor (_00954_, _00821_, _38494_);
  and (_00955_, _00821_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_00956_, _00955_, _00806_);
  or (_00957_, _00956_, _00954_);
  or (_00958_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_00959_, _00958_, _41894_);
  and (_39727_, _00959_, _00957_);
  nor (_00960_, _00821_, _38486_);
  and (_00961_, _00821_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_00962_, _00961_, _00806_);
  or (_00963_, _00962_, _00960_);
  or (_00964_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_00965_, _00964_, _41894_);
  and (_39729_, _00965_, _00963_);
  nor (_00966_, _00821_, _38479_);
  and (_00967_, _00821_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_00968_, _00967_, _00806_);
  or (_00969_, _00968_, _00966_);
  or (_00970_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_00971_, _00970_, _41894_);
  and (_39730_, _00971_, _00969_);
  nor (_00972_, _00821_, _38472_);
  and (_00973_, _00821_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_00974_, _00973_, _00806_);
  or (_00975_, _00974_, _00972_);
  or (_00976_, _40359_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_00977_, _00976_, _41894_);
  and (_39731_, _00977_, _00975_);
  nor (_00978_, _40632_, _40410_);
  nor (_00979_, _40551_, _40682_);
  and (_00980_, _00979_, _40467_);
  and (_00981_, _00980_, _00978_);
  not (_00982_, _40506_);
  nor (_00983_, _39187_, _39171_);
  and (_00984_, _39187_, _39171_);
  nor (_00985_, _00984_, _00983_);
  and (_00986_, _39159_, _39146_);
  nor (_00987_, _39159_, _39146_);
  or (_00988_, _00987_, _00986_);
  nor (_00989_, _00988_, _00985_);
  and (_00990_, _00988_, _00985_);
  nor (_00991_, _00990_, _00989_);
  nor (_00992_, _39211_, _39199_);
  and (_00993_, _39211_, _39199_);
  nor (_00994_, _00993_, _00992_);
  not (_00995_, _39134_);
  nor (_00996_, _39223_, _00995_);
  and (_00997_, _39223_, _00995_);
  nor (_00998_, _00997_, _00996_);
  nor (_00999_, _00998_, _00994_);
  and (_01000_, _00998_, _00994_);
  or (_01001_, _01000_, _00999_);
  or (_01002_, _01001_, _00991_);
  nand (_01003_, _01001_, _00991_);
  and (_01004_, _01003_, _01002_);
  or (_01005_, _01004_, _00982_);
  and (_01006_, _40586_, _40778_);
  or (_01007_, _40506_, _39080_);
  and (_01008_, _01007_, _01006_);
  and (_01009_, _01008_, _01005_);
  nor (_01010_, _40586_, _40778_);
  and (_01011_, _01010_, _40506_);
  and (_01012_, _01011_, _39070_);
  not (_01013_, _40586_);
  and (_01014_, _01013_, _40778_);
  or (_01015_, _40506_, _39087_);
  or (_01016_, _00982_, _38988_);
  and (_01017_, _01016_, _01015_);
  and (_01018_, _01017_, _01014_);
  and (_01019_, _01010_, _00982_);
  and (_01020_, _01019_, _38952_);
  or (_01021_, _01020_, _01018_);
  or (_01022_, _01021_, _01012_);
  or (_01023_, _00982_, _39032_);
  nor (_01024_, _01013_, _40778_);
  or (_01025_, _40506_, _39105_);
  and (_01026_, _01025_, _01024_);
  and (_01027_, _01026_, _01023_);
  or (_01028_, _01027_, _01022_);
  or (_01029_, _01028_, _01009_);
  and (_01030_, _01029_, _00981_);
  and (_01031_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_01032_, _01031_, _00982_);
  and (_01033_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01034_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01035_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_01036_, _01035_, _01034_);
  or (_01037_, _01036_, _01033_);
  or (_01038_, _01037_, _01032_);
  nor (_01039_, _40632_, _40467_);
  nor (_01040_, _40688_, _40410_);
  and (_01041_, _01040_, _40550_);
  and (_01042_, _01041_, _01039_);
  and (_01043_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_01044_, _01043_, _40506_);
  and (_01045_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01046_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01047_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_01048_, _01047_, _01046_);
  or (_01049_, _01048_, _01045_);
  or (_01050_, _01049_, _01044_);
  and (_01051_, _01050_, _01042_);
  and (_01052_, _01051_, _01038_);
  and (_01053_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_01054_, _01053_, _00982_);
  and (_01055_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_01056_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01057_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_01058_, _01057_, _01056_);
  or (_01059_, _01058_, _01055_);
  or (_01060_, _01059_, _01054_);
  not (_01061_, _40410_);
  and (_01062_, _00979_, _01061_);
  and (_01063_, _01062_, _01039_);
  and (_01064_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_01065_, _01064_, _40506_);
  and (_01066_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_01067_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01068_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_01069_, _01068_, _01067_);
  or (_01070_, _01069_, _01066_);
  or (_01071_, _01070_, _01065_);
  and (_01072_, _01071_, _01063_);
  and (_01073_, _01072_, _01060_);
  and (_01074_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_01075_, _01074_, _00982_);
  and (_01076_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_01077_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_01078_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_01079_, _01078_, _01077_);
  or (_01080_, _01079_, _01076_);
  or (_01081_, _01080_, _01075_);
  and (_01082_, _40632_, _01061_);
  nor (_01083_, _40688_, _40467_);
  and (_01084_, _01083_, _01082_);
  and (_01085_, _01084_, _40551_);
  and (_01086_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01087_, _01086_, _40506_);
  and (_01088_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_01089_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_01090_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01091_, _01090_, _01089_);
  or (_01092_, _01091_, _01088_);
  or (_01093_, _01092_, _01087_);
  and (_01094_, _01093_, _01085_);
  and (_01095_, _01094_, _01081_);
  or (_01096_, _01095_, _01073_);
  or (_01097_, _01096_, _01052_);
  not (_01098_, _38083_);
  and (_01099_, _42669_, _43221_);
  and (_01100_, _01099_, _01098_);
  nor (_01101_, _42643_, _37353_);
  and (_01102_, _37408_, _42642_);
  nor (_01103_, _01102_, _42665_);
  and (_01104_, _01103_, _01101_);
  and (_01105_, _38017_, _36785_);
  or (_01106_, _01105_, _42601_);
  or (_01107_, _01106_, _37233_);
  nor (_01108_, _01107_, _37786_);
  and (_01109_, _01108_, _01104_);
  and (_01110_, _01109_, _01100_);
  and (_01111_, _01110_, _42973_);
  and (_01112_, _01111_, _37659_);
  nor (_01113_, _01112_, _34314_);
  and (_01114_, _43156_, p0in_reg[0]);
  and (_01115_, _43152_, p0_in[0]);
  or (_01116_, _01115_, _01114_);
  or (_01117_, _01116_, _01113_);
  nand (_01118_, _01113_, _39483_);
  and (_01119_, _01118_, _01117_);
  and (_01120_, _01119_, _01006_);
  or (_01121_, _01120_, _00982_);
  and (_01122_, _43156_, p0in_reg[3]);
  and (_01123_, _43152_, p0_in[3]);
  or (_01124_, _01123_, _01122_);
  or (_01125_, _01124_, _01113_);
  nand (_01126_, _01113_, _39521_);
  and (_01127_, _01126_, _01125_);
  and (_01128_, _01127_, _01010_);
  and (_01129_, _43156_, p0in_reg[1]);
  and (_01130_, _43152_, p0_in[1]);
  or (_01131_, _01130_, _01129_);
  or (_01132_, _01131_, _01113_);
  not (_01133_, _01113_);
  or (_01134_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01135_, _01134_, _01132_);
  and (_01136_, _01135_, _01014_);
  and (_01137_, _43156_, p0in_reg[2]);
  and (_01138_, _43152_, p0_in[2]);
  or (_01139_, _01138_, _01137_);
  or (_01140_, _01139_, _01113_);
  or (_01141_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_01142_, _01141_, _01140_);
  and (_01143_, _01142_, _01024_);
  or (_01144_, _01143_, _01136_);
  or (_01145_, _01144_, _01128_);
  or (_01146_, _01145_, _01121_);
  and (_01147_, _40632_, _40467_);
  and (_01148_, _01147_, _01041_);
  and (_01149_, _43156_, p0in_reg[4]);
  and (_01150_, _43152_, p0_in[4]);
  or (_01151_, _01150_, _01149_);
  or (_01152_, _01151_, _01113_);
  or (_01153_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01154_, _01153_, _01152_);
  and (_01155_, _01154_, _01006_);
  or (_01156_, _01155_, _40506_);
  and (_01157_, _43156_, p0in_reg[7]);
  and (_01158_, _43152_, p0_in[7]);
  or (_01159_, _01158_, _01157_);
  or (_01160_, _01159_, _01113_);
  or (_01161_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_01162_, _01161_, _01160_);
  and (_01163_, _01162_, _01010_);
  and (_01164_, _43156_, p0in_reg[5]);
  and (_01165_, _43152_, p0_in[5]);
  or (_01166_, _01165_, _01164_);
  or (_01167_, _01166_, _01113_);
  or (_01168_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01169_, _01168_, _01167_);
  and (_01170_, _01169_, _01014_);
  and (_01171_, _43156_, p0in_reg[6]);
  and (_01172_, _43152_, p0_in[6]);
  or (_01173_, _01172_, _01171_);
  or (_01174_, _01173_, _01113_);
  or (_01175_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_01176_, _01175_, _01174_);
  and (_01177_, _01176_, _01024_);
  or (_01178_, _01177_, _01170_);
  or (_01179_, _01178_, _01163_);
  or (_01180_, _01179_, _01156_);
  and (_01181_, _01180_, _01148_);
  and (_01182_, _01181_, _01146_);
  and (_01183_, _43156_, p2in_reg[0]);
  and (_01184_, _43152_, p2_in[0]);
  or (_01185_, _01184_, _01183_);
  or (_01186_, _01185_, _01113_);
  or (_01187_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_01188_, _01187_, _01186_);
  and (_01189_, _01188_, _01006_);
  or (_01190_, _01189_, _00982_);
  and (_01191_, _43156_, p2in_reg[3]);
  and (_01192_, _43152_, p2_in[3]);
  or (_01193_, _01192_, _01191_);
  or (_01194_, _01193_, _01113_);
  or (_01195_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_01196_, _01195_, _01194_);
  and (_01197_, _01196_, _01010_);
  and (_01198_, _43156_, p2in_reg[2]);
  and (_01199_, _43152_, p2_in[2]);
  or (_01200_, _01199_, _01198_);
  or (_01201_, _01200_, _01113_);
  or (_01202_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_01203_, _01202_, _01201_);
  and (_01204_, _01203_, _01024_);
  and (_01205_, _43156_, p2in_reg[1]);
  and (_01206_, _43152_, p2_in[1]);
  or (_01207_, _01206_, _01205_);
  or (_01208_, _01207_, _01113_);
  or (_01209_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_01210_, _01209_, _01208_);
  and (_01211_, _01210_, _01014_);
  or (_01212_, _01211_, _01204_);
  or (_01213_, _01212_, _01197_);
  or (_01214_, _01213_, _01190_);
  and (_01215_, _01084_, _40550_);
  and (_01216_, _43156_, p2in_reg[4]);
  and (_01217_, _43152_, p2_in[4]);
  or (_01218_, _01217_, _01216_);
  or (_01219_, _01218_, _01113_);
  or (_01220_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_01221_, _01220_, _01219_);
  and (_01222_, _01221_, _01006_);
  or (_01223_, _01222_, _40506_);
  and (_01224_, _43156_, p2in_reg[7]);
  and (_01225_, _43152_, p2_in[7]);
  or (_01226_, _01225_, _01224_);
  or (_01227_, _01226_, _01113_);
  or (_01228_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_01229_, _01228_, _01227_);
  and (_01230_, _01229_, _01010_);
  and (_01231_, _43156_, p2in_reg[6]);
  and (_01232_, _43152_, p2_in[6]);
  or (_01233_, _01232_, _01231_);
  or (_01234_, _01233_, _01113_);
  or (_01235_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_01236_, _01235_, _01234_);
  and (_01237_, _01236_, _01024_);
  and (_01238_, _43156_, p2in_reg[5]);
  and (_01239_, _43152_, p2_in[5]);
  or (_01240_, _01239_, _01238_);
  or (_01241_, _01240_, _01113_);
  or (_01242_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01243_, _01242_, _01241_);
  and (_01244_, _01243_, _01014_);
  or (_01245_, _01244_, _01237_);
  or (_01246_, _01245_, _01230_);
  or (_01247_, _01246_, _01223_);
  and (_01248_, _01247_, _01215_);
  and (_01249_, _01248_, _01214_);
  or (_01250_, _01249_, _01182_);
  and (_01251_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_01252_, _01251_, _00982_);
  and (_01253_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_01254_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_01255_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_01256_, _01255_, _01254_);
  or (_01257_, _01256_, _01253_);
  or (_01258_, _01257_, _01252_);
  and (_01259_, _01147_, _01040_);
  and (_01260_, _01259_, _40551_);
  and (_01261_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_01262_, _01261_, _40506_);
  and (_01263_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_01264_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_01265_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_01266_, _01265_, _01264_);
  or (_01267_, _01266_, _01263_);
  or (_01268_, _01267_, _01262_);
  and (_01269_, _01268_, _01260_);
  and (_01270_, _01269_, _01258_);
  and (_01271_, _43156_, p1in_reg[1]);
  and (_01272_, _43152_, p1_in[1]);
  or (_01273_, _01272_, _01271_);
  or (_01274_, _01273_, _01113_);
  or (_01275_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_01276_, _01275_, _01274_);
  and (_01277_, _01276_, _01014_);
  or (_01278_, _01277_, _00982_);
  and (_01279_, _43156_, p1in_reg[3]);
  and (_01280_, _43152_, p1_in[3]);
  or (_01281_, _01280_, _01279_);
  or (_01282_, _01281_, _01113_);
  or (_01283_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_01284_, _01283_, _01282_);
  and (_01285_, _01284_, _01010_);
  and (_01286_, _43156_, p1in_reg[2]);
  and (_01287_, _43152_, p1_in[2]);
  or (_01288_, _01287_, _01286_);
  or (_01289_, _01288_, _01113_);
  or (_01290_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_01291_, _01290_, _01289_);
  and (_01292_, _01291_, _01024_);
  and (_01293_, _43156_, p1in_reg[0]);
  and (_01294_, _43152_, p1_in[0]);
  or (_01295_, _01294_, _01293_);
  or (_01296_, _01295_, _01113_);
  or (_01297_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_01298_, _01297_, _01296_);
  and (_01299_, _01298_, _01006_);
  or (_01300_, _01299_, _01292_);
  or (_01301_, _01300_, _01285_);
  or (_01302_, _01301_, _01278_);
  and (_01303_, _01082_, _00980_);
  and (_01304_, _43156_, p1in_reg[5]);
  and (_01305_, _43152_, p1_in[5]);
  or (_01306_, _01305_, _01304_);
  or (_01307_, _01306_, _01113_);
  or (_01308_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01309_, _01308_, _01307_);
  and (_01310_, _01309_, _01014_);
  or (_01311_, _01310_, _40506_);
  and (_01312_, _43156_, p1in_reg[7]);
  and (_01313_, _43152_, p1_in[7]);
  or (_01314_, _01313_, _01312_);
  or (_01315_, _01314_, _01113_);
  or (_01316_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_01317_, _01316_, _01315_);
  and (_01318_, _01317_, _01010_);
  and (_01319_, _43156_, p1in_reg[6]);
  and (_01320_, _43152_, p1_in[6]);
  or (_01321_, _01320_, _01319_);
  or (_01322_, _01321_, _01113_);
  or (_01323_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_01324_, _01323_, _01322_);
  and (_01325_, _01324_, _01024_);
  and (_01326_, _43156_, p1in_reg[4]);
  and (_01327_, _43152_, p1_in[4]);
  or (_01328_, _01327_, _01326_);
  or (_01329_, _01328_, _01113_);
  or (_01330_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01331_, _01330_, _01329_);
  and (_01332_, _01331_, _01006_);
  or (_01333_, _01332_, _01325_);
  or (_01334_, _01333_, _01318_);
  or (_01335_, _01334_, _01311_);
  and (_01336_, _01335_, _01303_);
  and (_01337_, _01336_, _01302_);
  or (_01338_, _01337_, _01270_);
  or (_01339_, _01338_, _01250_);
  or (_01340_, _01339_, _01097_);
  not (_01341_, _01215_);
  and (_01342_, _01062_, _40632_);
  nor (_01343_, _01342_, _01148_);
  and (_01344_, _01343_, _01341_);
  or (_01345_, _01042_, _00981_);
  nor (_01346_, _01345_, _01063_);
  nor (_01347_, _40550_, _40410_);
  and (_01348_, _40632_, _40682_);
  and (_01349_, _01348_, _01347_);
  and (_01350_, _40632_, _40688_);
  and (_01351_, _01350_, _01347_);
  nor (_01352_, _01351_, _01349_);
  and (_01353_, _01352_, _01346_);
  and (_01354_, _01353_, _01344_);
  nand (_01355_, _43271_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_01356_, _01355_, _01354_);
  and (_01357_, _43156_, p3in_reg[6]);
  and (_01358_, _43152_, p3_in[6]);
  or (_01359_, _01358_, _01357_);
  or (_01360_, _01359_, _01113_);
  or (_01361_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_01363_, _01361_, _01360_);
  nand (_01365_, _01363_, _01024_);
  and (_01367_, _01365_, _00982_);
  and (_01369_, _43156_, p3in_reg[7]);
  and (_01371_, _43152_, p3_in[7]);
  or (_01373_, _01371_, _01369_);
  or (_01375_, _01373_, _01113_);
  or (_01376_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_01377_, _01376_, _01375_);
  nand (_01378_, _01377_, _01010_);
  and (_01379_, _43156_, p3in_reg[5]);
  and (_01380_, _43152_, p3_in[5]);
  or (_01381_, _01380_, _01379_);
  or (_01383_, _01381_, _01113_);
  or (_01384_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01386_, _01384_, _01383_);
  nand (_01387_, _01386_, _01014_);
  and (_01388_, _43156_, p3in_reg[4]);
  and (_01390_, _43152_, p3_in[4]);
  or (_01391_, _01390_, _01388_);
  or (_01392_, _01391_, _01113_);
  or (_01394_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_01395_, _01394_, _01392_);
  nand (_01396_, _01395_, _01006_);
  and (_01398_, _01396_, _01387_);
  and (_01399_, _01398_, _01378_);
  and (_01400_, _01399_, _01367_);
  and (_01402_, _43156_, p3in_reg[2]);
  and (_01403_, _43152_, p3_in[2]);
  or (_01404_, _01403_, _01402_);
  or (_01406_, _01404_, _01113_);
  or (_01407_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_01408_, _01407_, _01406_);
  and (_01410_, _01408_, _01024_);
  or (_01411_, _01410_, _00982_);
  and (_01412_, _43156_, p3in_reg[3]);
  and (_01414_, _43152_, p3_in[3]);
  or (_01415_, _01414_, _01412_);
  or (_01416_, _01415_, _01113_);
  or (_01417_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_01418_, _01417_, _01416_);
  and (_01419_, _01418_, _01010_);
  and (_01420_, _43156_, p3in_reg[1]);
  and (_01421_, _43152_, p3_in[1]);
  or (_01422_, _01421_, _01420_);
  or (_01423_, _01422_, _01113_);
  or (_01424_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_01425_, _01424_, _01423_);
  and (_01426_, _01425_, _01014_);
  and (_01427_, _43156_, p3in_reg[0]);
  and (_01428_, _43152_, p3_in[0]);
  or (_01429_, _01428_, _01427_);
  or (_01430_, _01429_, _01113_);
  or (_01431_, _01133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_01432_, _01431_, _01430_);
  and (_01433_, _01432_, _01006_);
  or (_01434_, _01433_, _01426_);
  or (_01436_, _01434_, _01419_);
  or (_01437_, _01436_, _01411_);
  nand (_01439_, _01437_, _01342_);
  or (_01440_, _01439_, _01400_);
  nand (_01441_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_01443_, _01441_, _40506_);
  nand (_01444_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nand (_01445_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nand (_01447_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01448_, _01447_, _01445_);
  and (_01449_, _01448_, _01444_);
  and (_01451_, _01449_, _01443_);
  and (_01452_, _01024_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_01453_, _01452_, _40506_);
  and (_01455_, _01010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_01456_, _01014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01457_, _01006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01459_, _01457_, _01456_);
  or (_01460_, _01459_, _01455_);
  or (_01461_, _01460_, _01453_);
  nand (_01463_, _01461_, _01351_);
  or (_01464_, _01463_, _01451_);
  and (_01465_, _01464_, _01440_);
  or (_01467_, _01465_, _40467_);
  nand (_01468_, _01467_, _01356_);
  or (_01469_, _01468_, _01340_);
  or (_01470_, _01469_, _01030_);
  and (_01471_, _01042_, _39110_);
  nor (_01472_, _01356_, _29767_);
  nor (_01473_, _01472_, _01471_);
  and (_01474_, _01473_, _01470_);
  and (_01475_, _01019_, _39134_);
  and (_01476_, _01014_, _39211_);
  or (_01477_, _01476_, _40506_);
  and (_01478_, _01006_, _39199_);
  and (_01479_, _01024_, _39223_);
  or (_01480_, _01479_, _01478_);
  or (_01481_, _01480_, _01477_);
  and (_01482_, _01024_, _39171_);
  and (_01483_, _01014_, _39159_);
  or (_01484_, _01483_, _00982_);
  or (_01485_, _01484_, _01482_);
  and (_01486_, _01006_, _39146_);
  not (_01487_, _01010_);
  nor (_01489_, _01487_, _39187_);
  or (_01490_, _01489_, _01486_);
  or (_01492_, _01490_, _01485_);
  and (_01493_, _01492_, _01481_);
  or (_01494_, _01493_, _01475_);
  and (_01496_, _01494_, _01471_);
  not (_01497_, _01354_);
  nor (_01498_, _01344_, _01113_);
  not (_01500_, _01498_);
  and (_01501_, _43178_, _38931_);
  and (_01502_, _01501_, _01500_);
  and (_01504_, _01502_, _01497_);
  or (_01505_, _01504_, _01496_);
  or (_01506_, _01505_, _01474_);
  and (_01508_, _01019_, _40355_);
  or (_01509_, _40506_, _40598_);
  nand (_01510_, _40506_, _38502_);
  and (_01512_, _01510_, _01509_);
  and (_01513_, _01512_, _01024_);
  nand (_01514_, _00982_, _38486_);
  nand (_01516_, _40506_, _38518_);
  and (_01517_, _01516_, _01006_);
  and (_01518_, _01517_, _01514_);
  or (_01520_, _01518_, _01513_);
  not (_01521_, _38494_);
  and (_01522_, _01011_, _01521_);
  nand (_01523_, _00982_, _38479_);
  nand (_01524_, _40506_, _38509_);
  and (_01525_, _01524_, _01014_);
  and (_01526_, _01525_, _01523_);
  or (_01527_, _01526_, _01522_);
  or (_01528_, _01527_, _01520_);
  nor (_01529_, _01528_, _01508_);
  nand (_01530_, _01529_, _01504_);
  and (_01531_, _01530_, _41894_);
  and (_39761_, _01531_, _01506_);
  and (_01532_, _01006_, _40506_);
  and (_01533_, _01532_, _01042_);
  and (_01534_, _01533_, _39107_);
  and (_01535_, _01148_, _01011_);
  and (_01536_, _01535_, _38592_);
  and (_01537_, _01532_, _00981_);
  and (_01538_, _01537_, _38945_);
  or (_01539_, _01538_, _01536_);
  nor (_01541_, _01539_, _01534_);
  nor (_01542_, _01541_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_01544_, _01542_);
  not (_01545_, _38957_);
  nor (_01546_, _01019_, _01545_);
  and (_01548_, _01546_, _43178_);
  and (_01549_, _01532_, _01471_);
  nor (_01550_, _01549_, _01548_);
  and (_01552_, _01550_, _43275_);
  and (_01553_, _01552_, _01544_);
  and (_01554_, _40550_, _40506_);
  and (_01556_, _01554_, _01259_);
  and (_01557_, _01556_, _01024_);
  and (_01558_, _01557_, _38592_);
  or (_01560_, _01558_, rst);
  nor (_39762_, _01560_, _01553_);
  nand (_01561_, _01558_, _28496_);
  or (_01563_, _01553_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_01564_, _01557_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_01565_, _40682_, _40467_);
  and (_01567_, _01565_, _01082_);
  and (_01568_, _01532_, _40551_);
  and (_01569_, _01568_, _01567_);
  and (_01571_, _01569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_01572_, _01571_, _01564_);
  and (_01573_, _01568_, _01084_);
  and (_01574_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_01575_, _01568_, _01259_);
  and (_01576_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_01577_, _01576_, _01574_);
  or (_01578_, _01577_, _01572_);
  and (_01579_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_01580_, _01554_, _01006_);
  and (_01581_, _01565_, _00978_);
  and (_01582_, _01581_, _01580_);
  and (_01583_, _01582_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_01584_, _01583_, _01579_);
  and (_01585_, _01580_, _01567_);
  and (_01586_, _01585_, _01377_);
  and (_01587_, _01554_, _01014_);
  and (_01588_, _01587_, _01259_);
  and (_01589_, _01588_, _38542_);
  or (_01590_, _01589_, _01586_);
  or (_01591_, _01590_, _01584_);
  or (_01593_, _01591_, _01578_);
  and (_01594_, _01533_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01596_, _01580_, _01084_);
  and (_01597_, _01596_, _01229_);
  and (_01598_, _40688_, _40467_);
  and (_01600_, _01082_, _01598_);
  and (_01601_, _01600_, _01580_);
  and (_01602_, _01601_, _01317_);
  or (_01604_, _01602_, _01597_);
  and (_01605_, _01537_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01606_, _01580_, _01259_);
  and (_01608_, _01606_, _01162_);
  or (_01609_, _01608_, _01605_);
  or (_01610_, _01609_, _01604_);
  or (_01612_, _01610_, _01594_);
  nor (_01613_, _01612_, _01593_);
  nand (_01614_, _01613_, _01553_);
  and (_01616_, _01614_, _01563_);
  or (_01617_, _01616_, _01558_);
  and (_01618_, _01617_, _41894_);
  and (_39763_, _01618_, _01561_);
  and (_01620_, _01537_, _01004_);
  and (_01621_, _01557_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_01623_, _01532_, _01215_);
  and (_01624_, _01623_, _01188_);
  or (_01625_, _01624_, _01621_);
  and (_01626_, _01532_, _01148_);
  and (_01627_, _01626_, _01119_);
  and (_01628_, _01556_, _01014_);
  and (_01629_, _01628_, _40553_);
  or (_01630_, _01629_, _01627_);
  or (_01631_, _01630_, _01625_);
  and (_01632_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01633_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_01634_, _01582_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_01635_, _01532_, _01303_);
  and (_01636_, _01635_, _01298_);
  or (_01637_, _01636_, _01634_);
  or (_01638_, _01637_, _01633_);
  or (_01639_, _01638_, _01632_);
  and (_01640_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_01641_, _01569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01642_, _01585_, _01432_);
  and (_01643_, _01533_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_01645_, _01643_, _01642_);
  or (_01646_, _01645_, _01641_);
  or (_01648_, _01646_, _01640_);
  or (_01649_, _01648_, _01639_);
  nor (_01650_, _01649_, _01631_);
  nand (_01652_, _01650_, _01553_);
  or (_01653_, _01652_, _01620_);
  or (_01654_, _01553_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_01656_, _01654_, _01653_);
  or (_01657_, _01656_, _01558_);
  nand (_01658_, _01558_, _29679_);
  and (_01660_, _01658_, _41894_);
  and (_39825_, _01660_, _01657_);
  nand (_01661_, _01558_, _30358_);
  or (_01663_, _01553_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_01664_, _01557_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_01665_, _01569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_01667_, _01665_, _01664_);
  and (_01668_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_01669_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_01671_, _01669_, _01668_);
  or (_01672_, _01671_, _01667_);
  and (_01673_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_01675_, _01582_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_01676_, _01675_, _01673_);
  and (_01677_, _01585_, _01425_);
  and (_01678_, _01588_, _40706_);
  or (_01679_, _01678_, _01677_);
  or (_01680_, _01679_, _01676_);
  or (_01681_, _01680_, _01672_);
  and (_01682_, _01533_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01683_, _01596_, _01210_);
  and (_01684_, _01601_, _01276_);
  or (_01685_, _01684_, _01683_);
  and (_01686_, _01537_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_01687_, _01606_, _01135_);
  or (_01688_, _01687_, _01686_);
  or (_01689_, _01688_, _01685_);
  or (_01690_, _01689_, _01682_);
  nor (_01691_, _01690_, _01681_);
  nand (_01692_, _01691_, _01553_);
  and (_01693_, _01692_, _01663_);
  or (_01694_, _01693_, _01558_);
  and (_01695_, _01694_, _41894_);
  and (_39826_, _01695_, _01661_);
  not (_01697_, _01558_);
  and (_01699_, _01557_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_01700_, _01569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01701_, _01700_, _01699_);
  and (_01703_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_01704_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_01705_, _01704_, _01703_);
  or (_01707_, _01705_, _01701_);
  and (_01708_, _01582_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01709_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_01711_, _01709_, _01708_);
  and (_01712_, _01585_, _01408_);
  and (_01713_, _01588_, _40470_);
  or (_01715_, _01713_, _01712_);
  or (_01716_, _01715_, _01711_);
  or (_01717_, _01716_, _01707_);
  and (_01719_, _01533_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01720_, _01596_, _01203_);
  and (_01721_, _01601_, _01291_);
  or (_01723_, _01721_, _01720_);
  and (_01724_, _01537_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_01725_, _01606_, _01142_);
  or (_01727_, _01725_, _01724_);
  or (_01728_, _01727_, _01723_);
  or (_01729_, _01728_, _01719_);
  or (_01730_, _01729_, _01717_);
  and (_01731_, _01730_, _01553_);
  nor (_01732_, _01553_, _16436_);
  or (_01733_, _01732_, _01731_);
  and (_01734_, _01733_, _01697_);
  nor (_01735_, _01697_, _31069_);
  or (_01736_, _01735_, _01734_);
  and (_39828_, _01736_, _41894_);
  and (_01737_, _01569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_01738_, _01557_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_01739_, _01738_, _01737_);
  and (_01740_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_01741_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_01742_, _01741_, _01740_);
  or (_01743_, _01742_, _01739_);
  and (_01744_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_01745_, _01582_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_01746_, _01745_, _01744_);
  and (_01748_, _01585_, _01418_);
  and (_01749_, _01588_, _40515_);
  or (_01751_, _01749_, _01748_);
  or (_01752_, _01751_, _01746_);
  or (_01753_, _01752_, _01743_);
  and (_01755_, _01533_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01756_, _01596_, _01196_);
  and (_01757_, _01601_, _01284_);
  or (_01759_, _01757_, _01756_);
  and (_01760_, _01537_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_01761_, _01606_, _01127_);
  or (_01763_, _01761_, _01760_);
  or (_01764_, _01763_, _01759_);
  or (_01765_, _01764_, _01755_);
  or (_01767_, _01765_, _01753_);
  and (_01768_, _01767_, _01553_);
  nor (_01769_, _01553_, _17465_);
  or (_01771_, _01769_, _01768_);
  and (_01772_, _01771_, _01697_);
  nor (_01773_, _01697_, _31822_);
  or (_01775_, _01773_, _01772_);
  and (_39829_, _01775_, _41894_);
  and (_01776_, _01557_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_01778_, _01569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01779_, _01778_, _01776_);
  and (_01780_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_01781_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_01782_, _01781_, _01780_);
  or (_01783_, _01782_, _01779_);
  and (_01784_, _01582_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01785_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_01786_, _01785_, _01784_);
  and (_01787_, _01585_, _01395_);
  and (_01788_, _01588_, _40643_);
  or (_01789_, _01788_, _01787_);
  or (_01790_, _01789_, _01786_);
  or (_01791_, _01790_, _01783_);
  and (_01792_, _01533_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01793_, _01596_, _01221_);
  and (_01794_, _01601_, _01331_);
  or (_01795_, _01794_, _01793_);
  and (_01796_, _01537_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01797_, _01606_, _01154_);
  or (_01798_, _01797_, _01796_);
  or (_01800_, _01798_, _01795_);
  or (_01801_, _01800_, _01792_);
  or (_01803_, _01801_, _01791_);
  and (_01804_, _01803_, _01553_);
  nor (_01805_, _01553_, _16634_);
  or (_01807_, _01805_, _01804_);
  and (_01808_, _01807_, _01697_);
  nor (_01809_, _01697_, _32585_);
  or (_01811_, _01809_, _01808_);
  and (_39830_, _01811_, _41894_);
  and (_01812_, _01569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01814_, _01557_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_01815_, _01814_, _01812_);
  and (_01816_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_01818_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_01819_, _01818_, _01816_);
  or (_01820_, _01819_, _01815_);
  and (_01822_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_01823_, _01582_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_01824_, _01823_, _01822_);
  and (_01826_, _01585_, _01386_);
  and (_01827_, _01588_, _40448_);
  or (_01828_, _01827_, _01826_);
  or (_01830_, _01828_, _01824_);
  or (_01831_, _01830_, _01820_);
  and (_01832_, _01533_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01833_, _01596_, _01243_);
  and (_01834_, _01601_, _01309_);
  or (_01835_, _01834_, _01833_);
  and (_01836_, _01537_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01837_, _01606_, _01169_);
  or (_01838_, _01837_, _01836_);
  or (_01839_, _01838_, _01835_);
  or (_01840_, _01839_, _01832_);
  or (_01841_, _01840_, _01831_);
  and (_01842_, _01841_, _01553_);
  nor (_01843_, _01553_, _17617_);
  or (_01844_, _01843_, _01842_);
  and (_01845_, _01844_, _01697_);
  nor (_01846_, _01697_, _33379_);
  or (_01847_, _01846_, _01845_);
  and (_39831_, _01847_, _41894_);
  and (_01848_, _01557_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01849_, _01569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_01851_, _01849_, _01848_);
  and (_01852_, _01575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_01854_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_01855_, _01854_, _01852_);
  or (_01856_, _01855_, _01851_);
  and (_01858_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_01859_, _01582_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_01860_, _01859_, _01858_);
  and (_01862_, _01585_, _01363_);
  and (_01863_, _01588_, _40629_);
  or (_01864_, _01863_, _01862_);
  or (_01866_, _01864_, _01860_);
  or (_01867_, _01866_, _01856_);
  and (_01868_, _01533_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01870_, _01596_, _01236_);
  and (_01871_, _01601_, _01324_);
  or (_01872_, _01871_, _01870_);
  and (_01874_, _01537_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01875_, _01606_, _01176_);
  or (_01876_, _01875_, _01874_);
  or (_01878_, _01876_, _01872_);
  or (_01879_, _01878_, _01868_);
  or (_01880_, _01879_, _01867_);
  and (_01882_, _01880_, _01553_);
  nor (_01883_, _01553_, _16974_);
  or (_01884_, _01883_, _01882_);
  and (_01885_, _01884_, _01697_);
  nor (_01886_, _01697_, _34098_);
  or (_01887_, _01886_, _01885_);
  and (_39832_, _01887_, _41894_);
  and (_39876_, _40827_, _41894_);
  and (_39878_, _40965_, _41894_);
  nor (_39880_, _40506_, rst);
  and (_39895_, _40982_, _41894_);
  and (_39896_, _40997_, _41894_);
  and (_39897_, _41008_, _41894_);
  and (_39899_, _41016_, _41894_);
  and (_39900_, _41027_, _41894_);
  and (_39901_, _41038_, _41894_);
  and (_39902_, _41049_, _41894_);
  nor (_39903_, _40586_, rst);
  nor (_39904_, _40778_, rst);
  nor (_01888_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01890_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01891_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01890_);
  nor (_01893_, _01891_, _01888_);
  nor (_01894_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01895_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01890_);
  nor (_01897_, _01895_, _01894_);
  nor (_01898_, _01897_, _01893_);
  nor (_01899_, _00152_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01901_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01890_);
  nor (_01902_, _01901_, _01899_);
  and (_01903_, _01902_, _01898_);
  nor (_01905_, _00172_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01906_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01890_);
  nor (_01907_, _01906_, _01905_);
  and (_01909_, _01907_, _01903_);
  and (_01910_, _01909_, _42427_);
  not (_01911_, _42345_);
  not (_01913_, _01897_);
  nor (_01914_, _01913_, _01893_);
  not (_01915_, _01898_);
  and (_01917_, _01902_, _01915_);
  nor (_01918_, _01902_, _01915_);
  nor (_01919_, _01918_, _01917_);
  and (_01921_, _01907_, _01919_);
  and (_01922_, _01921_, _01914_);
  and (_01923_, _01922_, _01911_);
  not (_01924_, _42386_);
  and (_01925_, _01897_, _01893_);
  and (_01926_, _01921_, _01925_);
  and (_01927_, _01926_, _01924_);
  or (_01928_, _01927_, _01923_);
  not (_01929_, _42304_);
  and (_01930_, _01913_, _01893_);
  and (_01931_, _01921_, _01930_);
  and (_01932_, _01931_, _01929_);
  not (_01933_, _42263_);
  and (_01934_, _01907_, _01918_);
  and (_01935_, _01934_, _01933_);
  or (_01936_, _01935_, _01932_);
  or (_01937_, _01936_, _01928_);
  not (_01938_, _42222_);
  not (_01939_, _01919_);
  nor (_01940_, _01907_, _01917_);
  and (_01941_, _01907_, _01917_);
  nor (_01943_, _01941_, _01940_);
  and (_01944_, _01943_, _01939_);
  and (_01946_, _01944_, _01925_);
  and (_01947_, _01946_, _01938_);
  not (_01948_, _42181_);
  and (_01950_, _01914_, _01944_);
  and (_01951_, _01950_, _01948_);
  or (_01952_, _01951_, _01947_);
  not (_01954_, _42140_);
  and (_01955_, _01930_, _01944_);
  and (_01956_, _01955_, _01954_);
  not (_01958_, _42099_);
  nor (_01959_, _01907_, _01939_);
  and (_01960_, _01959_, _01898_);
  and (_01962_, _01960_, _01958_);
  or (_01963_, _01962_, _01956_);
  or (_01964_, _01963_, _01952_);
  or (_01966_, _01964_, _01937_);
  not (_01967_, _42017_);
  and (_01968_, _01959_, _01914_);
  and (_01970_, _01968_, _01967_);
  not (_01971_, _42058_);
  and (_01972_, _01959_, _01925_);
  and (_01974_, _01972_, _01971_);
  or (_01975_, _01974_, _01970_);
  not (_01976_, _41935_);
  nor (_01977_, _01943_, _01919_);
  and (_01978_, _01977_, _01898_);
  and (_01979_, _01978_, _01976_);
  not (_01980_, _41976_);
  and (_01981_, _01959_, _01930_);
  and (_01982_, _01981_, _01980_);
  or (_01983_, _01982_, _01979_);
  or (_01984_, _01983_, _01975_);
  not (_01985_, _41797_);
  and (_01986_, _01930_, _01977_);
  and (_01987_, _01986_, _01985_);
  not (_01988_, _41840_);
  and (_01989_, _01977_, _01914_);
  and (_01990_, _01989_, _01988_);
  not (_01991_, _41893_);
  and (_01992_, _01977_, _01925_);
  and (_01993_, _01992_, _01991_);
  or (_01994_, _01993_, _01990_);
  or (_01996_, _01994_, _01987_);
  or (_01997_, _01996_, _01984_);
  or (_01999_, _01997_, _01966_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01999_, _01910_);
  and (_02000_, _01989_, _42427_);
  and (_02002_, _01926_, _01929_);
  and (_02003_, _01922_, _01933_);
  or (_02004_, _02003_, _02002_);
  and (_02006_, _01986_, _01924_);
  and (_02007_, _01909_, _01911_);
  or (_02008_, _02007_, _02006_);
  or (_02010_, _02008_, _02004_);
  and (_02011_, _01934_, _01948_);
  and (_02012_, _01931_, _01938_);
  or (_02014_, _02012_, _02011_);
  and (_02015_, _01950_, _01958_);
  and (_02016_, _01946_, _01954_);
  or (_02018_, _02016_, _02015_);
  or (_02019_, _02018_, _02014_);
  or (_02020_, _02019_, _02010_);
  and (_02022_, _01968_, _01976_);
  and (_02023_, _01972_, _01980_);
  or (_02024_, _02023_, _02022_);
  and (_02026_, _01960_, _01967_);
  and (_02027_, _01955_, _01971_);
  or (_02028_, _02027_, _02026_);
  or (_02029_, _02028_, _02024_);
  and (_02030_, _01992_, _01985_);
  and (_02031_, _01981_, _01991_);
  and (_02032_, _01978_, _01988_);
  or (_02033_, _02032_, _02031_);
  or (_02034_, _02033_, _02030_);
  or (_02035_, _02034_, _02029_);
  or (_02036_, _02035_, _02020_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _02036_, _02000_);
  and (_02037_, _01986_, _42427_);
  and (_02038_, _01972_, _01967_);
  and (_02039_, _01960_, _01971_);
  or (_02040_, _02039_, _02038_);
  and (_02041_, _01968_, _01980_);
  and (_02042_, _01981_, _01976_);
  or (_02043_, _02042_, _02041_);
  or (_02044_, _02043_, _02040_);
  and (_02045_, _01989_, _01985_);
  and (_02047_, _01978_, _01991_);
  and (_02048_, _01992_, _01988_);
  or (_02050_, _02048_, _02047_);
  or (_02051_, _02050_, _02045_);
  or (_02052_, _02051_, _02044_);
  and (_02054_, _01922_, _01929_);
  and (_02055_, _01931_, _01933_);
  or (_02056_, _02055_, _02054_);
  and (_02058_, _01926_, _01911_);
  and (_02059_, _01909_, _01924_);
  or (_02060_, _02059_, _02058_);
  or (_02062_, _02060_, _02056_);
  and (_02063_, _01950_, _01954_);
  and (_02064_, _01955_, _01958_);
  or (_02066_, _02064_, _02063_);
  and (_02067_, _01946_, _01948_);
  and (_02068_, _01934_, _01938_);
  or (_02070_, _02068_, _02067_);
  or (_02071_, _02070_, _02066_);
  or (_02072_, _02071_, _02062_);
  or (_02074_, _02072_, _02052_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _02074_, _02037_);
  and (_02075_, _01992_, _42427_);
  and (_02077_, _01934_, _01954_);
  and (_02078_, _01946_, _01958_);
  and (_02079_, _01931_, _01948_);
  and (_02080_, _01922_, _01938_);
  or (_02081_, _02080_, _02079_);
  or (_02082_, _02081_, _02078_);
  or (_02083_, _02082_, _02077_);
  and (_02084_, _01989_, _01924_);
  and (_02085_, _01986_, _01911_);
  or (_02086_, _02085_, _02084_);
  and (_02087_, _01926_, _01933_);
  and (_02088_, _01909_, _01929_);
  or (_02089_, _02088_, _02087_);
  or (_02090_, _02089_, _02086_);
  or (_02091_, _02090_, _02083_);
  and (_02092_, _01981_, _01988_);
  and (_02093_, _01968_, _01991_);
  and (_02094_, _01978_, _01985_);
  or (_02095_, _02094_, _02093_);
  or (_02096_, _02095_, _02092_);
  and (_02097_, _01960_, _01980_);
  and (_02099_, _01972_, _01976_);
  or (_02100_, _02099_, _02097_);
  and (_02102_, _01950_, _01971_);
  and (_02103_, _01955_, _01967_);
  or (_02104_, _02103_, _02102_);
  or (_02106_, _02104_, _02100_);
  or (_02107_, _02106_, _02096_);
  or (_02108_, _02107_, _02091_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _02108_, _02075_);
  and (_02110_, _01989_, _42432_);
  not (_02111_, _42145_);
  and (_02113_, _01946_, _02111_);
  not (_02114_, _42104_);
  and (_02115_, _01950_, _02114_);
  or (_02117_, _02115_, _02113_);
  not (_02118_, _42186_);
  and (_02119_, _01934_, _02118_);
  not (_02121_, _42227_);
  and (_02122_, _01931_, _02121_);
  or (_02123_, _02122_, _02119_);
  or (_02125_, _02123_, _02117_);
  not (_02126_, _42309_);
  and (_02127_, _01926_, _02126_);
  not (_02129_, _42268_);
  and (_02130_, _01922_, _02129_);
  or (_02131_, _02130_, _02127_);
  not (_02132_, _42350_);
  and (_02133_, _01909_, _02132_);
  not (_02134_, _42391_);
  and (_02135_, _01986_, _02134_);
  or (_02136_, _02135_, _02133_);
  or (_02137_, _02136_, _02131_);
  or (_02138_, _02137_, _02125_);
  not (_02139_, _41981_);
  and (_02140_, _01972_, _02139_);
  not (_02141_, _41940_);
  and (_02142_, _01968_, _02141_);
  or (_02143_, _02142_, _02140_);
  not (_02144_, _42063_);
  and (_02145_, _01955_, _02144_);
  not (_02146_, _42022_);
  and (_02147_, _01960_, _02146_);
  or (_02148_, _02147_, _02145_);
  or (_02149_, _02148_, _02143_);
  not (_02151_, _41802_);
  and (_02152_, _01992_, _02151_);
  not (_02154_, _41899_);
  and (_02155_, _01981_, _02154_);
  not (_02156_, _41850_);
  and (_02158_, _01978_, _02156_);
  or (_02159_, _02158_, _02155_);
  or (_02160_, _02159_, _02152_);
  or (_02162_, _02160_, _02149_);
  or (_02163_, _02162_, _02138_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _02163_, _02110_);
  and (_02165_, _01989_, _42437_);
  not (_02166_, _42109_);
  and (_02167_, _01950_, _02166_);
  not (_02169_, _42150_);
  and (_02170_, _01946_, _02169_);
  or (_02171_, _02170_, _02167_);
  not (_02173_, _42191_);
  and (_02174_, _01934_, _02173_);
  not (_02175_, _42232_);
  and (_02177_, _01931_, _02175_);
  or (_02178_, _02177_, _02174_);
  or (_02179_, _02178_, _02171_);
  not (_02181_, _42314_);
  and (_02182_, _01926_, _02181_);
  not (_02183_, _42273_);
  and (_02184_, _01922_, _02183_);
  or (_02185_, _02184_, _02182_);
  not (_02186_, _42355_);
  and (_02187_, _01909_, _02186_);
  not (_02188_, _42396_);
  and (_02189_, _01986_, _02188_);
  or (_02190_, _02189_, _02187_);
  or (_02191_, _02190_, _02185_);
  or (_02192_, _02191_, _02179_);
  not (_02193_, _41986_);
  and (_02194_, _01972_, _02193_);
  not (_02195_, _41945_);
  and (_02196_, _01968_, _02195_);
  or (_02197_, _02196_, _02194_);
  not (_02198_, _42027_);
  and (_02199_, _01960_, _02198_);
  not (_02200_, _42068_);
  and (_02201_, _01955_, _02200_);
  or (_02202_, _02201_, _02199_);
  or (_02203_, _02202_, _02197_);
  not (_02204_, _41807_);
  and (_02205_, _01992_, _02204_);
  not (_02206_, _41904_);
  and (_02207_, _01981_, _02206_);
  not (_02208_, _41855_);
  and (_02209_, _01978_, _02208_);
  or (_02210_, _02209_, _02207_);
  or (_02211_, _02210_, _02205_);
  or (_02212_, _02211_, _02203_);
  or (_02213_, _02212_, _02192_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _02213_, _02165_);
  not (_02214_, _42401_);
  and (_02215_, _01986_, _02214_);
  not (_02216_, _42278_);
  and (_02217_, _01922_, _02216_);
  not (_02218_, _42319_);
  and (_02219_, _01926_, _02218_);
  or (_02220_, _02219_, _02217_);
  or (_02221_, _02220_, _02215_);
  not (_02222_, _42155_);
  and (_02223_, _01946_, _02222_);
  and (_02224_, _01989_, _42442_);
  or (_02225_, _02224_, _02223_);
  or (_02226_, _02225_, _02221_);
  not (_02227_, _42032_);
  and (_02228_, _01960_, _02227_);
  not (_02229_, _41950_);
  and (_02230_, _01968_, _02229_);
  not (_02231_, _41991_);
  and (_02232_, _01972_, _02231_);
  or (_02233_, _02232_, _02230_);
  or (_02234_, _02233_, _02228_);
  not (_02235_, _42073_);
  and (_02236_, _01955_, _02235_);
  not (_02237_, _41860_);
  and (_02238_, _01978_, _02237_);
  or (_02239_, _02238_, _02236_);
  or (_02240_, _02239_, _02234_);
  or (_02241_, _02240_, _02226_);
  not (_02242_, _42360_);
  and (_02243_, _01909_, _02242_);
  not (_02244_, _41812_);
  and (_02245_, _01992_, _02244_);
  not (_02246_, _41909_);
  and (_02247_, _01981_, _02246_);
  or (_02248_, _02247_, _02245_);
  not (_02249_, _42114_);
  and (_02250_, _01950_, _02249_);
  not (_02251_, _42237_);
  and (_02252_, _01931_, _02251_);
  not (_02253_, _42196_);
  and (_02254_, _01934_, _02253_);
  or (_02255_, _02254_, _02252_);
  or (_02256_, _02255_, _02250_);
  or (_02257_, _02256_, _02248_);
  or (_02258_, _02257_, _02243_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _02258_, _02241_);
  and (_02259_, _01989_, _42447_);
  not (_02260_, _42283_);
  and (_02261_, _01922_, _02260_);
  not (_02262_, _42324_);
  and (_02263_, _01926_, _02262_);
  or (_02264_, _02263_, _02261_);
  not (_02265_, _42406_);
  and (_02266_, _01986_, _02265_);
  not (_02267_, _42365_);
  and (_02268_, _01909_, _02267_);
  or (_02269_, _02268_, _02266_);
  or (_02270_, _02269_, _02264_);
  not (_02271_, _42201_);
  and (_02272_, _01934_, _02271_);
  not (_02273_, _42242_);
  and (_02274_, _01931_, _02273_);
  or (_02275_, _02274_, _02272_);
  not (_02276_, _42160_);
  and (_02277_, _01946_, _02276_);
  not (_02278_, _42119_);
  and (_02279_, _01950_, _02278_);
  or (_02280_, _02279_, _02277_);
  or (_02281_, _02280_, _02275_);
  or (_02282_, _02281_, _02270_);
  not (_02283_, _41817_);
  and (_02284_, _01992_, _02283_);
  not (_02285_, _41914_);
  and (_02286_, _01981_, _02285_);
  not (_02287_, _41865_);
  and (_02288_, _01978_, _02287_);
  or (_02289_, _02288_, _02286_);
  or (_02290_, _02289_, _02284_);
  not (_02291_, _41996_);
  and (_02292_, _01972_, _02291_);
  not (_02293_, _41955_);
  and (_02294_, _01968_, _02293_);
  or (_02295_, _02294_, _02292_);
  not (_02296_, _42078_);
  and (_02297_, _01955_, _02296_);
  not (_02298_, _42037_);
  and (_02299_, _01960_, _02298_);
  or (_02300_, _02299_, _02297_);
  or (_02301_, _02300_, _02295_);
  or (_02302_, _02301_, _02290_);
  or (_02303_, _02302_, _02282_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _02303_, _02259_);
  not (_02304_, _42411_);
  and (_02305_, _01986_, _02304_);
  not (_02306_, _42288_);
  and (_02307_, _01922_, _02306_);
  not (_02308_, _42329_);
  and (_02309_, _01926_, _02308_);
  or (_02310_, _02309_, _02307_);
  or (_02311_, _02310_, _02305_);
  not (_02312_, _42124_);
  and (_02313_, _01950_, _02312_);
  and (_02314_, _01989_, _42452_);
  or (_02315_, _02314_, _02313_);
  or (_02316_, _02315_, _02311_);
  not (_02317_, _42042_);
  and (_02318_, _01960_, _02317_);
  not (_02319_, _41960_);
  and (_02320_, _01968_, _02319_);
  not (_02321_, _42001_);
  and (_02322_, _01972_, _02321_);
  or (_02323_, _02322_, _02320_);
  or (_02324_, _02323_, _02318_);
  not (_02325_, _42083_);
  and (_02326_, _01955_, _02325_);
  not (_02327_, _41870_);
  and (_02328_, _01978_, _02327_);
  or (_02329_, _02328_, _02326_);
  or (_02330_, _02329_, _02324_);
  or (_02331_, _02330_, _02316_);
  not (_02332_, _42370_);
  and (_02333_, _01909_, _02332_);
  not (_02334_, _41822_);
  and (_02335_, _01992_, _02334_);
  not (_02336_, _41919_);
  and (_02337_, _01981_, _02336_);
  or (_02338_, _02337_, _02335_);
  not (_02339_, _42165_);
  and (_02340_, _01946_, _02339_);
  not (_02341_, _42247_);
  and (_02342_, _01931_, _02341_);
  not (_02343_, _42206_);
  and (_02344_, _01934_, _02343_);
  or (_02345_, _02344_, _02342_);
  or (_02346_, _02345_, _02340_);
  or (_02347_, _02346_, _02338_);
  or (_02348_, _02347_, _02333_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _02348_, _02331_);
  not (_02349_, _42416_);
  and (_02350_, _01986_, _02349_);
  not (_02351_, _42293_);
  and (_02352_, _01922_, _02351_);
  not (_02353_, _42334_);
  and (_02354_, _01926_, _02353_);
  or (_02355_, _02354_, _02352_);
  or (_02356_, _02355_, _02350_);
  not (_02357_, _42170_);
  and (_02358_, _01946_, _02357_);
  and (_02359_, _01989_, _42457_);
  or (_02360_, _02359_, _02358_);
  or (_02361_, _02360_, _02356_);
  not (_02362_, _42047_);
  and (_02363_, _01960_, _02362_);
  not (_02364_, _41965_);
  and (_02365_, _01968_, _02364_);
  not (_02366_, _42006_);
  and (_02367_, _01972_, _02366_);
  or (_02368_, _02367_, _02365_);
  or (_02369_, _02368_, _02363_);
  not (_02370_, _42088_);
  and (_02371_, _01955_, _02370_);
  not (_02372_, _41875_);
  and (_02373_, _01978_, _02372_);
  or (_02374_, _02373_, _02371_);
  or (_02375_, _02374_, _02369_);
  or (_02376_, _02375_, _02361_);
  not (_02377_, _42375_);
  and (_02378_, _01909_, _02377_);
  not (_02379_, _41827_);
  and (_02380_, _01992_, _02379_);
  not (_02381_, _41924_);
  and (_02382_, _01981_, _02381_);
  or (_02383_, _02382_, _02380_);
  not (_02384_, _42129_);
  and (_02385_, _01950_, _02384_);
  not (_02386_, _42252_);
  and (_02387_, _01931_, _02386_);
  not (_02388_, _42211_);
  and (_02389_, _01934_, _02388_);
  or (_02390_, _02389_, _02387_);
  or (_02391_, _02390_, _02385_);
  or (_02392_, _02391_, _02383_);
  or (_02393_, _02392_, _02378_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _02393_, _02376_);
  not (_02394_, _42421_);
  and (_02395_, _01986_, _02394_);
  not (_02396_, _42298_);
  and (_02397_, _01922_, _02396_);
  not (_02398_, _42339_);
  and (_02399_, _01926_, _02398_);
  or (_02400_, _02399_, _02397_);
  or (_02401_, _02400_, _02395_);
  not (_02402_, _42175_);
  and (_02403_, _01946_, _02402_);
  and (_02404_, _01989_, _42462_);
  or (_02405_, _02404_, _02403_);
  or (_02406_, _02405_, _02401_);
  not (_02407_, _42052_);
  and (_02408_, _01960_, _02407_);
  not (_02409_, _41970_);
  and (_02410_, _01968_, _02409_);
  not (_02411_, _42011_);
  and (_02412_, _01972_, _02411_);
  or (_02413_, _02412_, _02410_);
  or (_02414_, _02413_, _02408_);
  not (_02415_, _42093_);
  and (_02416_, _01955_, _02415_);
  not (_02417_, _41880_);
  and (_02418_, _01978_, _02417_);
  or (_02419_, _02418_, _02416_);
  or (_02420_, _02419_, _02414_);
  or (_02421_, _02420_, _02406_);
  not (_02422_, _42380_);
  and (_02423_, _01909_, _02422_);
  not (_02424_, _41832_);
  and (_02426_, _01992_, _02424_);
  not (_02427_, _41929_);
  and (_02428_, _01981_, _02427_);
  or (_02429_, _02428_, _02426_);
  not (_02430_, _42134_);
  and (_02431_, _01950_, _02430_);
  not (_02432_, _42257_);
  and (_02433_, _01931_, _02432_);
  not (_02434_, _42216_);
  and (_02435_, _01934_, _02434_);
  or (_02436_, _02435_, _02433_);
  or (_02437_, _02436_, _02431_);
  or (_02438_, _02437_, _02429_);
  or (_02439_, _02438_, _02423_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _02439_, _02421_);
  and (_02440_, _01909_, _42432_);
  and (_02441_, _01926_, _02134_);
  and (_02442_, _01922_, _02132_);
  or (_02443_, _02442_, _02441_);
  and (_02444_, _01931_, _02126_);
  and (_02445_, _01934_, _02129_);
  or (_02446_, _02445_, _02444_);
  or (_02447_, _02446_, _02443_);
  and (_02448_, _01946_, _02121_);
  and (_02449_, _01950_, _02118_);
  or (_02450_, _02449_, _02448_);
  and (_02451_, _01955_, _02111_);
  and (_02452_, _01960_, _02114_);
  or (_02453_, _02452_, _02451_);
  or (_02454_, _02453_, _02450_);
  or (_02455_, _02454_, _02447_);
  and (_02456_, _01968_, _02146_);
  and (_02457_, _01972_, _02144_);
  or (_02458_, _02457_, _02456_);
  and (_02459_, _01981_, _02139_);
  and (_02460_, _01978_, _02141_);
  or (_02461_, _02460_, _02459_);
  or (_02462_, _02461_, _02458_);
  and (_02463_, _01986_, _02151_);
  and (_02464_, _01989_, _02156_);
  and (_02465_, _01992_, _02154_);
  or (_02466_, _02465_, _02464_);
  or (_02467_, _02466_, _02463_);
  or (_02468_, _02467_, _02462_);
  or (_02469_, _02468_, _02455_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _02469_, _02440_);
  and (_02470_, _01909_, _42437_);
  and (_02471_, _01926_, _02188_);
  and (_02472_, _01922_, _02186_);
  or (_02473_, _02472_, _02471_);
  and (_02474_, _01931_, _02181_);
  and (_02475_, _01934_, _02183_);
  or (_02476_, _02475_, _02474_);
  or (_02477_, _02476_, _02473_);
  and (_02478_, _01950_, _02173_);
  and (_02479_, _01946_, _02175_);
  or (_02480_, _02479_, _02478_);
  and (_02481_, _01955_, _02169_);
  and (_02482_, _01960_, _02166_);
  or (_02483_, _02482_, _02481_);
  or (_02484_, _02483_, _02480_);
  or (_02485_, _02484_, _02477_);
  and (_02486_, _01972_, _02200_);
  and (_02487_, _01968_, _02198_);
  or (_02488_, _02487_, _02486_);
  and (_02489_, _01981_, _02193_);
  and (_02490_, _01978_, _02195_);
  or (_02491_, _02490_, _02489_);
  or (_02492_, _02491_, _02488_);
  and (_02493_, _01986_, _02204_);
  and (_02494_, _01992_, _02206_);
  and (_02495_, _01989_, _02208_);
  or (_02496_, _02495_, _02494_);
  or (_02497_, _02496_, _02493_);
  or (_02498_, _02497_, _02492_);
  or (_02499_, _02498_, _02485_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _02499_, _02470_);
  and (_02500_, _01909_, _42442_);
  and (_02501_, _01922_, _02242_);
  and (_02502_, _01926_, _02214_);
  or (_02503_, _02502_, _02501_);
  and (_02504_, _01931_, _02218_);
  and (_02505_, _01934_, _02216_);
  or (_02506_, _02505_, _02504_);
  or (_02507_, _02506_, _02503_);
  and (_02508_, _01946_, _02251_);
  and (_02509_, _01950_, _02253_);
  or (_02510_, _02509_, _02508_);
  and (_02511_, _01955_, _02222_);
  and (_02512_, _01960_, _02249_);
  or (_02513_, _02512_, _02511_);
  or (_02514_, _02513_, _02510_);
  or (_02515_, _02514_, _02507_);
  and (_02516_, _01972_, _02235_);
  and (_02517_, _01968_, _02227_);
  or (_02518_, _02517_, _02516_);
  and (_02519_, _01981_, _02231_);
  and (_02520_, _01978_, _02229_);
  or (_02521_, _02520_, _02519_);
  or (_02522_, _02521_, _02518_);
  and (_02523_, _01986_, _02244_);
  and (_02524_, _01992_, _02246_);
  and (_02525_, _01989_, _02237_);
  or (_02526_, _02525_, _02524_);
  or (_02527_, _02526_, _02523_);
  or (_02528_, _02527_, _02522_);
  or (_02529_, _02528_, _02515_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _02529_, _02500_);
  and (_02530_, _01909_, _42447_);
  and (_02531_, _01922_, _02267_);
  and (_02532_, _01926_, _02265_);
  or (_02533_, _02532_, _02531_);
  and (_02534_, _01931_, _02262_);
  and (_02535_, _01934_, _02260_);
  or (_02536_, _02535_, _02534_);
  or (_02537_, _02536_, _02533_);
  and (_02538_, _01946_, _02273_);
  and (_02539_, _01950_, _02271_);
  or (_02540_, _02539_, _02538_);
  and (_02541_, _01955_, _02276_);
  and (_02542_, _01960_, _02278_);
  or (_02543_, _02542_, _02541_);
  or (_02544_, _02543_, _02540_);
  or (_02545_, _02544_, _02537_);
  and (_02546_, _01968_, _02298_);
  and (_02547_, _01972_, _02296_);
  or (_02548_, _02547_, _02546_);
  and (_02549_, _01981_, _02291_);
  and (_02550_, _01978_, _02293_);
  or (_02551_, _02550_, _02549_);
  or (_02552_, _02551_, _02548_);
  and (_02553_, _01986_, _02283_);
  and (_02554_, _01992_, _02285_);
  and (_02555_, _01989_, _02287_);
  or (_02556_, _02555_, _02554_);
  or (_02557_, _02556_, _02553_);
  or (_02558_, _02557_, _02552_);
  or (_02559_, _02558_, _02545_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _02559_, _02530_);
  and (_02560_, _01909_, _42452_);
  and (_02561_, _01922_, _02332_);
  and (_02562_, _01926_, _02304_);
  or (_02563_, _02562_, _02561_);
  and (_02564_, _01931_, _02308_);
  and (_02565_, _01934_, _02306_);
  or (_02566_, _02565_, _02564_);
  or (_02567_, _02566_, _02563_);
  and (_02568_, _01946_, _02341_);
  and (_02569_, _01950_, _02343_);
  or (_02570_, _02569_, _02568_);
  and (_02571_, _01955_, _02339_);
  and (_02572_, _01960_, _02312_);
  or (_02573_, _02572_, _02571_);
  or (_02574_, _02573_, _02570_);
  or (_02575_, _02574_, _02567_);
  and (_02576_, _01968_, _02317_);
  and (_02577_, _01972_, _02325_);
  or (_02578_, _02577_, _02576_);
  and (_02579_, _01981_, _02321_);
  and (_02580_, _01978_, _02319_);
  or (_02581_, _02580_, _02579_);
  or (_02582_, _02581_, _02578_);
  and (_02583_, _01986_, _02334_);
  and (_02584_, _01992_, _02336_);
  and (_02585_, _01989_, _02327_);
  or (_02586_, _02585_, _02584_);
  or (_02587_, _02586_, _02583_);
  or (_02588_, _02587_, _02582_);
  or (_02589_, _02588_, _02575_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _02589_, _02560_);
  and (_02590_, _01909_, _42457_);
  and (_02591_, _01922_, _02377_);
  and (_02592_, _01926_, _02349_);
  or (_02593_, _02592_, _02591_);
  and (_02594_, _01931_, _02353_);
  and (_02595_, _01934_, _02351_);
  or (_02596_, _02595_, _02594_);
  or (_02597_, _02596_, _02593_);
  and (_02598_, _01946_, _02386_);
  and (_02599_, _01950_, _02388_);
  or (_02600_, _02599_, _02598_);
  and (_02601_, _01955_, _02357_);
  and (_02602_, _01960_, _02384_);
  or (_02603_, _02602_, _02601_);
  or (_02604_, _02603_, _02600_);
  or (_02605_, _02604_, _02597_);
  and (_02606_, _01972_, _02370_);
  and (_02607_, _01968_, _02362_);
  or (_02608_, _02607_, _02606_);
  and (_02609_, _01981_, _02366_);
  and (_02610_, _01978_, _02364_);
  or (_02611_, _02610_, _02609_);
  or (_02612_, _02611_, _02608_);
  and (_02613_, _01986_, _02379_);
  and (_02614_, _01992_, _02381_);
  and (_02615_, _01989_, _02372_);
  or (_02616_, _02615_, _02614_);
  or (_02617_, _02616_, _02613_);
  or (_02618_, _02617_, _02612_);
  or (_02619_, _02618_, _02605_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _02619_, _02590_);
  and (_02621_, _01909_, _42462_);
  and (_02622_, _01922_, _02422_);
  and (_02623_, _01926_, _02394_);
  or (_02624_, _02623_, _02622_);
  and (_02625_, _01931_, _02398_);
  and (_02626_, _01934_, _02396_);
  or (_02627_, _02626_, _02625_);
  or (_02628_, _02627_, _02624_);
  and (_02629_, _01946_, _02432_);
  and (_02630_, _01950_, _02434_);
  or (_02631_, _02630_, _02629_);
  and (_02632_, _01955_, _02402_);
  and (_02633_, _01960_, _02430_);
  or (_02634_, _02633_, _02632_);
  or (_02635_, _02634_, _02631_);
  or (_02636_, _02635_, _02628_);
  and (_02637_, _01972_, _02415_);
  and (_02638_, _01968_, _02407_);
  or (_02639_, _02638_, _02637_);
  and (_02640_, _01981_, _02411_);
  and (_02641_, _01978_, _02409_);
  or (_02642_, _02641_, _02640_);
  or (_02643_, _02642_, _02639_);
  and (_02644_, _01986_, _02424_);
  and (_02645_, _01992_, _02427_);
  and (_02646_, _01989_, _02417_);
  or (_02647_, _02646_, _02645_);
  or (_02648_, _02647_, _02644_);
  or (_02649_, _02648_, _02643_);
  or (_02650_, _02649_, _02636_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _02650_, _02621_);
  and (_02651_, _01992_, _42432_);
  and (_02652_, _01981_, _02156_);
  and (_02653_, _01978_, _02151_);
  and (_02654_, _01968_, _02154_);
  or (_02655_, _02654_, _02653_);
  or (_02656_, _02655_, _02652_);
  and (_02657_, _01955_, _02146_);
  and (_02658_, _01950_, _02144_);
  or (_02659_, _02658_, _02657_);
  and (_02660_, _01972_, _02141_);
  and (_02661_, _01960_, _02139_);
  or (_02662_, _02661_, _02660_);
  or (_02663_, _02662_, _02659_);
  or (_02664_, _02663_, _02656_);
  and (_02665_, _01946_, _02114_);
  and (_02666_, _01934_, _02111_);
  and (_02667_, _01931_, _02118_);
  and (_02668_, _01922_, _02121_);
  or (_02669_, _02668_, _02667_);
  or (_02670_, _02669_, _02666_);
  or (_02671_, _02670_, _02665_);
  and (_02672_, _01989_, _02134_);
  and (_02673_, _01986_, _02132_);
  or (_02674_, _02673_, _02672_);
  and (_02675_, _01926_, _02129_);
  and (_02676_, _01909_, _02126_);
  or (_02677_, _02676_, _02675_);
  or (_02678_, _02677_, _02674_);
  or (_02679_, _02678_, _02671_);
  or (_02680_, _02679_, _02664_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02680_, _02651_);
  and (_02681_, _01992_, _42437_);
  and (_02682_, _01989_, _02188_);
  or (_02683_, _02682_, _02681_);
  and (_02684_, _01986_, _02186_);
  and (_02685_, _01946_, _02166_);
  and (_02686_, _01934_, _02169_);
  and (_02687_, _01931_, _02173_);
  and (_02688_, _01922_, _02175_);
  or (_02689_, _02688_, _02687_);
  or (_02690_, _02689_, _02686_);
  or (_02691_, _02690_, _02685_);
  or (_02692_, _02691_, _02684_);
  or (_02693_, _02692_, _02683_);
  and (_02694_, _01968_, _02206_);
  and (_02695_, _01981_, _02208_);
  or (_02696_, _02695_, _02694_);
  and (_02697_, _01978_, _02204_);
  or (_02698_, _02697_, _02696_);
  and (_02699_, _01950_, _02200_);
  and (_02700_, _01955_, _02198_);
  or (_02701_, _02700_, _02699_);
  and (_02702_, _01960_, _02193_);
  and (_02703_, _01972_, _02195_);
  or (_02704_, _02703_, _02702_);
  or (_02705_, _02704_, _02701_);
  or (_02706_, _02705_, _02698_);
  and (_02707_, _01926_, _02183_);
  and (_02708_, _01909_, _02181_);
  or (_02709_, _02708_, _02707_);
  or (_02710_, _02709_, _02706_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02710_, _02693_);
  and (_02711_, _01986_, _02242_);
  and (_02712_, _01946_, _02249_);
  or (_02713_, _02712_, _02711_);
  and (_02714_, _01934_, _02222_);
  and (_02715_, _01922_, _02251_);
  and (_02716_, _01931_, _02253_);
  or (_02717_, _02716_, _02715_);
  or (_02718_, _02717_, _02714_);
  or (_02719_, _02718_, _02713_);
  and (_02720_, _01950_, _02235_);
  and (_02721_, _01981_, _02237_);
  and (_02722_, _01968_, _02246_);
  and (_02723_, _01978_, _02244_);
  or (_02724_, _02723_, _02722_);
  or (_02725_, _02724_, _02721_);
  or (_02726_, _02725_, _02720_);
  or (_02727_, _02726_, _02719_);
  and (_02728_, _01926_, _02216_);
  and (_02729_, _01989_, _02214_);
  and (_02730_, _01992_, _42442_);
  or (_02731_, _02730_, _02729_);
  or (_02732_, _02731_, _02728_);
  and (_02733_, _01909_, _02218_);
  and (_02734_, _01955_, _02227_);
  and (_02735_, _01960_, _02231_);
  and (_02736_, _01972_, _02229_);
  or (_02737_, _02736_, _02735_);
  or (_02738_, _02737_, _02734_);
  or (_02739_, _02738_, _02733_);
  or (_02740_, _02739_, _02732_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02740_, _02727_);
  and (_02741_, _01992_, _42447_);
  and (_02742_, _01989_, _02265_);
  and (_02743_, _01986_, _02267_);
  or (_02744_, _02743_, _02742_);
  and (_02745_, _01909_, _02262_);
  and (_02746_, _01926_, _02260_);
  or (_02747_, _02746_, _02745_);
  or (_02748_, _02747_, _02744_);
  and (_02749_, _01931_, _02271_);
  and (_02750_, _01922_, _02273_);
  or (_02751_, _02750_, _02749_);
  and (_02752_, _01934_, _02276_);
  and (_02753_, _01946_, _02278_);
  or (_02754_, _02753_, _02752_);
  or (_02755_, _02754_, _02751_);
  or (_02756_, _02755_, _02748_);
  and (_02757_, _01981_, _02287_);
  and (_02758_, _01968_, _02285_);
  and (_02759_, _01978_, _02283_);
  or (_02760_, _02759_, _02758_);
  or (_02761_, _02760_, _02757_);
  and (_02762_, _01972_, _02293_);
  and (_02763_, _01960_, _02291_);
  or (_02764_, _02763_, _02762_);
  and (_02765_, _01950_, _02296_);
  and (_02766_, _01955_, _02298_);
  or (_02767_, _02766_, _02765_);
  or (_02768_, _02767_, _02764_);
  or (_02769_, _02768_, _02761_);
  or (_02770_, _02769_, _02756_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02770_, _02741_);
  and (_02771_, _01992_, _42452_);
  and (_02772_, _01981_, _02327_);
  and (_02773_, _01968_, _02336_);
  and (_02774_, _01978_, _02334_);
  or (_02775_, _02774_, _02773_);
  or (_02776_, _02775_, _02772_);
  and (_02777_, _01972_, _02319_);
  and (_02778_, _01960_, _02321_);
  or (_02779_, _02778_, _02777_);
  and (_02780_, _01950_, _02325_);
  and (_02781_, _01955_, _02317_);
  or (_02782_, _02781_, _02780_);
  or (_02783_, _02782_, _02779_);
  or (_02784_, _02783_, _02776_);
  and (_02785_, _01946_, _02312_);
  and (_02786_, _01934_, _02339_);
  and (_02787_, _01931_, _02343_);
  and (_02788_, _01922_, _02341_);
  or (_02789_, _02788_, _02787_);
  or (_02790_, _02789_, _02786_);
  or (_02791_, _02790_, _02785_);
  and (_02792_, _01989_, _02304_);
  and (_02793_, _01986_, _02332_);
  or (_02794_, _02793_, _02792_);
  and (_02795_, _01926_, _02306_);
  and (_02796_, _01909_, _02308_);
  or (_02797_, _02796_, _02795_);
  or (_02798_, _02797_, _02794_);
  or (_02799_, _02798_, _02791_);
  or (_02800_, _02799_, _02784_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02800_, _02771_);
  and (_02801_, _01992_, _42457_);
  and (_02802_, _01989_, _02349_);
  and (_02803_, _01986_, _02377_);
  or (_02804_, _02803_, _02802_);
  and (_02805_, _01926_, _02351_);
  and (_02806_, _01909_, _02353_);
  or (_02807_, _02806_, _02805_);
  or (_02808_, _02807_, _02804_);
  and (_02809_, _01922_, _02386_);
  and (_02810_, _01931_, _02388_);
  or (_02811_, _02810_, _02809_);
  and (_02812_, _01946_, _02384_);
  and (_02813_, _01934_, _02357_);
  or (_02815_, _02813_, _02812_);
  or (_02816_, _02815_, _02811_);
  or (_02817_, _02816_, _02808_);
  and (_02818_, _01981_, _02372_);
  and (_02819_, _01968_, _02381_);
  and (_02820_, _01978_, _02379_);
  or (_02821_, _02820_, _02819_);
  or (_02822_, _02821_, _02818_);
  and (_02823_, _01972_, _02364_);
  and (_02824_, _01960_, _02366_);
  or (_02825_, _02824_, _02823_);
  and (_02826_, _01950_, _02370_);
  and (_02827_, _01955_, _02362_);
  or (_02828_, _02827_, _02826_);
  or (_02829_, _02828_, _02825_);
  or (_02830_, _02829_, _02822_);
  or (_02831_, _02830_, _02817_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02831_, _02801_);
  and (_02832_, _01992_, _42462_);
  and (_02833_, _01989_, _02394_);
  and (_02834_, _01986_, _02422_);
  or (_02835_, _02834_, _02833_);
  and (_02836_, _01926_, _02396_);
  and (_02837_, _01909_, _02398_);
  or (_02838_, _02837_, _02836_);
  or (_02839_, _02838_, _02835_);
  and (_02840_, _01931_, _02434_);
  and (_02841_, _01922_, _02432_);
  or (_02842_, _02841_, _02840_);
  and (_02843_, _01946_, _02430_);
  and (_02844_, _01934_, _02402_);
  or (_02845_, _02844_, _02843_);
  or (_02846_, _02845_, _02842_);
  or (_02847_, _02846_, _02839_);
  and (_02848_, _01981_, _02417_);
  and (_02849_, _01968_, _02427_);
  and (_02850_, _01978_, _02424_);
  or (_02851_, _02850_, _02849_);
  or (_02852_, _02851_, _02848_);
  and (_02853_, _01972_, _02409_);
  and (_02854_, _01960_, _02411_);
  or (_02855_, _02854_, _02853_);
  and (_02856_, _01955_, _02407_);
  and (_02857_, _01950_, _02415_);
  or (_02858_, _02857_, _02856_);
  or (_02859_, _02858_, _02855_);
  or (_02860_, _02859_, _02852_);
  or (_02861_, _02860_, _02847_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02861_, _02832_);
  and (_02862_, _01986_, _42432_);
  and (_02863_, _01950_, _02111_);
  and (_02864_, _01955_, _02114_);
  or (_02865_, _02864_, _02863_);
  and (_02866_, _01946_, _02118_);
  and (_02867_, _01934_, _02121_);
  or (_02868_, _02867_, _02866_);
  or (_02869_, _02868_, _02865_);
  and (_02870_, _01931_, _02129_);
  and (_02871_, _01922_, _02126_);
  or (_02872_, _02871_, _02870_);
  and (_02873_, _01926_, _02132_);
  and (_02874_, _01909_, _02134_);
  or (_02875_, _02874_, _02873_);
  or (_02876_, _02875_, _02872_);
  or (_02877_, _02876_, _02869_);
  and (_02878_, _01960_, _02144_);
  and (_02879_, _01972_, _02146_);
  or (_02880_, _02879_, _02878_);
  and (_02881_, _01968_, _02139_);
  and (_02882_, _01981_, _02141_);
  or (_02883_, _02882_, _02881_);
  or (_02884_, _02883_, _02880_);
  and (_02885_, _01989_, _02151_);
  and (_02886_, _01992_, _02156_);
  and (_02887_, _01978_, _02154_);
  or (_02888_, _02887_, _02886_);
  or (_02889_, _02888_, _02885_);
  or (_02890_, _02889_, _02884_);
  or (_02891_, _02890_, _02877_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _02891_, _02862_);
  and (_02892_, _01986_, _42437_);
  and (_02893_, _01931_, _02183_);
  and (_02894_, _01922_, _02181_);
  or (_02895_, _02894_, _02893_);
  and (_02896_, _01926_, _02186_);
  and (_02897_, _01909_, _02188_);
  or (_02898_, _02897_, _02896_);
  or (_02899_, _02898_, _02895_);
  and (_02900_, _01946_, _02173_);
  and (_02901_, _01934_, _02175_);
  or (_02902_, _02901_, _02900_);
  and (_02903_, _01950_, _02169_);
  and (_02904_, _01955_, _02166_);
  or (_02905_, _02904_, _02903_);
  or (_02906_, _02905_, _02902_);
  or (_02907_, _02906_, _02899_);
  and (_02908_, _01960_, _02200_);
  and (_02909_, _01972_, _02198_);
  or (_02910_, _02909_, _02908_);
  and (_02911_, _01968_, _02193_);
  and (_02912_, _01981_, _02195_);
  or (_02913_, _02912_, _02911_);
  or (_02914_, _02913_, _02910_);
  and (_02915_, _01989_, _02204_);
  and (_02916_, _01992_, _02208_);
  and (_02917_, _01978_, _02206_);
  or (_02918_, _02917_, _02916_);
  or (_02919_, _02918_, _02915_);
  or (_02920_, _02919_, _02914_);
  or (_02921_, _02920_, _02907_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _02921_, _02892_);
  and (_02922_, _01986_, _42442_);
  and (_02923_, _01972_, _02227_);
  and (_02924_, _01960_, _02235_);
  or (_02925_, _02924_, _02923_);
  and (_02926_, _01968_, _02231_);
  and (_02927_, _01981_, _02229_);
  or (_02928_, _02927_, _02926_);
  or (_02929_, _02928_, _02925_);
  and (_02930_, _01989_, _02244_);
  and (_02931_, _01978_, _02246_);
  and (_02932_, _01992_, _02237_);
  or (_02933_, _02932_, _02931_);
  or (_02934_, _02933_, _02930_);
  or (_02935_, _02934_, _02929_);
  and (_02936_, _01946_, _02253_);
  and (_02937_, _01934_, _02251_);
  or (_02938_, _02937_, _02936_);
  and (_02939_, _01955_, _02249_);
  and (_02940_, _01950_, _02222_);
  or (_02941_, _02940_, _02939_);
  or (_02942_, _02941_, _02938_);
  and (_02943_, _01931_, _02216_);
  and (_02944_, _01922_, _02218_);
  or (_02945_, _02944_, _02943_);
  and (_02946_, _01926_, _02242_);
  and (_02947_, _01909_, _02214_);
  or (_02948_, _02947_, _02946_);
  or (_02949_, _02948_, _02945_);
  or (_02950_, _02949_, _02942_);
  or (_02951_, _02950_, _02935_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _02951_, _02922_);
  and (_02952_, _01986_, _42447_);
  and (_02953_, _01972_, _02298_);
  and (_02954_, _01960_, _02296_);
  or (_02955_, _02954_, _02953_);
  and (_02956_, _01981_, _02293_);
  and (_02957_, _01968_, _02291_);
  or (_02958_, _02957_, _02956_);
  or (_02959_, _02958_, _02955_);
  and (_02960_, _01989_, _02283_);
  and (_02961_, _01978_, _02285_);
  and (_02962_, _01992_, _02287_);
  or (_02963_, _02962_, _02961_);
  or (_02964_, _02963_, _02960_);
  or (_02965_, _02964_, _02959_);
  and (_02966_, _01931_, _02260_);
  and (_02967_, _01922_, _02262_);
  or (_02968_, _02967_, _02966_);
  and (_02969_, _01909_, _02265_);
  and (_02971_, _01926_, _02267_);
  or (_02972_, _02971_, _02969_);
  or (_02973_, _02972_, _02968_);
  and (_02974_, _01946_, _02271_);
  and (_02975_, _01934_, _02273_);
  or (_02976_, _02975_, _02974_);
  and (_02977_, _01955_, _02278_);
  and (_02978_, _01950_, _02276_);
  or (_02979_, _02978_, _02977_);
  or (_02980_, _02979_, _02976_);
  or (_02982_, _02980_, _02973_);
  or (_02983_, _02982_, _02965_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02983_, _02952_);
  and (_02984_, _01986_, _42452_);
  and (_02985_, _01931_, _02306_);
  and (_02986_, _01922_, _02308_);
  or (_02987_, _02986_, _02985_);
  and (_02988_, _01926_, _02332_);
  and (_02989_, _01909_, _02304_);
  or (_02990_, _02989_, _02988_);
  or (_02991_, _02990_, _02987_);
  and (_02992_, _01946_, _02343_);
  and (_02993_, _01934_, _02341_);
  or (_02994_, _02993_, _02992_);
  and (_02995_, _01950_, _02339_);
  and (_02996_, _01955_, _02312_);
  or (_02997_, _02996_, _02995_);
  or (_02998_, _02997_, _02994_);
  or (_02999_, _02998_, _02991_);
  and (_03000_, _01960_, _02325_);
  and (_03002_, _01972_, _02317_);
  or (_03003_, _03002_, _03000_);
  and (_03004_, _01968_, _02321_);
  and (_03005_, _01981_, _02319_);
  or (_03006_, _03005_, _03004_);
  or (_03007_, _03006_, _03003_);
  and (_03008_, _01989_, _02334_);
  and (_03009_, _01992_, _02327_);
  and (_03010_, _01978_, _02336_);
  or (_03011_, _03010_, _03009_);
  or (_03013_, _03011_, _03008_);
  or (_03014_, _03013_, _03007_);
  or (_03015_, _03014_, _02999_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _03015_, _02984_);
  and (_03016_, _01986_, _42457_);
  and (_03017_, _01931_, _02351_);
  and (_03018_, _01922_, _02353_);
  or (_03019_, _03018_, _03017_);
  and (_03020_, _01926_, _02377_);
  and (_03021_, _01909_, _02349_);
  or (_03023_, _03021_, _03020_);
  or (_03024_, _03023_, _03019_);
  and (_03025_, _01946_, _02388_);
  and (_03026_, _01934_, _02386_);
  or (_03027_, _03026_, _03025_);
  and (_03028_, _01955_, _02384_);
  and (_03029_, _01950_, _02357_);
  or (_03030_, _03029_, _03028_);
  or (_03031_, _03030_, _03027_);
  or (_03032_, _03031_, _03024_);
  and (_03033_, _01960_, _02370_);
  and (_03034_, _01972_, _02362_);
  or (_03035_, _03034_, _03033_);
  and (_03036_, _01981_, _02364_);
  and (_03037_, _01968_, _02366_);
  or (_03038_, _03037_, _03036_);
  or (_03039_, _03038_, _03035_);
  and (_03040_, _01989_, _02379_);
  and (_03041_, _01992_, _02372_);
  and (_03042_, _01978_, _02381_);
  or (_03044_, _03042_, _03041_);
  or (_03045_, _03044_, _03040_);
  or (_03046_, _03045_, _03039_);
  or (_03047_, _03046_, _03032_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _03047_, _03016_);
  and (_03048_, _01986_, _42462_);
  and (_03049_, _01931_, _02396_);
  and (_03050_, _01922_, _02398_);
  or (_03051_, _03050_, _03049_);
  and (_03052_, _01926_, _02422_);
  and (_03054_, _01909_, _02394_);
  or (_03055_, _03054_, _03052_);
  or (_03056_, _03055_, _03051_);
  and (_03057_, _01946_, _02434_);
  and (_03058_, _01934_, _02432_);
  or (_03059_, _03058_, _03057_);
  and (_03060_, _01955_, _02430_);
  and (_03061_, _01950_, _02402_);
  or (_03062_, _03061_, _03060_);
  or (_03063_, _03062_, _03059_);
  or (_03065_, _03063_, _03056_);
  and (_03066_, _01960_, _02415_);
  and (_03067_, _01972_, _02407_);
  or (_03068_, _03067_, _03066_);
  and (_03069_, _01981_, _02409_);
  and (_03070_, _01968_, _02411_);
  or (_03071_, _03070_, _03069_);
  or (_03072_, _03071_, _03068_);
  and (_03073_, _01989_, _02424_);
  and (_03074_, _01992_, _02417_);
  and (_03076_, _01978_, _02427_);
  or (_03077_, _03076_, _03074_);
  or (_03078_, _03077_, _03073_);
  or (_03079_, _03078_, _03072_);
  or (_03080_, _03079_, _03065_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _03080_, _03048_);
  nand (_03081_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_03082_, \oc8051_golden_model_1.PC [3]);
  or (_03083_, \oc8051_golden_model_1.PC [2], _03082_);
  or (_03084_, _03083_, _03081_);
  or (_03086_, _03084_, _42298_);
  not (_03087_, \oc8051_golden_model_1.PC [1]);
  or (_03088_, _03087_, \oc8051_golden_model_1.PC [0]);
  or (_03089_, _03088_, _03083_);
  or (_03090_, _03089_, _42257_);
  and (_03091_, _03090_, _03086_);
  not (_03092_, \oc8051_golden_model_1.PC [2]);
  or (_03093_, _03092_, \oc8051_golden_model_1.PC [3]);
  or (_03094_, _03093_, _03081_);
  or (_03095_, _03094_, _42134_);
  or (_03097_, _03093_, _03088_);
  or (_03098_, _03097_, _42093_);
  and (_03099_, _03098_, _03095_);
  and (_03100_, _03099_, _03091_);
  and (_03101_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  and (_03102_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and (_03103_, _03102_, _03101_);
  nand (_03104_, _03103_, _42462_);
  nand (_03105_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_03106_, _03105_, _03088_);
  or (_03108_, _03106_, _42421_);
  and (_03109_, _03108_, _03104_);
  or (_03110_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_03111_, _03110_, _03081_);
  or (_03112_, _03111_, _41970_);
  or (_03113_, _03110_, _03088_);
  or (_03114_, _03113_, _41929_);
  and (_03115_, _03114_, _03112_);
  and (_03116_, _03115_, _03109_);
  and (_03117_, _03116_, _03100_);
  not (_03119_, \oc8051_golden_model_1.PC [0]);
  or (_03120_, \oc8051_golden_model_1.PC [1], _03119_);
  or (_03121_, _03120_, _03105_);
  or (_03122_, _03121_, _42380_);
  or (_03123_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_03124_, _03123_, _03105_);
  or (_03125_, _03124_, _42339_);
  and (_03126_, _03125_, _03122_);
  or (_03127_, _03110_, _03123_);
  or (_03128_, _03127_, _41832_);
  or (_03130_, _03110_, _03120_);
  or (_03131_, _03130_, _41880_);
  and (_03132_, _03131_, _03128_);
  and (_03133_, _03132_, _03126_);
  or (_03134_, _03120_, _03083_);
  or (_03135_, _03134_, _42216_);
  or (_03136_, _03123_, _03083_);
  or (_03137_, _03136_, _42175_);
  and (_03138_, _03137_, _03135_);
  or (_03139_, _03120_, _03093_);
  or (_03140_, _03139_, _42052_);
  or (_03141_, _03123_, _03093_);
  or (_03142_, _03141_, _42011_);
  and (_03143_, _03142_, _03140_);
  and (_03144_, _03143_, _03138_);
  and (_03145_, _03144_, _03133_);
  and (_03146_, _03145_, _03117_);
  or (_03147_, _03084_, _42263_);
  or (_03148_, _03089_, _42222_);
  and (_03149_, _03148_, _03147_);
  or (_03150_, _03094_, _42099_);
  or (_03151_, _03097_, _42058_);
  and (_03152_, _03151_, _03150_);
  and (_03153_, _03152_, _03149_);
  nand (_03154_, _03103_, _42427_);
  or (_03155_, _03106_, _42386_);
  and (_03156_, _03155_, _03154_);
  or (_03157_, _03111_, _41935_);
  or (_03158_, _03113_, _41893_);
  and (_03159_, _03158_, _03157_);
  and (_03160_, _03159_, _03156_);
  and (_03161_, _03160_, _03153_);
  or (_03162_, _03121_, _42345_);
  or (_03163_, _03124_, _42304_);
  and (_03164_, _03163_, _03162_);
  or (_03165_, _03127_, _41797_);
  or (_03166_, _03130_, _41840_);
  and (_03167_, _03166_, _03165_);
  and (_03168_, _03167_, _03164_);
  or (_03169_, _03134_, _42181_);
  or (_03170_, _03136_, _42140_);
  and (_03171_, _03170_, _03169_);
  or (_03172_, _03139_, _42017_);
  or (_03173_, _03141_, _41976_);
  and (_03174_, _03173_, _03172_);
  and (_03175_, _03174_, _03171_);
  and (_03176_, _03175_, _03168_);
  and (_03177_, _03176_, _03161_);
  and (_03178_, _03177_, _03146_);
  or (_03179_, _03084_, _42288_);
  or (_03180_, _03089_, _42247_);
  and (_03181_, _03180_, _03179_);
  or (_03182_, _03094_, _42124_);
  or (_03183_, _03097_, _42083_);
  and (_03184_, _03183_, _03182_);
  and (_03185_, _03184_, _03181_);
  nand (_03186_, _03103_, _42452_);
  or (_03187_, _03106_, _42411_);
  and (_03188_, _03187_, _03186_);
  or (_03189_, _03111_, _41960_);
  or (_03190_, _03113_, _41919_);
  and (_03191_, _03190_, _03189_);
  and (_03192_, _03191_, _03188_);
  and (_03193_, _03192_, _03185_);
  or (_03194_, _03121_, _42370_);
  or (_03195_, _03124_, _42329_);
  and (_03196_, _03195_, _03194_);
  or (_03197_, _03127_, _41822_);
  or (_03198_, _03130_, _41870_);
  and (_03199_, _03198_, _03197_);
  and (_03200_, _03199_, _03196_);
  or (_03201_, _03134_, _42206_);
  or (_03202_, _03136_, _42165_);
  and (_03203_, _03202_, _03201_);
  or (_03204_, _03139_, _42042_);
  or (_03205_, _03141_, _42001_);
  and (_03206_, _03205_, _03204_);
  and (_03207_, _03206_, _03203_);
  and (_03208_, _03207_, _03200_);
  and (_03209_, _03208_, _03193_);
  or (_03210_, _03084_, _42293_);
  or (_03211_, _03089_, _42252_);
  and (_03212_, _03211_, _03210_);
  or (_03213_, _03094_, _42129_);
  or (_03214_, _03097_, _42088_);
  and (_03215_, _03214_, _03213_);
  and (_03216_, _03215_, _03212_);
  nand (_03217_, _03103_, _42457_);
  or (_03218_, _03106_, _42416_);
  and (_03219_, _03218_, _03217_);
  or (_03221_, _03111_, _41965_);
  or (_03222_, _03113_, _41924_);
  and (_03223_, _03222_, _03221_);
  and (_03224_, _03223_, _03219_);
  and (_03225_, _03224_, _03216_);
  or (_03226_, _03121_, _42375_);
  or (_03227_, _03124_, _42334_);
  and (_03228_, _03227_, _03226_);
  or (_03229_, _03127_, _41827_);
  or (_03230_, _03130_, _41875_);
  and (_03231_, _03230_, _03229_);
  and (_03232_, _03231_, _03228_);
  or (_03233_, _03134_, _42211_);
  or (_03234_, _03136_, _42170_);
  and (_03235_, _03234_, _03233_);
  or (_03236_, _03139_, _42047_);
  or (_03237_, _03141_, _42006_);
  and (_03238_, _03237_, _03236_);
  and (_03239_, _03238_, _03235_);
  and (_03240_, _03239_, _03232_);
  nand (_03241_, _03240_, _03225_);
  or (_03242_, _03241_, _03209_);
  not (_03243_, _03242_);
  and (_03244_, _03243_, _03178_);
  or (_03245_, _03084_, _42268_);
  or (_03246_, _03089_, _42227_);
  and (_03247_, _03246_, _03245_);
  or (_03248_, _03094_, _42104_);
  or (_03249_, _03097_, _42063_);
  and (_03250_, _03249_, _03248_);
  and (_03251_, _03250_, _03247_);
  nand (_03252_, _03103_, _42432_);
  or (_03253_, _03106_, _42391_);
  and (_03254_, _03253_, _03252_);
  or (_03255_, _03111_, _41940_);
  or (_03256_, _03113_, _41899_);
  and (_03257_, _03256_, _03255_);
  and (_03258_, _03257_, _03254_);
  and (_03259_, _03258_, _03251_);
  or (_03260_, _03121_, _42350_);
  or (_03261_, _03124_, _42309_);
  and (_03262_, _03261_, _03260_);
  or (_03263_, _03127_, _41802_);
  or (_03264_, _03130_, _41850_);
  and (_03265_, _03264_, _03263_);
  and (_03266_, _03265_, _03262_);
  or (_03267_, _03134_, _42186_);
  or (_03268_, _03136_, _42145_);
  and (_03269_, _03268_, _03267_);
  or (_03270_, _03139_, _42022_);
  or (_03271_, _03141_, _41981_);
  and (_03272_, _03271_, _03270_);
  and (_03273_, _03272_, _03269_);
  and (_03274_, _03273_, _03266_);
  and (_03275_, _03274_, _03259_);
  or (_03276_, _03084_, _42273_);
  or (_03277_, _03089_, _42232_);
  and (_03278_, _03277_, _03276_);
  or (_03279_, _03094_, _42109_);
  or (_03280_, _03097_, _42068_);
  and (_03281_, _03280_, _03279_);
  and (_03282_, _03281_, _03278_);
  nand (_03283_, _03103_, _42437_);
  or (_03284_, _03106_, _42396_);
  and (_03285_, _03284_, _03283_);
  or (_03286_, _03111_, _41945_);
  or (_03287_, _03113_, _41904_);
  and (_03288_, _03287_, _03286_);
  and (_03289_, _03288_, _03285_);
  and (_03290_, _03289_, _03282_);
  or (_03291_, _03121_, _42355_);
  or (_03292_, _03124_, _42314_);
  and (_03293_, _03292_, _03291_);
  or (_03294_, _03127_, _41807_);
  or (_03295_, _03130_, _41855_);
  and (_03296_, _03295_, _03294_);
  and (_03297_, _03296_, _03293_);
  or (_03298_, _03134_, _42191_);
  or (_03299_, _03136_, _42150_);
  and (_03300_, _03299_, _03298_);
  or (_03301_, _03139_, _42027_);
  or (_03302_, _03141_, _41986_);
  and (_03303_, _03302_, _03301_);
  and (_03304_, _03303_, _03300_);
  and (_03305_, _03304_, _03297_);
  nand (_03306_, _03305_, _03290_);
  not (_03307_, _03306_);
  and (_03308_, _03307_, _03275_);
  or (_03309_, _03084_, _42278_);
  or (_03310_, _03089_, _42237_);
  and (_03311_, _03310_, _03309_);
  or (_03312_, _03094_, _42114_);
  or (_03313_, _03097_, _42073_);
  and (_03314_, _03313_, _03312_);
  and (_03315_, _03314_, _03311_);
  nand (_03316_, _03103_, _42442_);
  or (_03317_, _03106_, _42401_);
  and (_03318_, _03317_, _03316_);
  or (_03319_, _03111_, _41950_);
  or (_03320_, _03113_, _41909_);
  and (_03321_, _03320_, _03319_);
  and (_03322_, _03321_, _03318_);
  and (_03323_, _03322_, _03315_);
  or (_03324_, _03121_, _42360_);
  or (_03325_, _03124_, _42319_);
  and (_03326_, _03325_, _03324_);
  or (_03327_, _03127_, _41812_);
  or (_03328_, _03130_, _41860_);
  and (_03329_, _03328_, _03327_);
  and (_03330_, _03329_, _03326_);
  or (_03331_, _03134_, _42196_);
  or (_03332_, _03136_, _42155_);
  and (_03333_, _03332_, _03331_);
  or (_03334_, _03139_, _42032_);
  or (_03335_, _03141_, _41991_);
  and (_03336_, _03335_, _03334_);
  and (_03337_, _03336_, _03333_);
  and (_03338_, _03337_, _03330_);
  nand (_03339_, _03338_, _03323_);
  or (_03340_, _03084_, _42283_);
  or (_03341_, _03089_, _42242_);
  and (_03342_, _03341_, _03340_);
  or (_03343_, _03094_, _42119_);
  or (_03344_, _03097_, _42078_);
  and (_03345_, _03344_, _03343_);
  and (_03346_, _03345_, _03342_);
  nand (_03347_, _03103_, _42447_);
  or (_03348_, _03106_, _42406_);
  and (_03349_, _03348_, _03347_);
  or (_03350_, _03111_, _41955_);
  or (_03351_, _03113_, _41914_);
  and (_03352_, _03351_, _03350_);
  and (_03353_, _03352_, _03349_);
  and (_03354_, _03353_, _03346_);
  or (_03355_, _03121_, _42365_);
  or (_03356_, _03124_, _42324_);
  and (_03357_, _03356_, _03355_);
  or (_03358_, _03127_, _41817_);
  or (_03359_, _03130_, _41865_);
  and (_03360_, _03359_, _03358_);
  and (_03361_, _03360_, _03357_);
  or (_03362_, _03134_, _42201_);
  or (_03363_, _03136_, _42160_);
  and (_03364_, _03363_, _03362_);
  or (_03365_, _03139_, _42037_);
  or (_03366_, _03141_, _41996_);
  and (_03367_, _03366_, _03365_);
  and (_03368_, _03367_, _03364_);
  and (_03369_, _03368_, _03361_);
  nand (_03370_, _03369_, _03354_);
  or (_03371_, _03370_, _03339_);
  not (_03372_, _03371_);
  and (_03373_, _03372_, _03308_);
  and (_03374_, _03373_, _03244_);
  not (_03375_, _03374_);
  or (_03376_, _03306_, _03275_);
  or (_03377_, _03376_, _03371_);
  not (_03378_, _03377_);
  and (_03379_, _03240_, _03225_);
  or (_03380_, _03379_, _03209_);
  not (_03381_, _03380_);
  and (_03382_, _03381_, _03178_);
  and (_03383_, _03382_, _03378_);
  not (_03384_, _03383_);
  nand (_03385_, _03145_, _03117_);
  and (_03386_, _03177_, _03385_);
  and (_03387_, _03386_, _03243_);
  and (_03388_, _03387_, _03378_);
  nand (_03389_, _03208_, _03193_);
  or (_03390_, _03241_, _03389_);
  not (_03391_, _03390_);
  and (_03392_, _03391_, _03386_);
  and (_03393_, _03392_, _03378_);
  nor (_03394_, _03393_, _03388_);
  and (_03395_, _03394_, _03384_);
  or (_03396_, _03177_, _03385_);
  nor (_03397_, _03396_, _03390_);
  and (_03398_, _03397_, _03378_);
  not (_03399_, _03398_);
  and (_03400_, _03386_, _03381_);
  and (_03401_, _03400_, _03378_);
  or (_03402_, _03379_, _03389_);
  not (_03403_, _03402_);
  and (_03404_, _03403_, _03386_);
  and (_03405_, _03404_, _03378_);
  nor (_03406_, _03405_, _03401_);
  and (_03407_, _03406_, _03399_);
  and (_03408_, _03407_, _03395_);
  and (_03409_, _03403_, _03178_);
  and (_03410_, _03409_, _03378_);
  not (_03411_, _03410_);
  and (_03412_, _03391_, _03178_);
  and (_03413_, _03412_, _03378_);
  and (_03414_, _03378_, _03244_);
  nor (_03415_, _03414_, _03413_);
  and (_03416_, _03415_, _03411_);
  and (_03417_, _03416_, _03408_);
  nor (_03418_, _03417_, _03087_);
  not (_03419_, _03418_);
  not (_03420_, _03275_);
  and (_03422_, _03306_, _03420_);
  and (_03423_, _03422_, _03372_);
  nor (_03424_, _03396_, _03242_);
  and (_03425_, _03424_, _03423_);
  not (_03426_, _03425_);
  or (_03427_, _03396_, _03380_);
  or (_03428_, _03427_, _03377_);
  or (_03429_, _03177_, _03146_);
  or (_03430_, _03429_, _03242_);
  or (_03431_, _03430_, _03377_);
  and (_03432_, _03431_, _03428_);
  or (_03433_, _03429_, _03390_);
  or (_03434_, _03433_, _03377_);
  or (_03435_, _03429_, _03402_);
  or (_03436_, _03435_, _03377_);
  and (_03437_, _03436_, _03434_);
  or (_03438_, _03429_, _03380_);
  or (_03439_, _03438_, _03377_);
  or (_03440_, _03396_, _03402_);
  or (_03441_, _03440_, _03377_);
  and (_03442_, _03441_, _03439_);
  and (_03443_, _03442_, _03437_);
  and (_03444_, _03443_, _03432_);
  or (_03445_, _03444_, \oc8051_golden_model_1.PC [1]);
  nand (_03446_, _03443_, _03432_);
  nand (_03447_, _03123_, _03081_);
  or (_03448_, _03447_, _03446_);
  nand (_03449_, _03448_, _03445_);
  nand (_03450_, _03449_, _03426_);
  not (_03451_, _03376_);
  not (_03452_, _03370_);
  and (_03453_, _03452_, _03339_);
  and (_03454_, _03453_, _03451_);
  and (_03455_, _03454_, _03397_);
  and (_03456_, _03424_, _03378_);
  nor (_03457_, _03456_, _03455_);
  not (_03458_, _03457_);
  and (_03459_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  and (_03460_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_03461_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_03462_, _03461_, _03460_);
  and (_03463_, _03462_, _03459_);
  nor (_03464_, _03462_, _03459_);
  nor (_03465_, _03464_, _03463_);
  and (_03466_, _03465_, _03425_);
  nor (_03467_, _03466_, _03458_);
  nand (_03468_, _03467_, _03450_);
  and (_03469_, _03423_, _03397_);
  nor (_03470_, _03457_, _03087_);
  nor (_03471_, _03470_, _03469_);
  nand (_03472_, _03471_, _03468_);
  and (_03473_, \oc8051_golden_model_1.ACC [0], _03119_);
  not (_03474_, \oc8051_golden_model_1.ACC [1]);
  nor (_03475_, _03447_, _03474_);
  and (_03476_, _03447_, _03474_);
  nor (_03477_, _03476_, _03475_);
  and (_03478_, _03477_, _03473_);
  not (_03479_, _03469_);
  nor (_03480_, _03477_, _03473_);
  or (_03481_, _03480_, _03479_);
  or (_03482_, _03481_, _03478_);
  and (_03483_, _03482_, _03417_);
  nand (_03484_, _03483_, _03472_);
  and (_03485_, _03484_, _03419_);
  or (_03486_, _03444_, _03119_);
  or (_03487_, _03446_, \oc8051_golden_model_1.PC [0]);
  nand (_03488_, _03487_, _03486_);
  and (_03489_, _03488_, _03426_);
  nor (_03490_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03491_, _03490_, _03459_);
  and (_03492_, _03491_, _03425_);
  or (_03493_, _03492_, _03458_);
  or (_03494_, _03493_, _03489_);
  nor (_03495_, _03457_, \oc8051_golden_model_1.PC [0]);
  nor (_03496_, _03495_, _03469_);
  nand (_03497_, _03496_, _03494_);
  not (_03498_, \oc8051_golden_model_1.ACC [0]);
  and (_03499_, _03498_, \oc8051_golden_model_1.PC [0]);
  or (_03500_, _03473_, _03479_);
  or (_03501_, _03500_, _03499_);
  and (_03502_, _03501_, _03417_);
  nand (_03503_, _03502_, _03497_);
  nor (_03504_, _03417_, \oc8051_golden_model_1.PC [0]);
  not (_03505_, _03504_);
  and (_03506_, _03505_, _03503_);
  and (_03507_, _03506_, _03485_);
  and (_03508_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03509_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03510_, _03509_, _03508_);
  not (_03511_, _03510_);
  nor (_03512_, _03511_, _03416_);
  not (_03513_, _03512_);
  or (_03514_, _03458_, _03446_);
  and (_03515_, _03514_, _03511_);
  and (_03516_, _03101_, \oc8051_golden_model_1.PC [2]);
  and (_03517_, _03081_, _03092_);
  nor (_03518_, _03517_, _03516_);
  nor (_03519_, _03518_, _03425_);
  and (_03520_, _03519_, _03444_);
  nor (_03521_, _03463_, _03460_);
  and (_03522_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_03523_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_03524_, _03523_, _03522_);
  not (_03525_, _03524_);
  nor (_03526_, _03525_, _03521_);
  and (_03527_, _03525_, _03521_);
  nor (_03528_, _03527_, _03526_);
  not (_03529_, _03528_);
  and (_03530_, _03529_, _03425_);
  or (_03531_, _03530_, _03520_);
  and (_03532_, _03531_, _03457_);
  or (_03533_, _03532_, _03469_);
  or (_03534_, _03533_, _03515_);
  nor (_03535_, _03478_, _03475_);
  and (_03536_, _03518_, \oc8051_golden_model_1.ACC [2]);
  nor (_03537_, _03518_, \oc8051_golden_model_1.ACC [2]);
  nor (_03538_, _03537_, _03536_);
  not (_03539_, _03538_);
  nor (_03540_, _03539_, _03535_);
  and (_03541_, _03539_, _03535_);
  nor (_03542_, _03541_, _03540_);
  and (_03543_, _03542_, _03469_);
  not (_03544_, _03543_);
  and (_03545_, _03544_, _03408_);
  nand (_03546_, _03545_, _03534_);
  or (_03547_, _03510_, _03417_);
  nand (_03548_, _03547_, _03546_);
  nand (_03549_, _03548_, _03513_);
  and (_03550_, _03102_, \oc8051_golden_model_1.PC [1]);
  nor (_03551_, _03508_, \oc8051_golden_model_1.PC [3]);
  nor (_03552_, _03551_, _03550_);
  nor (_03553_, _03552_, _03417_);
  not (_03554_, _03553_);
  nor (_03555_, _03552_, _03457_);
  not (_03556_, _03094_);
  nor (_03557_, _03516_, _03082_);
  nor (_03558_, _03557_, _03556_);
  not (_03559_, _03558_);
  or (_03560_, _03446_, _03559_);
  or (_03561_, _03552_, _03444_);
  and (_03562_, _03561_, _03560_);
  nand (_03563_, _03562_, _03426_);
  nor (_03564_, _03526_, _03522_);
  and (_03565_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03566_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03567_, _03566_, _03565_);
  not (_03568_, _03567_);
  nor (_03569_, _03568_, _03564_);
  and (_03570_, _03568_, _03564_);
  nor (_03571_, _03570_, _03569_);
  nand (_03572_, _03571_, _03425_);
  and (_03573_, _03572_, _03457_);
  nand (_03574_, _03573_, _03563_);
  nand (_03575_, _03574_, _03479_);
  or (_03576_, _03575_, _03555_);
  nor (_03577_, _03540_, _03536_);
  nor (_03578_, _03558_, \oc8051_golden_model_1.ACC [3]);
  and (_03579_, _03558_, \oc8051_golden_model_1.ACC [3]);
  nor (_03580_, _03579_, _03578_);
  and (_03581_, _03580_, _03577_);
  nor (_03582_, _03580_, _03577_);
  nor (_03583_, _03582_, _03581_);
  and (_03584_, _03583_, _03469_);
  not (_03585_, _03584_);
  and (_03586_, _03585_, _03417_);
  nand (_03587_, _03586_, _03576_);
  nand (_03588_, _03587_, _03554_);
  and (_03589_, _03588_, _03549_);
  and (_03590_, _03589_, _03507_);
  nand (_03591_, _03590_, _01958_);
  nand (_03592_, _03484_, _03419_);
  and (_03593_, _03506_, _03592_);
  and (_03594_, _03548_, _03513_);
  and (_03595_, _03588_, _03594_);
  and (_03596_, _03595_, _03593_);
  nand (_03597_, _03596_, _01988_);
  and (_03598_, _03597_, _03591_);
  and (_03599_, _03587_, _03554_);
  and (_03600_, _03599_, _03549_);
  nand (_03601_, _03505_, _03503_);
  and (_03602_, _03601_, _03485_);
  and (_03603_, _03602_, _03600_);
  nand (_03604_, _03603_, _01924_);
  and (_03605_, _03595_, _03507_);
  nand (_03606_, _03605_, _01976_);
  and (_03607_, _03606_, _03604_);
  and (_03608_, _03607_, _03598_);
  and (_03609_, _03600_, _03593_);
  nand (_03610_, _03609_, _01911_);
  and (_03611_, _03601_, _03592_);
  and (_03612_, _03611_, _03600_);
  nand (_03613_, _03612_, _01929_);
  and (_03614_, _03613_, _03610_);
  and (_03615_, _03593_, _03589_);
  nand (_03616_, _03615_, _01967_);
  and (_03617_, _03611_, _03589_);
  nand (_03618_, _03617_, _01980_);
  and (_03619_, _03618_, _03616_);
  and (_03620_, _03619_, _03614_);
  and (_03621_, _03620_, _03608_);
  and (_03623_, _03599_, _03594_);
  and (_03624_, _03623_, _03602_);
  nand (_03625_, _03624_, _01938_);
  and (_03626_, _03623_, _03611_);
  nand (_03627_, _03626_, _01954_);
  and (_03628_, _03627_, _03625_);
  and (_03629_, _03611_, _03595_);
  nand (_03630_, _03629_, _01985_);
  and (_03631_, _03602_, _03595_);
  nand (_03632_, _03631_, _01991_);
  and (_03633_, _03632_, _03630_);
  and (_03634_, _03633_, _03628_);
  and (_03635_, _03600_, _03507_);
  nand (_03636_, _03635_, _42427_);
  and (_03637_, _03602_, _03589_);
  nand (_03638_, _03637_, _01971_);
  and (_03639_, _03638_, _03636_);
  and (_03640_, _03623_, _03507_);
  nand (_03641_, _03640_, _01933_);
  and (_03642_, _03623_, _03593_);
  nand (_03643_, _03642_, _01948_);
  and (_03644_, _03643_, _03641_);
  and (_03645_, _03644_, _03639_);
  and (_03646_, _03645_, _03634_);
  nand (_03647_, _03646_, _03621_);
  nand (_03648_, _03640_, _02260_);
  nand (_03649_, _03596_, _02287_);
  and (_03650_, _03649_, _03648_);
  nand (_03651_, _03635_, _42447_);
  nand (_03652_, _03615_, _02298_);
  and (_03653_, _03652_, _03651_);
  and (_03654_, _03653_, _03650_);
  nand (_03655_, _03624_, _02273_);
  nand (_03656_, _03642_, _02271_);
  and (_03657_, _03656_, _03655_);
  nand (_03658_, _03603_, _02265_);
  nand (_03659_, _03605_, _02293_);
  and (_03660_, _03659_, _03658_);
  and (_03661_, _03660_, _03657_);
  and (_03662_, _03661_, _03654_);
  nand (_03663_, _03590_, _02278_);
  nand (_03664_, _03637_, _02296_);
  and (_03665_, _03664_, _03663_);
  nand (_03666_, _03617_, _02291_);
  nand (_03667_, _03629_, _02283_);
  and (_03668_, _03667_, _03666_);
  and (_03669_, _03668_, _03665_);
  nand (_03670_, _03626_, _02276_);
  nand (_03671_, _03631_, _02285_);
  and (_03672_, _03671_, _03670_);
  nand (_03673_, _03609_, _02267_);
  nand (_03674_, _03612_, _02262_);
  and (_03675_, _03674_, _03673_);
  and (_03676_, _03675_, _03672_);
  and (_03677_, _03676_, _03669_);
  and (_03678_, _03677_, _03662_);
  or (_03679_, _03678_, _03647_);
  nor (_03680_, _03679_, _03375_);
  nor (_03681_, _03647_, _03375_);
  not (_03682_, _03681_);
  not (_03683_, \oc8051_golden_model_1.SP [0]);
  and (_03684_, _03383_, _03683_);
  nand (_03685_, _03605_, _02141_);
  nand (_03686_, _03631_, _02154_);
  and (_03687_, _03686_, _03685_);
  nand (_03688_, _03637_, _02144_);
  nand (_03689_, _03617_, _02139_);
  and (_03690_, _03689_, _03688_);
  and (_03691_, _03690_, _03687_);
  nand (_03692_, _03609_, _02132_);
  nand (_03693_, _03642_, _02118_);
  and (_03694_, _03693_, _03692_);
  nand (_03695_, _03640_, _02129_);
  nand (_03696_, _03626_, _02111_);
  and (_03697_, _03696_, _03695_);
  and (_03698_, _03697_, _03694_);
  and (_03699_, _03698_, _03691_);
  nand (_03700_, _03629_, _02151_);
  nand (_03701_, _03596_, _02156_);
  and (_03702_, _03701_, _03700_);
  nand (_03703_, _03590_, _02114_);
  nand (_03704_, _03615_, _02146_);
  and (_03705_, _03704_, _03703_);
  and (_03706_, _03705_, _03702_);
  nand (_03707_, _03635_, _42432_);
  nand (_03708_, _03603_, _02134_);
  and (_03709_, _03708_, _03707_);
  nand (_03710_, _03612_, _02126_);
  nand (_03711_, _03624_, _02121_);
  and (_03712_, _03711_, _03710_);
  and (_03713_, _03712_, _03709_);
  and (_03714_, _03713_, _03706_);
  and (_03715_, _03714_, _03699_);
  not (_03716_, _03715_);
  not (_03717_, _03339_);
  and (_03718_, _03370_, _03307_);
  and (_03719_, _03718_, _03717_);
  not (_03720_, _03397_);
  nor (_03721_, _03647_, _03720_);
  and (_03722_, _03721_, _03719_);
  not (_03723_, _03722_);
  and (_03724_, _03370_, _03339_);
  not (_03725_, _03724_);
  nor (_03726_, _03725_, _03308_);
  and (_03727_, _03721_, _03726_);
  and (_03728_, _03370_, _03717_);
  and (_03729_, _03728_, _03306_);
  and (_03730_, _03724_, _03308_);
  nor (_03731_, _03730_, _03729_);
  not (_03732_, _03731_);
  and (_03733_, _03721_, _03732_);
  nor (_03734_, _03733_, _03727_);
  and (_03735_, _03734_, _03723_);
  and (_03736_, _03453_, _03306_);
  and (_03737_, _03736_, _03397_);
  not (_03738_, _03737_);
  nor (_03739_, _03738_, _03647_);
  and (_03740_, _03721_, _03454_);
  nor (_03741_, _03740_, _03739_);
  and (_03742_, _03741_, _03735_);
  nor (_03743_, _03742_, _03716_);
  and (_03744_, _03306_, _03275_);
  and (_03745_, _03744_, _03372_);
  and (_03746_, _03745_, _03424_);
  not (_03747_, _03746_);
  nor (_03748_, _03747_, _03679_);
  nor (_03749_, _03428_, _03683_);
  not (_03750_, _03749_);
  not (_03751_, _03427_);
  and (_03752_, _03745_, _03751_);
  not (_03753_, _03752_);
  nor (_03754_, _03753_, _03679_);
  nor (_03755_, _03753_, _03647_);
  not (_03756_, _03755_);
  not (_03757_, _03433_);
  and (_03758_, _03757_, _03373_);
  and (_03759_, _03745_, _03757_);
  not (_03760_, _03759_);
  nor (_03761_, _03760_, _03679_);
  not (_03762_, _03430_);
  and (_03763_, _03745_, _03762_);
  not (_03764_, _03763_);
  or (_03765_, _03764_, _03679_);
  not (_03766_, _03435_);
  and (_03767_, _03724_, _03451_);
  and (_03768_, _03767_, _03766_);
  and (_03769_, _03768_, _03683_);
  not (_03770_, _03768_);
  not (_03771_, _03439_);
  and (_03772_, _03454_, _03412_);
  and (_03773_, _03454_, _03244_);
  not (_03774_, _03773_);
  and (_03775_, _03409_, _03373_);
  not (_03776_, _03775_);
  and (_03777_, _03745_, _03409_);
  not (_03778_, _03777_);
  and (_03779_, _03454_, _03409_);
  and (_03780_, _03615_, _02407_);
  and (_03781_, _03605_, _02409_);
  nor (_03782_, _03781_, _03780_);
  and (_03783_, _03609_, _02422_);
  and (_03784_, _03642_, _02434_);
  nor (_03785_, _03784_, _03783_);
  and (_03786_, _03785_, _03782_);
  and (_03787_, _03631_, _02427_);
  and (_03788_, _03596_, _02417_);
  nor (_03789_, _03788_, _03787_);
  and (_03790_, _03637_, _02415_);
  and (_03791_, _03617_, _02411_);
  nor (_03792_, _03791_, _03790_);
  and (_03793_, _03792_, _03789_);
  and (_03794_, _03793_, _03786_);
  and (_03795_, _03612_, _02398_);
  and (_03796_, _03640_, _02396_);
  nor (_03797_, _03796_, _03795_);
  and (_03798_, _03635_, _42462_);
  and (_03799_, _03603_, _02394_);
  nor (_03800_, _03799_, _03798_);
  and (_03801_, _03800_, _03797_);
  and (_03802_, _03590_, _02430_);
  and (_03803_, _03629_, _02424_);
  nor (_03804_, _03803_, _03802_);
  and (_03805_, _03624_, _02432_);
  and (_03806_, _03626_, _02402_);
  nor (_03807_, _03806_, _03805_);
  and (_03808_, _03807_, _03804_);
  and (_03809_, _03808_, _03801_);
  and (_03810_, _03809_, _03794_);
  nor (_03811_, _03810_, _03647_);
  not (_03812_, _03678_);
  and (_03813_, _03812_, _03647_);
  nor (_03814_, _03813_, _03811_);
  and (_03815_, _03745_, _03400_);
  and (_03816_, _03745_, _03397_);
  nor (_03817_, _03816_, _03815_);
  not (_03818_, _03817_);
  and (_03819_, _03818_, _03814_);
  not (_03820_, _03455_);
  not (_03821_, _03440_);
  and (_03822_, _03728_, _03744_);
  and (_03824_, _03822_, _03821_);
  and (_03825_, _03728_, _03451_);
  and (_03826_, _03825_, _03821_);
  or (_03827_, _03826_, _03824_);
  and (_03828_, _03724_, _03306_);
  and (_03829_, _03828_, _03821_);
  nor (_03830_, _03829_, _03827_);
  and (_03831_, _03728_, _03308_);
  and (_03832_, _03831_, _03821_);
  not (_03833_, _03832_);
  and (_03834_, _03728_, _03422_);
  and (_03835_, _03834_, _03821_);
  and (_03836_, _03724_, _03307_);
  and (_03837_, _03836_, _03821_);
  nor (_03838_, _03837_, _03835_);
  and (_03839_, _03838_, _03833_);
  and (_03840_, _03839_, _03830_);
  not (_03841_, _03840_);
  and (_03842_, _03841_, _03678_);
  and (_03843_, _03751_, _03373_);
  nor (_03844_, _03843_, _03752_);
  nor (_03845_, _03844_, _03814_);
  nand (_03846_, _03763_, _03814_);
  not (_03847_, \oc8051_golden_model_1.SP [3]);
  and (_03848_, _03762_, _03373_);
  nand (_03849_, _03848_, _03847_);
  and (_03850_, _03454_, _03762_);
  and (_03851_, _03454_, _03766_);
  nor (_03852_, _03851_, _03850_);
  nor (_03853_, _03852_, _03678_);
  and (_03854_, _03454_, _03757_);
  not (_03855_, _03854_);
  nor (_03856_, _03848_, _03763_);
  not (_03857_, _03856_);
  and (_03858_, _03852_, \oc8051_golden_model_1.PSW [3]);
  or (_03859_, _03858_, _03857_);
  and (_03860_, _03859_, _03855_);
  or (_03861_, _03860_, _03853_);
  and (_03862_, _03861_, _03849_);
  and (_03863_, _03862_, _03846_);
  nor (_03864_, _03855_, _03678_);
  or (_03865_, _03864_, _03863_);
  and (_03866_, _03865_, _03760_);
  or (_03867_, _03814_, _03760_);
  and (_03868_, _03454_, _03751_);
  nor (_03869_, _03868_, _03758_);
  nand (_03870_, _03869_, _03867_);
  or (_03871_, _03870_, _03866_);
  or (_03872_, _03869_, _03812_);
  and (_03873_, _03844_, _03872_);
  and (_03874_, _03873_, _03871_);
  or (_03875_, _03874_, _03841_);
  nor (_03876_, _03875_, _03845_);
  nor (_03877_, _03876_, _03842_);
  and (_03878_, _03821_, _03373_);
  and (_03879_, _03745_, _03821_);
  nor (_03880_, _03879_, _03878_);
  not (_03881_, _03880_);
  nor (_03882_, _03881_, _03877_);
  and (_03883_, _03454_, _03424_);
  and (_03884_, _03881_, _03814_);
  nor (_03885_, _03884_, _03883_);
  not (_03886_, _03885_);
  nor (_03887_, _03886_, _03882_);
  not (_03888_, _03883_);
  nor (_03889_, _03888_, _03678_);
  or (_03890_, _03889_, _03887_);
  and (_03891_, _03890_, _03747_);
  nor (_03892_, _03814_, _03747_);
  or (_03893_, _03892_, _03891_);
  and (_03894_, _03893_, _03820_);
  and (_03895_, _03724_, _03744_);
  and (_03896_, _03895_, _03751_);
  and (_03897_, _03423_, _03404_);
  nor (_03898_, _03897_, _03896_);
  and (_03899_, _03745_, _03244_);
  not (_03900_, _03899_);
  and (_03901_, _03745_, _03412_);
  nor (_03902_, _03901_, _03374_);
  and (_03903_, _03454_, _03400_);
  nor (_03904_, _03775_, _03903_);
  and (_03905_, _03904_, _03902_);
  and (_03906_, _03905_, _03900_);
  and (_03907_, _03906_, _03898_);
  and (_03908_, _03423_, _03387_);
  not (_03909_, _03908_);
  and (_03910_, _03724_, _03422_);
  and (_03911_, _03910_, _03751_);
  nor (_03912_, _03911_, _03850_);
  and (_03913_, _03382_, _03373_);
  and (_03914_, _03423_, _03392_);
  nor (_03915_, _03914_, _03913_);
  and (_03916_, _03915_, _03912_);
  and (_03917_, _03916_, _03909_);
  not (_03918_, _03868_);
  and (_03919_, _03453_, _03308_);
  and (_03920_, _03919_, _03751_);
  and (_03921_, _03424_, _03373_);
  nor (_03922_, _03921_, _03920_);
  and (_03923_, _03922_, _03918_);
  and (_03924_, _03729_, _03751_);
  and (_03925_, _03736_, _03751_);
  nor (_03926_, _03925_, _03924_);
  and (_03927_, _03836_, _03751_);
  and (_03928_, _03719_, _03751_);
  nor (_03929_, _03928_, _03927_);
  and (_03930_, _03929_, _03926_);
  and (_03931_, _03930_, _03923_);
  and (_03932_, _03931_, _03917_);
  and (_03933_, _03932_, _03907_);
  nor (_03934_, _03933_, _03510_);
  not (_03935_, _03518_);
  and (_03936_, _03933_, _03935_);
  nor (_03937_, _03936_, _03934_);
  not (_03938_, _03552_);
  nor (_03939_, _03933_, _03938_);
  and (_03940_, _03933_, _03559_);
  nor (_03941_, _03940_, _03939_);
  not (_03942_, _03941_);
  and (_03943_, _03942_, _03937_);
  nor (_03944_, _03933_, _03119_);
  and (_03945_, _03933_, _03119_);
  nor (_03946_, _03945_, _03944_);
  nor (_03947_, _03933_, \oc8051_golden_model_1.PC [1]);
  not (_03948_, _03447_);
  and (_03949_, _03933_, _03948_);
  nor (_03950_, _03949_, _03947_);
  nor (_03951_, _03950_, _03946_);
  and (_03952_, _03951_, _03943_);
  and (_03953_, _03952_, _42447_);
  not (_03954_, _03946_);
  and (_03955_, _03950_, _03954_);
  nor (_03956_, _03941_, _03937_);
  and (_03957_, _03956_, _03955_);
  and (_03958_, _03957_, _02271_);
  nor (_03959_, _03958_, _03953_);
  and (_03960_, _03941_, _03937_);
  and (_03961_, _03960_, _03955_);
  and (_03962_, _03961_, _02298_);
  and (_03963_, _03946_, \oc8051_golden_model_1.PC [1]);
  nor (_03964_, _03942_, _03937_);
  and (_03965_, _03964_, _03963_);
  and (_03966_, _03965_, _02283_);
  nor (_03967_, _03966_, _03962_);
  and (_03968_, _03967_, _03959_);
  and (_03969_, _03960_, _03951_);
  and (_03970_, _03969_, _02278_);
  and (_03971_, _03960_, _03963_);
  and (_03972_, _03971_, _02291_);
  nor (_03973_, _03972_, _03970_);
  and (_03974_, _03955_, _03943_);
  and (_03975_, _03974_, _02267_);
  and (_03976_, _03963_, _03943_);
  and (_03977_, _03976_, _02262_);
  nor (_03978_, _03977_, _03975_);
  and (_03979_, _03978_, _03973_);
  and (_03980_, _03979_, _03968_);
  and (_03981_, _03946_, _03087_);
  and (_03982_, _03956_, _03981_);
  and (_03983_, _03982_, _02273_);
  and (_03984_, _03956_, _03963_);
  and (_03985_, _03984_, _02276_);
  nor (_03986_, _03985_, _03983_);
  and (_03987_, _03964_, _03951_);
  and (_03988_, _03987_, _02293_);
  and (_03989_, _03964_, _03955_);
  and (_03990_, _03989_, _02287_);
  nor (_03991_, _03990_, _03988_);
  and (_03992_, _03991_, _03986_);
  and (_03993_, _03981_, _03943_);
  and (_03994_, _03993_, _02265_);
  and (_03995_, _03960_, _03981_);
  and (_03996_, _03995_, _02296_);
  nor (_03997_, _03996_, _03994_);
  and (_03998_, _03956_, _03951_);
  and (_03999_, _03998_, _02260_);
  and (_04000_, _03964_, _03981_);
  and (_04001_, _04000_, _02285_);
  nor (_04002_, _04001_, _03999_);
  and (_04003_, _04002_, _03997_);
  and (_04004_, _04003_, _03992_);
  and (_04005_, _04004_, _03980_);
  nor (_04006_, _04005_, _03820_);
  nor (_04007_, _04006_, _03818_);
  not (_04008_, _04007_);
  nor (_04009_, _04008_, _03894_);
  nor (_04010_, _04009_, _03819_);
  and (_04011_, _03745_, _03392_);
  nor (_04012_, _04011_, _03914_);
  and (_04013_, _03454_, _03392_);
  not (_04014_, _04013_);
  and (_04015_, _04014_, _04012_);
  and (_04016_, _03454_, _03404_);
  not (_04017_, _04016_);
  and (_04018_, _03745_, _03404_);
  nor (_04019_, _04018_, _03897_);
  and (_04020_, _04019_, _04017_);
  and (_04021_, _04020_, _04015_);
  and (_04022_, _03454_, _03382_);
  not (_04023_, _04022_);
  and (_04025_, _03454_, _03387_);
  not (_04026_, _04025_);
  and (_04027_, _03745_, _03387_);
  nor (_04028_, _04027_, _03908_);
  and (_04029_, _04028_, _04026_);
  and (_04030_, _04029_, _04023_);
  and (_04031_, _04030_, _04021_);
  not (_04032_, _04031_);
  nor (_04033_, _04032_, _04010_);
  and (_04034_, _03745_, _03382_);
  and (_04035_, _04032_, _03678_);
  nor (_04036_, _04035_, _04034_);
  not (_04037_, _04036_);
  nor (_04038_, _04037_, _04033_);
  and (_04039_, _04034_, \oc8051_golden_model_1.SP [3]);
  or (_04040_, _04039_, _03913_);
  or (_04041_, _04040_, _04038_);
  nand (_04042_, _03814_, _03913_);
  and (_04043_, _04042_, _04041_);
  nor (_04044_, _04043_, _03779_);
  and (_04045_, _03779_, _03678_);
  nor (_04046_, _04045_, _04044_);
  and (_04047_, _04046_, _03778_);
  and (_04048_, _03777_, \oc8051_golden_model_1.SP [3]);
  or (_04049_, _04048_, _04047_);
  and (_04050_, _04049_, _03776_);
  nor (_04051_, _03776_, _03814_);
  or (_04052_, _04051_, _04050_);
  and (_04053_, _04052_, _03774_);
  nor (_04054_, _03774_, _03678_);
  or (_04055_, _04054_, _04053_);
  and (_04056_, _04055_, _03375_);
  nor (_04057_, _03814_, _03375_);
  nor (_04058_, _04057_, _04056_);
  nor (_04059_, _04058_, _03772_);
  not (_04060_, _03772_);
  nor (_04061_, _04060_, _03678_);
  nor (_04062_, _04061_, _04059_);
  and (_04063_, _03635_, _42457_);
  and (_04064_, _03617_, _02366_);
  nor (_04065_, _04064_, _04063_);
  and (_04066_, _03609_, _02377_);
  and (_04067_, _03626_, _02357_);
  nor (_04068_, _04067_, _04066_);
  and (_04069_, _04068_, _04065_);
  and (_04070_, _03596_, _02372_);
  and (_04071_, _03631_, _02381_);
  nor (_04072_, _04071_, _04070_);
  and (_04073_, _03640_, _02351_);
  and (_04074_, _03605_, _02364_);
  nor (_04075_, _04074_, _04073_);
  and (_04076_, _04075_, _04072_);
  and (_04077_, _04076_, _04069_);
  and (_04078_, _03603_, _02349_);
  and (_04079_, _03612_, _02353_);
  nor (_04080_, _04079_, _04078_);
  and (_04081_, _03642_, _02388_);
  and (_04082_, _03590_, _02384_);
  nor (_04083_, _04082_, _04081_);
  and (_04084_, _04083_, _04080_);
  and (_04085_, _03624_, _02386_);
  and (_04086_, _03637_, _02370_);
  nor (_04087_, _04086_, _04085_);
  and (_04088_, _03615_, _02362_);
  and (_04089_, _03629_, _02379_);
  nor (_04090_, _04089_, _04088_);
  and (_04091_, _04090_, _04087_);
  and (_04092_, _04091_, _04084_);
  and (_04093_, _04092_, _04077_);
  nor (_04094_, _04093_, _03647_);
  and (_04095_, _04094_, _03374_);
  not (_04096_, _04095_);
  not (_04097_, _03913_);
  nor (_04098_, _03775_, _03763_);
  and (_04099_, _04098_, _04097_);
  nor (_04100_, _03759_, _03746_);
  and (_04101_, _04100_, _03817_);
  and (_04102_, _03880_, _03844_);
  and (_04103_, _04102_, _04101_);
  and (_04104_, _04103_, _04099_);
  not (_04105_, _04104_);
  and (_04106_, _04105_, _04094_);
  not (_04107_, _04106_);
  and (_04108_, _03640_, _02216_);
  and (_04109_, _03590_, _02249_);
  nor (_04110_, _04109_, _04108_);
  and (_04111_, _03637_, _02235_);
  and (_04112_, _03629_, _02244_);
  nor (_04113_, _04112_, _04111_);
  and (_04114_, _04113_, _04110_);
  and (_04115_, _03609_, _02242_);
  and (_04116_, _03603_, _02214_);
  nor (_04117_, _04116_, _04115_);
  and (_04118_, _03635_, _42442_);
  and (_04119_, _03605_, _02229_);
  nor (_04120_, _04119_, _04118_);
  and (_04121_, _04120_, _04117_);
  and (_04122_, _04121_, _04114_);
  and (_04123_, _03615_, _02227_);
  and (_04124_, _03617_, _02231_);
  nor (_04126_, _04124_, _04123_);
  and (_04127_, _03624_, _02251_);
  and (_04128_, _03596_, _02237_);
  nor (_04129_, _04128_, _04127_);
  and (_04130_, _04129_, _04126_);
  and (_04131_, _03612_, _02218_);
  and (_04132_, _03631_, _02246_);
  nor (_04133_, _04132_, _04131_);
  and (_04134_, _03642_, _02253_);
  and (_04135_, _03626_, _02222_);
  nor (_04136_, _04135_, _04134_);
  and (_04137_, _04136_, _04133_);
  and (_04138_, _04137_, _04130_);
  and (_04139_, _04138_, _04122_);
  not (_04140_, _03779_);
  nor (_04141_, _03883_, _03854_);
  and (_04142_, _04141_, _04140_);
  and (_04143_, _03869_, _03852_);
  nor (_04144_, _03773_, _03772_);
  and (_04145_, _04144_, _04143_);
  and (_04146_, _04145_, _04142_);
  and (_04147_, _04146_, _04031_);
  and (_04148_, _04147_, _03840_);
  nor (_04149_, _04148_, _04139_);
  and (_04150_, _03952_, _42442_);
  and (_04151_, _03961_, _02227_);
  nor (_04152_, _04151_, _04150_);
  and (_04153_, _03974_, _02242_);
  and (_04154_, _03957_, _02253_);
  nor (_04155_, _04154_, _04153_);
  and (_04156_, _04155_, _04152_);
  and (_04157_, _03998_, _02216_);
  and (_04158_, _03987_, _02229_);
  nor (_04159_, _04158_, _04157_);
  and (_04160_, _03965_, _02244_);
  and (_04161_, _04000_, _02246_);
  nor (_04162_, _04161_, _04160_);
  and (_04163_, _04162_, _04159_);
  and (_04164_, _04163_, _04156_);
  and (_04165_, _03993_, _02214_);
  and (_04166_, _03976_, _02218_);
  nor (_04167_, _04166_, _04165_);
  and (_04168_, _03984_, _02222_);
  and (_04169_, _03995_, _02235_);
  nor (_04170_, _04169_, _04168_);
  and (_04171_, _04170_, _04167_);
  and (_04172_, _03982_, _02251_);
  and (_04173_, _03969_, _02249_);
  nor (_04174_, _04173_, _04172_);
  and (_04175_, _03971_, _02231_);
  and (_04176_, _03989_, _02237_);
  nor (_04177_, _04176_, _04175_);
  and (_04178_, _04177_, _04174_);
  and (_04179_, _04178_, _04171_);
  and (_04180_, _04179_, _04164_);
  nor (_04181_, _04180_, _03820_);
  not (_04182_, \oc8051_golden_model_1.SP [2]);
  nor (_04183_, _04034_, _03777_);
  nor (_04184_, _04183_, _04182_);
  not (_04185_, _04184_);
  nand (_04186_, _03724_, _03387_);
  and (_04187_, _03828_, _03751_);
  and (_04188_, _03828_, _03757_);
  nor (_04189_, _04188_, _04187_);
  and (_04190_, _03828_, _03424_);
  and (_04191_, _03828_, _03397_);
  nor (_04192_, _04191_, _04190_);
  and (_04193_, _04192_, _04189_);
  and (_04194_, _04193_, _04186_);
  and (_04195_, _04194_, _04185_);
  and (_04196_, _03836_, _03244_);
  and (_04197_, _03828_, _03412_);
  nor (_04198_, _04197_, _04196_);
  and (_04199_, _03836_, _03412_);
  and (_04200_, _03828_, _03244_);
  nor (_04201_, _04200_, _04199_);
  and (_04202_, _04201_, _04198_);
  and (_04203_, _03828_, _03382_);
  and (_04204_, _03836_, _03404_);
  nor (_04205_, _04204_, _04203_);
  and (_04206_, _03828_, _03409_);
  and (_04207_, _03836_, _03392_);
  nor (_04208_, _04207_, _04206_);
  and (_04209_, _04208_, _04205_);
  and (_04210_, _03386_, _03209_);
  and (_04211_, _04210_, _03828_);
  and (_04212_, _03836_, _03424_);
  nor (_04213_, _04212_, _04211_);
  and (_04214_, _03836_, _03397_);
  and (_04215_, _03836_, _03409_);
  nor (_04216_, _04215_, _04214_);
  and (_04217_, _04216_, _04213_);
  and (_04218_, _04217_, _04209_);
  and (_04219_, _04218_, _04202_);
  and (_04220_, _03730_, _03382_);
  not (_04221_, _04220_);
  and (_04222_, _03848_, \oc8051_golden_model_1.SP [2]);
  and (_04223_, _03730_, _03766_);
  nor (_04224_, _04223_, _04222_);
  and (_04225_, _04224_, _04221_);
  and (_04227_, _03836_, _03757_);
  nor (_04228_, _03725_, _03430_);
  nor (_04229_, _04228_, _04227_);
  and (_04230_, _03828_, _03766_);
  nor (_04231_, _04230_, _03927_);
  and (_04232_, _04231_, _04229_);
  and (_04233_, _03767_, _03382_);
  nor (_04234_, _04233_, _03768_);
  and (_04235_, _04234_, _04232_);
  and (_04236_, _04235_, _04225_);
  and (_04237_, _04236_, _04219_);
  and (_04238_, _04237_, _04195_);
  not (_04239_, _04238_);
  nor (_04240_, _04239_, _04181_);
  not (_04241_, _04240_);
  nor (_04242_, _04241_, _04149_);
  and (_04243_, _04242_, _04107_);
  and (_04244_, _04243_, _04096_);
  not (_04245_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_04246_, _03715_, _04060_);
  not (_04247_, _04246_);
  nor (_04248_, _03715_, _03888_);
  nor (_04249_, _03880_, _03679_);
  nor (_04250_, _03715_, _03918_);
  or (_04251_, _03715_, _03855_);
  nor (_04252_, _03715_, _03852_);
  and (_04253_, _03744_, _03453_);
  nor (_04254_, _04253_, _03831_);
  not (_04255_, _03822_);
  nor (_04256_, _03730_, _03454_);
  and (_04257_, _04256_, _04255_);
  and (_04258_, _04257_, _04254_);
  nor (_04259_, _04258_, _03435_);
  not (_04260_, _04259_);
  not (_04261_, _03438_);
  and (_04262_, _04253_, _04261_);
  and (_04263_, _03895_, _03766_);
  nor (_04264_, _04263_, _04262_);
  and (_04265_, _03728_, _03762_);
  nor (_04266_, _04265_, _04228_);
  not (_04267_, _04266_);
  and (_04268_, _04267_, _03744_);
  and (_04269_, _03831_, _03762_);
  nor (_04270_, _04269_, _03850_);
  and (_04271_, _03730_, _03762_);
  and (_04272_, _04253_, _03762_);
  nor (_04273_, _04272_, _04271_);
  and (_04274_, _04273_, _04270_);
  not (_04275_, _04274_);
  nor (_04276_, _04275_, _04268_);
  and (_04277_, _04276_, _04264_);
  and (_04278_, _04277_, _04260_);
  or (_04279_, _04278_, _04252_);
  nand (_04280_, _04279_, _03764_);
  nand (_04281_, _03765_, _04280_);
  and (_04282_, _03728_, _03757_);
  and (_04283_, _04282_, _03306_);
  nor (_04284_, _04283_, _04188_);
  nor (_04285_, _04284_, _03420_);
  not (_04286_, _04285_);
  and (_04287_, _03831_, _03757_);
  and (_04288_, _03848_, _03683_);
  nor (_04289_, _04288_, _04287_);
  not (_04290_, _03730_);
  nor (_04291_, _04253_, _03454_);
  and (_04292_, _04291_, _04290_);
  nor (_04293_, _04292_, _03433_);
  not (_04294_, _04293_);
  and (_04295_, _04294_, _04289_);
  and (_04296_, _04295_, _04286_);
  nand (_04297_, _04296_, _04281_);
  nand (_04298_, _04297_, _04251_);
  and (_04299_, _04298_, _03760_);
  or (_04300_, _03761_, _04299_);
  and (_04301_, _03715_, _03758_);
  nor (_04302_, _03927_, _03924_);
  or (_04303_, _04302_, _03420_);
  and (_04304_, _04253_, _03751_);
  not (_04305_, _04304_);
  and (_04306_, _03831_, _03751_);
  or (_04307_, _04306_, _03868_);
  nor (_04308_, _04307_, _03896_);
  and (_04309_, _04308_, _04305_);
  and (_04310_, _04309_, _04303_);
  not (_04311_, _04310_);
  nor (_04312_, _04311_, _04301_);
  and (_04313_, _04312_, _04300_);
  or (_04314_, _04313_, _04250_);
  nand (_04315_, _04314_, _03844_);
  nor (_04316_, _03844_, _03679_);
  nor (_04317_, _04316_, _03841_);
  nand (_04318_, _04317_, _04315_);
  and (_04319_, _03715_, _03841_);
  and (_04320_, _04253_, _03821_);
  nor (_04321_, _04320_, _03881_);
  not (_04322_, _04321_);
  nor (_04323_, _04322_, _04319_);
  and (_04324_, _04323_, _04318_);
  or (_04325_, _04324_, _04249_);
  nor (_04326_, _04212_, _04190_);
  nor (_04328_, _04326_, _03420_);
  not (_04329_, _04328_);
  and (_04330_, _03736_, _03424_);
  and (_04331_, _04330_, _03275_);
  not (_04332_, _04331_);
  and (_04333_, _03822_, _03424_);
  not (_04334_, _04333_);
  and (_04335_, _03831_, _03424_);
  nor (_04336_, _04335_, _03883_);
  and (_04337_, _04336_, _04334_);
  and (_04338_, _04337_, _04332_);
  and (_04339_, _04338_, _04329_);
  and (_04340_, _04339_, _04325_);
  or (_04341_, _04340_, _04248_);
  and (_04342_, _04341_, _03747_);
  or (_04343_, _04342_, _03748_);
  and (_04344_, _03730_, _03397_);
  not (_04345_, _04344_);
  nor (_04346_, _03895_, _03454_);
  and (_04347_, _04346_, _04255_);
  and (_04348_, _04347_, _04254_);
  or (_04349_, _04348_, _03720_);
  and (_04350_, _04349_, _04345_);
  and (_04351_, _04350_, _04343_);
  and (_04352_, _03952_, _42432_);
  and (_04353_, _03989_, _02156_);
  nor (_04354_, _04353_, _04352_);
  and (_04355_, _03998_, _02129_);
  and (_04356_, _03965_, _02151_);
  nor (_04357_, _04356_, _04355_);
  and (_04358_, _04357_, _04354_);
  and (_04359_, _03957_, _02118_);
  and (_04360_, _04000_, _02154_);
  nor (_04361_, _04360_, _04359_);
  and (_04362_, _03995_, _02144_);
  and (_04363_, _03971_, _02139_);
  nor (_04364_, _04363_, _04362_);
  and (_04365_, _04364_, _04361_);
  and (_04366_, _04365_, _04358_);
  and (_04367_, _03961_, _02146_);
  and (_04368_, _03987_, _02141_);
  nor (_04369_, _04368_, _04367_);
  and (_04370_, _03974_, _02132_);
  and (_04371_, _03982_, _02121_);
  nor (_04372_, _04371_, _04370_);
  and (_04373_, _04372_, _04369_);
  and (_04374_, _03993_, _02134_);
  and (_04375_, _03984_, _02111_);
  nor (_04376_, _04375_, _04374_);
  and (_04377_, _03976_, _02126_);
  and (_04378_, _03969_, _02114_);
  nor (_04379_, _04378_, _04377_);
  and (_04380_, _04379_, _04376_);
  and (_04381_, _04380_, _04373_);
  and (_04382_, _04381_, _04366_);
  nor (_04383_, _04382_, _03820_);
  or (_04384_, _04383_, _04351_);
  and (_04385_, _03816_, _03679_);
  and (_04386_, _04253_, _03400_);
  nor (_04387_, _04386_, _03815_);
  not (_04388_, _04387_);
  nor (_04389_, _04388_, _04385_);
  and (_04390_, _04389_, _04384_);
  not (_04391_, _03815_);
  nor (_04392_, _04391_, _03679_);
  or (_04393_, _04392_, _04390_);
  and (_04394_, _03822_, _03404_);
  not (_04395_, _04394_);
  and (_04396_, _03895_, _03404_);
  and (_04397_, _03831_, _03404_);
  nor (_04398_, _04397_, _04396_);
  and (_04399_, _04398_, _04395_);
  and (_04400_, _03730_, _03404_);
  and (_04401_, _04253_, _03404_);
  nor (_04402_, _04401_, _04400_);
  and (_04403_, _04402_, _04399_);
  and (_04404_, _04403_, _04393_);
  nor (_04405_, _03716_, _04020_);
  and (_04406_, _03730_, _03387_);
  not (_04407_, _04406_);
  and (_04408_, _03895_, _03387_);
  and (_04409_, _03831_, _03387_);
  nor (_04410_, _04409_, _04408_);
  and (_04411_, _04410_, _04407_);
  and (_04412_, _03822_, _03387_);
  and (_04413_, _04253_, _03387_);
  nor (_04414_, _04413_, _04412_);
  and (_04415_, _04414_, _04411_);
  not (_04416_, _04415_);
  nor (_04417_, _04416_, _04405_);
  and (_04418_, _04417_, _04404_);
  nor (_04419_, _03716_, _04029_);
  not (_04420_, _03392_);
  and (_04421_, _03370_, _03275_);
  and (_04422_, _04421_, _03339_);
  nor (_04423_, _04422_, _03822_);
  and (_04424_, _04423_, _04254_);
  nor (_04425_, _04424_, _04420_);
  nor (_04426_, _04425_, _04419_);
  and (_04427_, _04426_, _04418_);
  nor (_04429_, _03716_, _04015_);
  and (_04430_, _03895_, _03382_);
  nor (_04431_, _04430_, _04022_);
  and (_04432_, _03822_, _03382_);
  not (_04433_, _04432_);
  and (_04434_, _03831_, _03382_);
  and (_04435_, _04253_, _03382_);
  nor (_04436_, _04435_, _04434_);
  and (_04437_, _04436_, _04433_);
  and (_04438_, _04437_, _04221_);
  and (_04439_, _04438_, _04431_);
  not (_04440_, _04439_);
  nor (_04441_, _04440_, _04429_);
  and (_04442_, _04441_, _04427_);
  nor (_04443_, _03715_, _04023_);
  or (_04444_, _04443_, _04442_);
  and (_04445_, _04034_, _03683_);
  nor (_04446_, _04445_, _03913_);
  and (_04447_, _04446_, _04444_);
  nor (_04448_, _04097_, _03679_);
  or (_04449_, _04448_, _04447_);
  and (_04450_, _03822_, _03409_);
  not (_04451_, _04450_);
  not (_04452_, _03409_);
  and (_04453_, _04346_, _04290_);
  nor (_04454_, _04453_, _04452_);
  and (_04455_, _04253_, _03409_);
  and (_04456_, _03831_, _03409_);
  or (_04457_, _04456_, _04455_);
  nor (_04458_, _04457_, _04454_);
  and (_04459_, _04458_, _04451_);
  and (_04460_, _04459_, _04449_);
  nor (_04461_, _03715_, _04140_);
  or (_04462_, _04461_, _04460_);
  and (_04463_, _03777_, _03683_);
  nor (_04464_, _04463_, _03775_);
  and (_04465_, _04464_, _04462_);
  nor (_04466_, _03776_, _03679_);
  or (_04467_, _04466_, _04465_);
  nand (_04468_, _03724_, _03244_);
  or (_04469_, _04468_, _03420_);
  and (_04470_, _03822_, _03244_);
  and (_04471_, _04253_, _03244_);
  and (_04472_, _03831_, _03244_);
  or (_04473_, _04472_, _03773_);
  or (_04474_, _04473_, _04471_);
  nor (_04475_, _04474_, _04470_);
  and (_04476_, _04475_, _04469_);
  and (_04477_, _04476_, _04467_);
  nor (_04478_, _03715_, _03774_);
  or (_04479_, _04478_, _04477_);
  and (_04480_, _04479_, _03375_);
  or (_04481_, _04480_, _03680_);
  nand (_04482_, _03412_, _03370_);
  not (_04483_, _04482_);
  nand (_04484_, _04483_, _03744_);
  and (_04485_, _03728_, _03412_);
  nand (_04486_, _04485_, _03308_);
  and (_04487_, _04486_, _04060_);
  and (_04488_, _03730_, _03412_);
  and (_04489_, _04253_, _03412_);
  nor (_04490_, _04489_, _04488_);
  and (_04491_, _04490_, _04487_);
  and (_04492_, _04491_, _04484_);
  nand (_04493_, _04492_, _04481_);
  nand (_04494_, _04493_, _04247_);
  or (_04495_, _04494_, _04245_);
  and (_04496_, _03590_, _02312_);
  and (_04497_, _03605_, _02319_);
  nor (_04498_, _04497_, _04496_);
  and (_04499_, _03603_, _02304_);
  and (_04500_, _03642_, _02343_);
  nor (_04501_, _04500_, _04499_);
  and (_04502_, _04501_, _04498_);
  and (_04503_, _03631_, _02336_);
  and (_04504_, _03596_, _02327_);
  nor (_04505_, _04504_, _04503_);
  and (_04506_, _03637_, _02325_);
  and (_04507_, _03617_, _02321_);
  nor (_04508_, _04507_, _04506_);
  and (_04509_, _04508_, _04505_);
  and (_04510_, _04509_, _04502_);
  and (_04511_, _03612_, _02308_);
  and (_04512_, _03640_, _02306_);
  nor (_04513_, _04512_, _04511_);
  and (_04514_, _03635_, _42452_);
  and (_04515_, _03609_, _02332_);
  nor (_04516_, _04515_, _04514_);
  and (_04517_, _04516_, _04513_);
  and (_04518_, _03615_, _02317_);
  and (_04519_, _03629_, _02334_);
  nor (_04520_, _04519_, _04518_);
  and (_04521_, _03624_, _02341_);
  and (_04522_, _03626_, _02339_);
  nor (_04523_, _04522_, _04521_);
  and (_04524_, _04523_, _04520_);
  and (_04525_, _04524_, _04517_);
  and (_04526_, _04525_, _04510_);
  nor (_04527_, _04526_, _03647_);
  and (_04528_, _04527_, _04105_);
  not (_04530_, _04528_);
  and (_04531_, _04527_, _03374_);
  not (_04532_, _04531_);
  and (_04533_, _03635_, _42437_);
  and (_04534_, _03640_, _02183_);
  nor (_04535_, _04534_, _04533_);
  and (_04536_, _03637_, _02200_);
  and (_04537_, _03596_, _02208_);
  nor (_04538_, _04537_, _04536_);
  and (_04539_, _04538_, _04535_);
  and (_04540_, _03603_, _02188_);
  and (_04541_, _03612_, _02181_);
  nor (_04542_, _04541_, _04540_);
  and (_04543_, _03624_, _02175_);
  and (_04544_, _03626_, _02169_);
  nor (_04545_, _04544_, _04543_);
  and (_04546_, _04545_, _04542_);
  and (_04547_, _04546_, _04539_);
  and (_04548_, _03617_, _02193_);
  and (_04549_, _03605_, _02195_);
  nor (_04550_, _04549_, _04548_);
  and (_04551_, _03590_, _02166_);
  and (_04552_, _03615_, _02198_);
  nor (_04553_, _04552_, _04551_);
  and (_04554_, _04553_, _04550_);
  and (_04555_, _03609_, _02186_);
  and (_04556_, _03642_, _02173_);
  nor (_04557_, _04556_, _04555_);
  and (_04558_, _03629_, _02204_);
  and (_04559_, _03631_, _02206_);
  nor (_04560_, _04559_, _04558_);
  and (_04561_, _04560_, _04557_);
  and (_04562_, _04561_, _04554_);
  and (_04563_, _04562_, _04547_);
  nor (_04564_, _04563_, _04148_);
  and (_04565_, _03969_, _02166_);
  and (_04566_, _03965_, _02204_);
  nor (_04567_, _04566_, _04565_);
  and (_04568_, _03984_, _02169_);
  and (_04569_, _03987_, _02195_);
  nor (_04570_, _04569_, _04568_);
  and (_04571_, _04570_, _04567_);
  and (_04572_, _03998_, _02183_);
  and (_04573_, _03989_, _02208_);
  nor (_04574_, _04573_, _04572_);
  and (_04575_, _03952_, _42437_);
  and (_04576_, _03976_, _02181_);
  nor (_04577_, _04576_, _04575_);
  and (_04578_, _04577_, _04574_);
  and (_04579_, _04578_, _04571_);
  and (_04580_, _03993_, _02188_);
  and (_04581_, _04000_, _02206_);
  nor (_04582_, _04581_, _04580_);
  and (_04583_, _03957_, _02173_);
  and (_04584_, _03995_, _02200_);
  nor (_04585_, _04584_, _04583_);
  and (_04586_, _04585_, _04582_);
  and (_04587_, _03982_, _02175_);
  and (_04588_, _03961_, _02198_);
  nor (_04589_, _04588_, _04587_);
  and (_04590_, _03974_, _02186_);
  and (_04591_, _03971_, _02193_);
  nor (_04592_, _04591_, _04590_);
  and (_04593_, _04592_, _04589_);
  and (_04594_, _04593_, _04586_);
  and (_04595_, _04594_, _04579_);
  nor (_04596_, _04595_, _03820_);
  and (_04597_, _03828_, _03762_);
  nor (_04598_, _04597_, _04206_);
  and (_04599_, _03828_, _03387_);
  and (_04600_, _03386_, _03379_);
  and (_04601_, _03729_, _04600_);
  nor (_04602_, _04601_, _04599_);
  and (_04603_, _04602_, _04598_);
  and (_04604_, _04603_, _04193_);
  not (_04605_, \oc8051_golden_model_1.SP [1]);
  nor (_04606_, _03848_, _03777_);
  nor (_04607_, _04606_, _04605_);
  not (_04608_, _03729_);
  not (_04609_, _03424_);
  and (_04610_, _03435_, _04609_);
  nor (_04611_, _03397_, _03404_);
  and (_04612_, _04611_, _04610_);
  nor (_04613_, _04612_, _04608_);
  nor (_04614_, _04613_, _04607_);
  and (_04615_, _04614_, _04604_);
  and (_04616_, _03834_, _03382_);
  not (_04617_, _04616_);
  and (_04618_, _04034_, \oc8051_golden_model_1.SP [1]);
  nor (_04619_, _04618_, _04283_);
  and (_04620_, _04619_, _04617_);
  and (_04621_, _03834_, _03409_);
  nor (_04622_, _04621_, _04450_);
  nor (_04623_, _04432_, _04197_);
  and (_04624_, _04623_, _04622_);
  nor (_04625_, _04230_, _03924_);
  nor (_04626_, _04211_, _04203_);
  and (_04627_, _04626_, _04625_);
  and (_04628_, _03729_, _03762_);
  and (_04629_, _03729_, _03412_);
  nor (_04631_, _04629_, _04628_);
  and (_04632_, _03729_, _03244_);
  nor (_04633_, _04632_, _04200_);
  and (_04634_, _04633_, _04631_);
  and (_04635_, _04634_, _04627_);
  and (_04636_, _04635_, _04624_);
  and (_04637_, _04636_, _04620_);
  and (_04638_, _04637_, _04615_);
  not (_04639_, _04638_);
  nor (_04640_, _04639_, _04596_);
  not (_04641_, _04640_);
  nor (_04642_, _04641_, _04564_);
  and (_04643_, _04642_, _04532_);
  and (_04644_, _04643_, _04530_);
  not (_04645_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_04646_, _04493_, _04247_);
  or (_04647_, _04646_, _04645_);
  and (_04648_, _04647_, _04644_);
  nand (_04649_, _04648_, _04495_);
  not (_04650_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_04651_, _04646_, _04650_);
  not (_04652_, _04644_);
  not (_04653_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_04654_, _04494_, _04653_);
  and (_04655_, _04654_, _04652_);
  nand (_04656_, _04655_, _04651_);
  nand (_04657_, _04656_, _04649_);
  nand (_04658_, _04657_, _04244_);
  not (_04659_, _04244_);
  not (_04660_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_04661_, _04646_, _04660_);
  not (_04662_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_04663_, _04494_, _04662_);
  and (_04664_, _04663_, _04652_);
  nand (_04665_, _04664_, _04661_);
  not (_04666_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_04667_, _04494_, _04666_);
  not (_04668_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_04669_, _04646_, _04668_);
  and (_04670_, _04669_, _04644_);
  nand (_04671_, _04670_, _04667_);
  nand (_04672_, _04671_, _04665_);
  nand (_04673_, _04672_, _04659_);
  nand (_04674_, _04673_, _04658_);
  nand (_04675_, _04674_, _04062_);
  not (_04676_, _04062_);
  nand (_04677_, _04494_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_04678_, _04646_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_04679_, _04678_, _04652_);
  nand (_04680_, _04679_, _04677_);
  not (_04681_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_04682_, _04494_, _04681_);
  nand (_04683_, _04494_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_04684_, _04683_, _04644_);
  nand (_04685_, _04684_, _04682_);
  nand (_04686_, _04685_, _04680_);
  nand (_04687_, _04686_, _04244_);
  nand (_04688_, _04494_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_04689_, _04646_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_04690_, _04689_, _04652_);
  nand (_04691_, _04690_, _04688_);
  nand (_04692_, _04646_, \oc8051_golden_model_1.IRAM[12] [0]);
  nand (_04693_, _04494_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_04694_, _04693_, _04644_);
  nand (_04695_, _04694_, _04692_);
  nand (_04696_, _04695_, _04691_);
  nand (_04697_, _04696_, _04659_);
  nand (_04698_, _04697_, _04687_);
  nand (_04699_, _04698_, _04676_);
  and (_04700_, _04699_, _04675_);
  and (_04701_, _04700_, _03771_);
  nor (_04702_, _03919_, _03378_);
  and (_04703_, _04702_, _04254_);
  nor (_04704_, _04703_, _03438_);
  not (_04705_, _04704_);
  nor (_04706_, _04705_, _04701_);
  and (_04707_, _03910_, _03766_);
  not (_04708_, _04707_);
  nor (_04709_, _04708_, _03647_);
  and (_04710_, _04709_, _03715_);
  nor (_04711_, _04710_, _04706_);
  and (_04712_, _04711_, _03770_);
  nor (_04713_, _04712_, _03769_);
  and (_04714_, _04421_, _03762_);
  nor (_04715_, _04714_, _04713_);
  and (_04716_, _03736_, _03762_);
  not (_04717_, _04716_);
  nor (_04718_, _04717_, _04700_);
  not (_04719_, _04718_);
  and (_04720_, _04719_, _04715_);
  nor (_04721_, _03764_, _03647_);
  not (_04722_, _03850_);
  nor (_04723_, _04722_, _03647_);
  and (_04724_, _04723_, _03715_);
  nor (_04725_, _04724_, _04721_);
  and (_04726_, _04725_, _04720_);
  not (_04727_, _04726_);
  and (_04728_, _04727_, _03765_);
  nor (_04729_, _03431_, _03683_);
  nor (_04730_, _04729_, _04728_);
  and (_04732_, _04421_, _03757_);
  not (_04733_, _03848_);
  nor (_04734_, _04733_, _03647_);
  and (_04735_, _04734_, _03715_);
  nor (_04736_, _04735_, _04732_);
  and (_04737_, _04736_, _04730_);
  and (_04738_, _03736_, _03757_);
  not (_04739_, _04738_);
  nor (_04740_, _04739_, _04700_);
  not (_04741_, _04740_);
  and (_04742_, _04741_, _04737_);
  nor (_04743_, _03760_, _03647_);
  nor (_04744_, _03855_, _03647_);
  and (_04745_, _04744_, _03715_);
  nor (_04746_, _04745_, _04743_);
  and (_04747_, _04746_, _04742_);
  nor (_04748_, _04747_, _03761_);
  or (_04749_, _04748_, _03758_);
  nand (_04750_, _03758_, _03683_);
  nand (_04751_, _04750_, _04749_);
  and (_04752_, _04751_, _03756_);
  nor (_04753_, _04752_, _03754_);
  or (_04754_, _03832_, _03824_);
  and (_04755_, _04422_, _03821_);
  or (_04756_, _04755_, _04754_);
  nor (_04757_, _04756_, _04753_);
  and (_04758_, _04757_, _03750_);
  nor (_04759_, _03747_, _03647_);
  and (_04760_, _03453_, _03422_);
  and (_04761_, _04760_, _03821_);
  nor (_04762_, _04761_, _04320_);
  nor (_04763_, _04762_, _04700_);
  nor (_04764_, _04763_, _04759_);
  and (_04765_, _04764_, _04758_);
  nor (_04766_, _04765_, _03748_);
  nor (_04767_, _04766_, _03456_);
  and (_04768_, _03456_, _03683_);
  nor (_04769_, _04768_, _04767_);
  and (_04770_, _04421_, _03400_);
  or (_04771_, _04770_, _04769_);
  nor (_04772_, _04771_, _03743_);
  and (_04773_, _03736_, _03400_);
  not (_04774_, _04773_);
  nor (_04775_, _04774_, _04700_);
  not (_04776_, _04775_);
  and (_04777_, _04776_, _04772_);
  not (_04778_, _03903_);
  nor (_04779_, _04778_, _03647_);
  and (_04780_, _04779_, _03715_);
  nor (_04781_, _04780_, _03401_);
  and (_04782_, _04781_, _04777_);
  and (_04783_, _03401_, _03683_);
  nor (_04784_, _04783_, _04782_);
  not (_04785_, _04027_);
  nor (_04786_, _04785_, _03647_);
  not (_04787_, _04786_);
  nor (_04788_, _03909_, _03647_);
  not (_04789_, _04788_);
  not (_04790_, _03897_);
  nor (_04791_, _04790_, _03647_);
  not (_04792_, _04018_);
  nor (_04793_, _04792_, _03647_);
  nor (_04794_, _04793_, _04791_);
  and (_04795_, _04794_, _04789_);
  and (_04796_, _04795_, _04787_);
  nor (_04797_, _04796_, _03716_);
  nor (_04798_, _04797_, _03388_);
  not (_04799_, _04798_);
  nor (_04800_, _04799_, _04784_);
  and (_04801_, _03388_, _03683_);
  nor (_04802_, _04801_, _04800_);
  nor (_04803_, _04012_, _03647_);
  and (_04804_, _04803_, _03715_);
  nor (_04805_, _04804_, _03383_);
  not (_04806_, _04805_);
  nor (_04807_, _04806_, _04802_);
  nor (_04808_, _04807_, _03684_);
  and (_04809_, _04421_, _03244_);
  nor (_04810_, _04809_, _04808_);
  nor (_04811_, _03774_, _03647_);
  and (_04812_, _03736_, _03244_);
  not (_04813_, _04812_);
  nor (_04814_, _04813_, _04700_);
  nor (_04815_, _04814_, _04811_);
  and (_04816_, _04815_, _04810_);
  and (_04817_, _04811_, _03716_);
  nor (_04818_, _04817_, _04816_);
  nor (_04819_, _03899_, _03414_);
  nor (_04820_, _04819_, _03683_);
  nor (_04821_, _04820_, _04818_);
  and (_04822_, _04821_, _03682_);
  nor (_04823_, _04822_, _03680_);
  and (_04824_, _04421_, _03412_);
  nor (_04825_, _04824_, _04823_);
  and (_04826_, _03736_, _03412_);
  not (_04827_, _04826_);
  nor (_04828_, _04827_, _04700_);
  not (_04829_, _04828_);
  and (_04830_, _04829_, _04825_);
  nor (_04831_, _04060_, _03647_);
  and (_04832_, _04831_, _03715_);
  not (_04833_, _04832_);
  and (_04834_, _04833_, _04830_);
  not (_04835_, _04563_);
  and (_04836_, _04831_, _04835_);
  and (_04837_, _04605_, \oc8051_golden_model_1.SP [0]);
  and (_04838_, \oc8051_golden_model_1.SP [1], _03683_);
  nor (_04839_, _04838_, _04837_);
  not (_04840_, _04839_);
  and (_04841_, _04840_, _03383_);
  and (_04842_, _04779_, _04835_);
  and (_04843_, _04527_, _03746_);
  and (_04844_, _04840_, _03758_);
  not (_04845_, _03758_);
  and (_04846_, _04723_, _04835_);
  and (_04847_, _03736_, _04261_);
  not (_04848_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_04849_, _04494_, _04848_);
  not (_04850_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_04851_, _04646_, _04850_);
  and (_04852_, _04851_, _04644_);
  nand (_04853_, _04852_, _04849_);
  not (_04854_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_04855_, _04646_, _04854_);
  not (_04856_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_04857_, _04494_, _04856_);
  and (_04858_, _04857_, _04652_);
  nand (_04859_, _04858_, _04855_);
  nand (_04860_, _04859_, _04853_);
  nand (_04861_, _04860_, _04244_);
  not (_04862_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_04863_, _04646_, _04862_);
  not (_04864_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_04865_, _04494_, _04864_);
  and (_04866_, _04865_, _04652_);
  nand (_04867_, _04866_, _04863_);
  not (_04868_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_04869_, _04494_, _04868_);
  not (_04870_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_04871_, _04646_, _04870_);
  and (_04872_, _04871_, _04644_);
  nand (_04873_, _04872_, _04869_);
  nand (_04874_, _04873_, _04867_);
  nand (_04875_, _04874_, _04659_);
  nand (_04876_, _04875_, _04861_);
  nand (_04877_, _04876_, _04062_);
  nand (_04878_, _04494_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_04879_, _04646_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_04880_, _04879_, _04652_);
  nand (_04881_, _04880_, _04878_);
  nand (_04882_, _04646_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_04883_, _04494_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_04884_, _04883_, _04644_);
  nand (_04885_, _04884_, _04882_);
  nand (_04886_, _04885_, _04881_);
  nand (_04887_, _04886_, _04244_);
  nand (_04888_, _04494_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_04889_, _04646_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_04890_, _04889_, _04652_);
  nand (_04891_, _04890_, _04888_);
  nand (_04892_, _04646_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_04893_, _04494_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_04894_, _04893_, _04644_);
  nand (_04895_, _04894_, _04892_);
  nand (_04896_, _04895_, _04891_);
  nand (_04897_, _04896_, _04659_);
  nand (_04898_, _04897_, _04887_);
  nand (_04899_, _04898_, _04676_);
  and (_04900_, _04899_, _04877_);
  nor (_04901_, _04900_, _03439_);
  or (_04902_, _04901_, _04847_);
  and (_04903_, _04709_, _04563_);
  or (_04904_, _04903_, _04902_);
  and (_04905_, _04839_, _03768_);
  and (_04906_, _03718_, _03762_);
  nor (_04907_, _04906_, _04905_);
  not (_04908_, _04907_);
  nor (_04909_, _04908_, _04904_);
  nor (_04910_, _04900_, _04717_);
  nor (_04911_, _04910_, _04723_);
  and (_04912_, _04911_, _04909_);
  nor (_04913_, _04912_, _04846_);
  and (_04914_, _04526_, _04721_);
  or (_04915_, _04914_, _04913_);
  nor (_04916_, _04840_, _03431_);
  or (_04917_, _04916_, _04915_);
  and (_04918_, _04734_, _04563_);
  and (_04919_, _03718_, _03757_);
  nor (_04920_, _04919_, _04918_);
  not (_04921_, _04920_);
  nor (_04922_, _04921_, _04917_);
  nor (_04923_, _04900_, _04739_);
  nor (_04924_, _04923_, _04744_);
  and (_04925_, _04924_, _04922_);
  and (_04926_, _04744_, _04835_);
  nor (_04927_, _04926_, _04925_);
  and (_04928_, _04526_, _04743_);
  nor (_04929_, _04928_, _04927_);
  and (_04930_, _04929_, _04845_);
  nor (_04931_, _04930_, _04844_);
  and (_04932_, _03755_, _04526_);
  or (_04933_, _04932_, _04931_);
  and (_04934_, _03718_, _03821_);
  nor (_04935_, _04840_, _03428_);
  nor (_04936_, _04935_, _04934_);
  not (_04937_, _04936_);
  nor (_04938_, _04937_, _04933_);
  and (_04939_, _03736_, _03821_);
  not (_04940_, _04939_);
  nor (_04941_, _04900_, _04940_);
  nor (_04942_, _04941_, _04759_);
  and (_04943_, _04942_, _04938_);
  nor (_04944_, _04943_, _04843_);
  nor (_04945_, _04944_, _03456_);
  and (_04946_, _04840_, _03456_);
  nor (_04947_, _04946_, _04945_);
  nor (_04948_, _03742_, _04835_);
  and (_04949_, _03718_, _03400_);
  nor (_04950_, _04949_, _04948_);
  not (_04951_, _04950_);
  nor (_04952_, _04951_, _04947_);
  nor (_04953_, _04900_, _04774_);
  nor (_04954_, _04953_, _04779_);
  and (_04955_, _04954_, _04952_);
  nor (_04956_, _04955_, _04842_);
  nor (_04957_, _04956_, _03401_);
  and (_04958_, _04840_, _03401_);
  nor (_04959_, _04958_, _04957_);
  nor (_04960_, _04796_, _04835_);
  nor (_04961_, _04960_, _03388_);
  not (_04962_, _04961_);
  nor (_04963_, _04962_, _04959_);
  and (_04964_, _04840_, _03388_);
  nor (_04965_, _04964_, _04963_);
  and (_04966_, _04803_, _04563_);
  nor (_04967_, _04966_, _03383_);
  not (_04968_, _04967_);
  nor (_04969_, _04968_, _04965_);
  nor (_04970_, _04969_, _04841_);
  and (_04971_, _03718_, _03244_);
  nor (_04972_, _04971_, _04970_);
  nor (_04973_, _04900_, _04813_);
  nor (_04974_, _04973_, _04811_);
  and (_04975_, _04974_, _04972_);
  and (_04976_, _04811_, _04835_);
  nor (_04977_, _04976_, _04975_);
  nor (_04978_, _04840_, _04819_);
  nor (_04979_, _04978_, _04977_);
  and (_04980_, _04979_, _03682_);
  nor (_04981_, _04980_, _04531_);
  and (_04982_, _03719_, _03412_);
  nor (_04983_, _04982_, _04199_);
  not (_04984_, _04983_);
  nor (_04985_, _04984_, _04981_);
  nor (_04986_, _04900_, _04827_);
  nor (_04987_, _04986_, _04831_);
  and (_04988_, _04987_, _04985_);
  nor (_04989_, _04988_, _04836_);
  not (_04990_, _00000_);
  nor (_04991_, _04723_, _04709_);
  nor (_04992_, _04803_, _03739_);
  and (_04993_, _04992_, _04991_);
  nor (_04994_, _04779_, _04721_);
  nor (_04995_, _03755_, _04734_);
  and (_04996_, _04995_, _04994_);
  and (_04997_, _04996_, _04993_);
  and (_04998_, _04997_, _04795_);
  nor (_04999_, _03740_, _03727_);
  nor (_05000_, _03733_, _03722_);
  and (_05001_, _05000_, _04999_);
  nor (_05002_, _04831_, _03681_);
  nor (_05003_, _04786_, _04744_);
  and (_05004_, _05003_, _05002_);
  not (_05005_, _04743_);
  not (_05006_, _03454_);
  nand (_05007_, _04702_, _05006_);
  and (_05008_, _05007_, _04261_);
  nor (_05009_, _03719_, _03736_);
  nor (_05010_, _05009_, _03438_);
  or (_05011_, _05010_, _05008_);
  not (_05012_, _05011_);
  and (_05013_, _04265_, _03307_);
  nor (_05014_, _05013_, _03827_);
  not (_05015_, _03308_);
  and (_05016_, _03728_, _03400_);
  and (_05017_, _05016_, _05015_);
  and (_05018_, _04485_, _03451_);
  nor (_05019_, _05018_, _05017_);
  and (_05020_, _05019_, _05014_);
  nor (_05021_, _04287_, _03768_);
  and (_05022_, _04282_, _05015_);
  not (_05023_, _05022_);
  and (_05024_, _05023_, _04631_);
  and (_05025_, _05024_, _05021_);
  and (_05026_, _05025_, _05020_);
  and (_05027_, _05026_, _05012_);
  and (_05028_, _04202_, _03838_);
  nor (_05029_, _04227_, _03832_);
  and (_05030_, _05029_, _04717_);
  and (_05031_, _03910_, _03400_);
  nor (_05032_, _05031_, _04228_);
  and (_05033_, _03831_, _03400_);
  nor (_05034_, _05033_, _04738_);
  and (_05035_, _05034_, _05032_);
  and (_05036_, _05035_, _05030_);
  and (_05037_, _03831_, _03412_);
  nor (_05038_, _04826_, _05037_);
  and (_05039_, _04422_, _03400_);
  and (_05040_, _03767_, _03400_);
  or (_05041_, _05040_, _05039_);
  not (_05042_, _05041_);
  and (_05043_, _05042_, _05038_);
  and (_05044_, _05043_, _05036_);
  not (_05045_, _03431_);
  nor (_05046_, _05045_, _03401_);
  and (_05047_, _05046_, _04819_);
  nor (_05048_, _03388_, _03383_);
  not (_05049_, _03428_);
  nor (_05050_, _03456_, _05049_);
  and (_05051_, _05050_, _05048_);
  and (_05052_, _05051_, _05047_);
  and (_05053_, _03719_, _03244_);
  nor (_05054_, _05053_, _04632_);
  nor (_05055_, _04939_, _03829_);
  and (_05056_, _05055_, _05054_);
  nor (_05057_, _04812_, _03758_);
  nor (_05058_, _04773_, _04188_);
  and (_05059_, _05058_, _05057_);
  and (_05060_, _05059_, _05056_);
  and (_05061_, _05060_, _05052_);
  and (_05062_, _05061_, _05044_);
  and (_05063_, _05062_, _05028_);
  and (_05064_, _05063_, _05027_);
  and (_05065_, _05064_, _05005_);
  nor (_05066_, _04811_, _04759_);
  and (_05067_, _05066_, _05065_);
  and (_05068_, _05067_, _05004_);
  and (_05069_, _05068_, _05001_);
  and (_05070_, _05069_, _04998_);
  nor (_05071_, _05070_, _04990_);
  not (_05072_, _05071_);
  nor (_05073_, _05072_, _04989_);
  and (_05074_, _05073_, _04834_);
  and (_05075_, _04646_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_05076_, _04494_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_05077_, _05076_, _05075_);
  and (_05078_, _05077_, _04644_);
  and (_05079_, _04494_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_05080_, _04646_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_05081_, _05080_, _05079_);
  and (_05082_, _05081_, _04652_);
  or (_05083_, _05082_, _05078_);
  nor (_05084_, _05083_, _04659_);
  and (_05085_, _04646_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_05086_, _04494_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_05087_, _05086_, _05085_);
  and (_05088_, _05087_, _04644_);
  and (_05089_, _04494_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_05090_, _04646_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_05091_, _05090_, _05089_);
  and (_05092_, _05091_, _04652_);
  or (_05093_, _05092_, _05088_);
  nor (_05094_, _05093_, _04244_);
  nor (_05095_, _05094_, _05084_);
  nor (_05096_, _05095_, _04676_);
  and (_05097_, _04646_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_05098_, _04494_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_05099_, _05098_, _05097_);
  and (_05100_, _05099_, _04644_);
  and (_05101_, _04494_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_05102_, _04646_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_05103_, _05102_, _05101_);
  and (_05104_, _05103_, _04652_);
  or (_05105_, _05104_, _05100_);
  nor (_05106_, _05105_, _04659_);
  and (_05107_, _04646_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_05108_, _04494_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_05109_, _05108_, _05107_);
  and (_05110_, _05109_, _04644_);
  and (_05111_, _04494_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_05112_, _04646_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_05113_, _05112_, _05111_);
  and (_05114_, _05113_, _04652_);
  or (_05115_, _05114_, _05110_);
  nor (_05116_, _05115_, _04244_);
  nor (_05117_, _05116_, _05106_);
  nor (_05118_, _05117_, _04062_);
  nor (_05119_, _05118_, _05096_);
  nor (_05120_, _05119_, _04813_);
  nor (_05121_, _05119_, _04774_);
  or (_05122_, _05119_, _04762_);
  and (_05123_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_05124_, _05123_, \oc8051_golden_model_1.SP [2]);
  nor (_05125_, _05124_, \oc8051_golden_model_1.SP [3]);
  and (_05126_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_05127_, _05126_, \oc8051_golden_model_1.SP [3]);
  and (_05128_, _05127_, \oc8051_golden_model_1.SP [0]);
  nor (_05129_, _05128_, _05125_);
  and (_05130_, _05129_, _05049_);
  not (_05131_, _04762_);
  not (_05132_, _04734_);
  and (_05133_, _05129_, _03768_);
  nor (_05134_, _05119_, _03439_);
  not (_05135_, \oc8051_golden_model_1.PSW [3]);
  and (_05136_, _03439_, _05135_);
  nor (_05137_, _05136_, _04709_);
  not (_05138_, _05137_);
  nor (_05139_, _05138_, _05134_);
  nor (_05140_, _04708_, _03679_);
  nor (_05141_, _05140_, _05139_);
  nor (_05142_, _05141_, _03768_);
  or (_05143_, _05142_, _04716_);
  nor (_05144_, _05143_, _05133_);
  nor (_05145_, _05119_, _04717_);
  nor (_05146_, _05145_, _04723_);
  not (_05147_, _05146_);
  nor (_05148_, _05147_, _05144_);
  nor (_05149_, _04722_, _03679_);
  or (_05150_, _05149_, _04721_);
  nor (_05151_, _05150_, _05148_);
  not (_05152_, _04721_);
  nor (_05153_, _05152_, _03811_);
  nor (_05154_, _05153_, _05151_);
  and (_05155_, _05154_, _03431_);
  and (_05156_, _05129_, _05045_);
  or (_05157_, _05156_, _05155_);
  and (_05158_, _05157_, _05132_);
  and (_05159_, _04734_, _03812_);
  nor (_05160_, _05159_, _04738_);
  not (_05161_, _05160_);
  nor (_05162_, _05161_, _05158_);
  nor (_05163_, _05119_, _04739_);
  nor (_05164_, _05163_, _04744_);
  not (_05165_, _05164_);
  nor (_05166_, _05165_, _05162_);
  and (_05167_, _04744_, _03812_);
  or (_05168_, _05167_, _04743_);
  nor (_05169_, _05168_, _05166_);
  and (_05170_, _03810_, _04743_);
  nor (_05171_, _05170_, _05169_);
  and (_05172_, _05171_, _04845_);
  and (_05173_, _05129_, _03758_);
  nor (_05174_, _05173_, _05172_);
  nor (_05175_, _05174_, _03755_);
  nor (_05176_, _03756_, _03814_);
  or (_05177_, _05176_, _05175_);
  and (_05178_, _05177_, _03428_);
  or (_05179_, _05178_, _05131_);
  nor (_05180_, _05179_, _05130_);
  nor (_05181_, _05180_, _04759_);
  and (_05182_, _05181_, _05122_);
  not (_05183_, _04759_);
  nor (_05184_, _05183_, _03814_);
  nor (_05185_, _05184_, _05182_);
  nor (_05186_, _05185_, _03456_);
  and (_05187_, _05129_, _03456_);
  not (_05188_, _05187_);
  and (_05189_, _05188_, _03742_);
  not (_05190_, _05189_);
  nor (_05191_, _05190_, _05186_);
  nor (_05192_, _03742_, _03812_);
  nor (_05193_, _05192_, _05191_);
  nor (_05194_, _05193_, _04773_);
  or (_05195_, _05194_, _04779_);
  nor (_05196_, _05195_, _05121_);
  and (_05197_, _04779_, _03812_);
  nor (_05198_, _05197_, _05196_);
  nor (_05199_, _05198_, _03401_);
  and (_05200_, _05129_, _03401_);
  not (_05201_, _05200_);
  and (_05202_, _05201_, _04796_);
  not (_05203_, _05202_);
  nor (_05204_, _05203_, _05199_);
  nor (_05205_, _04796_, _03812_);
  nor (_05206_, _05205_, _03388_);
  not (_05207_, _05206_);
  nor (_05208_, _05207_, _05204_);
  and (_05209_, _05129_, _03388_);
  nor (_05210_, _05209_, _04803_);
  not (_05211_, _05210_);
  nor (_05212_, _05211_, _05208_);
  and (_05213_, _04803_, _03678_);
  nor (_05214_, _05213_, _03383_);
  not (_05215_, _05214_);
  nor (_05216_, _05215_, _05212_);
  and (_05217_, _05129_, _03383_);
  nor (_05218_, _05217_, _04812_);
  not (_05219_, _05218_);
  nor (_05220_, _05219_, _05216_);
  or (_05221_, _05220_, _04811_);
  nor (_05222_, _05221_, _05120_);
  not (_05223_, _04819_);
  and (_05224_, _04811_, _03812_);
  nor (_05225_, _05224_, _05223_);
  not (_05226_, _05225_);
  nor (_05227_, _05226_, _05222_);
  nor (_05228_, _05129_, _04819_);
  nor (_05229_, _05228_, _03681_);
  not (_05230_, _05229_);
  nor (_05231_, _05230_, _05227_);
  not (_05232_, _03810_);
  and (_05233_, _03681_, _05232_);
  nor (_05234_, _05233_, _04826_);
  not (_05235_, _05234_);
  nor (_05236_, _05235_, _05231_);
  nor (_05237_, _05119_, _04827_);
  nor (_05238_, _05237_, _04831_);
  not (_05239_, _05238_);
  nor (_05240_, _05239_, _05236_);
  nor (_05241_, _04060_, _03679_);
  nor (_05242_, _05241_, _05240_);
  not (_05243_, _04139_);
  and (_05244_, _04831_, _05243_);
  not (_05245_, _05054_);
  nor (_05246_, _05123_, \oc8051_golden_model_1.SP [2]);
  nor (_05247_, _05246_, _05124_);
  and (_05248_, _05247_, _03383_);
  and (_05249_, _04779_, _05243_);
  nor (_05250_, _03742_, _05243_);
  and (_05251_, _04094_, _03746_);
  nor (_05252_, _05247_, _03428_);
  and (_05253_, _05247_, _03758_);
  and (_05254_, _04723_, _05243_);
  not (_05255_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_05256_, _04494_, _05255_);
  not (_05257_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_05258_, _04646_, _05257_);
  and (_05259_, _05258_, _04644_);
  nand (_05260_, _05259_, _05256_);
  not (_05261_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_05262_, _04646_, _05261_);
  not (_05263_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_05264_, _04494_, _05263_);
  and (_05265_, _05264_, _04652_);
  nand (_05266_, _05265_, _05262_);
  nand (_05267_, _05266_, _05260_);
  nand (_05268_, _05267_, _04244_);
  not (_05269_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_05270_, _04646_, _05269_);
  not (_05271_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_05272_, _04494_, _05271_);
  and (_05273_, _05272_, _04652_);
  nand (_05274_, _05273_, _05270_);
  not (_05275_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_05276_, _04494_, _05275_);
  not (_05277_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_05278_, _04646_, _05277_);
  and (_05279_, _05278_, _04644_);
  nand (_05280_, _05279_, _05276_);
  nand (_05281_, _05280_, _05274_);
  nand (_05282_, _05281_, _04659_);
  nand (_05283_, _05282_, _05268_);
  nand (_05284_, _05283_, _04062_);
  nand (_05285_, _04494_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_05286_, _04646_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_05287_, _05286_, _04652_);
  nand (_05288_, _05287_, _05285_);
  nand (_05289_, _04646_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_05290_, _04494_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_05291_, _05290_, _04644_);
  nand (_05292_, _05291_, _05289_);
  nand (_05293_, _05292_, _05288_);
  nand (_05294_, _05293_, _04244_);
  nand (_05295_, _04494_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_05296_, _04646_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_05297_, _05296_, _04652_);
  nand (_05298_, _05297_, _05295_);
  nand (_05299_, _04646_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_05300_, _04494_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_05301_, _05300_, _04644_);
  nand (_05302_, _05301_, _05299_);
  nand (_05303_, _05302_, _05298_);
  nand (_05304_, _05303_, _04659_);
  nand (_05305_, _05304_, _05294_);
  nand (_05306_, _05305_, _04676_);
  and (_05307_, _05306_, _05284_);
  nand (_05308_, _05307_, _03378_);
  and (_05309_, _05308_, _05008_);
  and (_05310_, _04709_, _04139_);
  or (_05311_, _05310_, _05309_);
  not (_05312_, _05247_);
  and (_05313_, _05312_, _03768_);
  nor (_05314_, _05313_, _04265_);
  not (_05315_, _05314_);
  nor (_05316_, _05315_, _05311_);
  nor (_05317_, _05307_, _04717_);
  nor (_05318_, _05317_, _04723_);
  and (_05319_, _05318_, _05316_);
  nor (_05320_, _05319_, _05254_);
  and (_05321_, _04721_, _04093_);
  or (_05322_, _05321_, _05320_);
  nor (_05323_, _05247_, _03431_);
  nor (_05324_, _05323_, _04734_);
  not (_05325_, _05324_);
  nor (_05326_, _05325_, _05322_);
  and (_05327_, _04734_, _05243_);
  nor (_05328_, _05327_, _05326_);
  nor (_05329_, _05328_, _04282_);
  nor (_05330_, _05307_, _04739_);
  nor (_05331_, _05330_, _04744_);
  and (_05332_, _05331_, _05329_);
  and (_05333_, _04744_, _05243_);
  nor (_05334_, _05333_, _05332_);
  and (_05335_, _04093_, _04743_);
  nor (_05336_, _05335_, _05334_);
  and (_05337_, _05336_, _04845_);
  nor (_05338_, _05337_, _05253_);
  and (_05339_, _03755_, _04093_);
  or (_05340_, _05339_, _05338_);
  and (_05341_, _03728_, _03821_);
  or (_05342_, _05341_, _05340_);
  nor (_05343_, _05342_, _05252_);
  nor (_05344_, _05307_, _04762_);
  nor (_05345_, _05344_, _04759_);
  and (_05346_, _05345_, _05343_);
  nor (_05347_, _05346_, _05251_);
  nor (_05348_, _05347_, _03456_);
  and (_05349_, _05247_, _03456_);
  nor (_05350_, _05349_, _05348_);
  or (_05351_, _05350_, _05016_);
  nor (_05352_, _05351_, _05250_);
  nor (_05353_, _05307_, _04774_);
  nor (_05354_, _05353_, _04779_);
  and (_05355_, _05354_, _05352_);
  nor (_05356_, _05355_, _05249_);
  nor (_05357_, _05356_, _03401_);
  and (_05358_, _05247_, _03401_);
  nor (_05359_, _05358_, _05357_);
  nor (_05360_, _04796_, _05243_);
  nor (_05361_, _05360_, _03388_);
  not (_05362_, _05361_);
  nor (_05363_, _05362_, _05359_);
  and (_05364_, _05247_, _03388_);
  nor (_05365_, _05364_, _05363_);
  and (_05366_, _04803_, _04139_);
  nor (_05367_, _05366_, _03383_);
  not (_05368_, _05367_);
  nor (_05369_, _05368_, _05365_);
  nor (_05370_, _05369_, _05248_);
  nor (_05371_, _05370_, _05245_);
  nor (_05372_, _05307_, _04813_);
  nor (_05373_, _05372_, _04811_);
  and (_05374_, _05373_, _05371_);
  and (_05375_, _04811_, _05243_);
  nor (_05376_, _05375_, _05374_);
  nor (_05377_, _05247_, _04819_);
  nor (_05378_, _05377_, _05376_);
  and (_05379_, _05378_, _03682_);
  nor (_05380_, _05379_, _04095_);
  nor (_05381_, _05380_, _04485_);
  nor (_05382_, _05307_, _04827_);
  nor (_05383_, _05382_, _04831_);
  and (_05384_, _05383_, _05381_);
  nor (_05385_, _05384_, _05244_);
  nor (_05386_, _05385_, _05072_);
  not (_05387_, _05386_);
  nor (_05388_, _05387_, _05242_);
  and (_05389_, _05388_, _05074_);
  or (_05390_, _05389_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_05391_, _05126_, _03683_);
  nor (_05392_, _05247_, _04838_);
  nor (_05393_, _05392_, _05391_);
  and (_05394_, _05127_, _03683_);
  nor (_05395_, _05391_, _05129_);
  nor (_05396_, _05395_, _05394_);
  and (_05397_, _44002_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_05398_, _05397_);
  and (_05399_, _05052_, _03770_);
  nor (_05400_, _05399_, _05398_);
  and (_05401_, _05400_, _05396_);
  and (_05402_, _05401_, _05393_);
  and (_05403_, _05402_, _04837_);
  not (_05404_, _05403_);
  and (_05405_, _05404_, _05390_);
  not (_05406_, _04989_);
  nor (_05407_, _05398_, _05070_);
  and (_05408_, _05407_, _04834_);
  and (_05409_, _05408_, _05406_);
  not (_05410_, _05385_);
  not (_05411_, _05407_);
  nor (_05412_, _05411_, _05242_);
  and (_05413_, _05412_, _05410_);
  and (_05414_, _05413_, _05409_);
  not (_05415_, _05414_);
  and (_05416_, _04139_, _03678_);
  and (_05417_, _04563_, _03715_);
  and (_05418_, _05417_, _05416_);
  not (_05419_, _04526_);
  and (_05420_, _05419_, _04093_);
  not (_05421_, _03647_);
  nor (_05422_, _03810_, _05421_);
  and (_05423_, _05422_, _05420_);
  and (_05424_, _05423_, _05418_);
  and (_05425_, _05424_, \oc8051_golden_model_1.PSW [7]);
  not (_05426_, _04093_);
  and (_05427_, _04526_, _05426_);
  and (_05428_, _05422_, _05427_);
  and (_05429_, _05428_, _05418_);
  and (_05430_, _05429_, \oc8051_golden_model_1.ACC [7]);
  nor (_05431_, _05430_, _05425_);
  and (_05432_, _05417_, _04139_);
  and (_05433_, _05432_, _03812_);
  and (_05434_, _03810_, _03647_);
  nor (_05435_, _04526_, _04093_);
  and (_05436_, _05435_, _05434_);
  and (_05437_, _05436_, _05433_);
  and (_05438_, _05437_, \oc8051_golden_model_1.IP [7]);
  and (_05439_, _05435_, _05422_);
  and (_05440_, _05439_, _05418_);
  and (_05441_, _05440_, \oc8051_golden_model_1.B [7]);
  nor (_05442_, _05441_, _05438_);
  and (_05443_, _05442_, _05431_);
  and (_05444_, _04526_, _04093_);
  nand (_05445_, _05444_, _05434_);
  not (_05446_, _05433_);
  nor (_05447_, _05446_, _05445_);
  and (_05448_, _05447_, \oc8051_golden_model_1.TCON [7]);
  nor (_05449_, _04139_, _03678_);
  nand (_05450_, _05449_, _05417_);
  nor (_05451_, _05450_, _05445_);
  and (_05452_, _05451_, \oc8051_golden_model_1.TH0 [7]);
  nor (_05453_, _05452_, _05448_);
  and (_05454_, _05420_, _05434_);
  and (_05455_, _05418_, _05454_);
  and (_05456_, _05455_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_05457_, _04563_, _03715_);
  not (_05458_, _05457_);
  nand (_05459_, _04139_, _03812_);
  or (_05460_, _05459_, _05458_);
  nor (_05461_, _05460_, _05445_);
  and (_05462_, _05461_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05463_, _05462_, _05456_);
  and (_05464_, _05463_, _05453_);
  and (_05465_, _05454_, _05433_);
  and (_05466_, _05465_, \oc8051_golden_model_1.SCON [7]);
  and (_05467_, _04563_, _03716_);
  nand (_05468_, _05449_, _05467_);
  nor (_05469_, _05468_, _05445_);
  and (_05470_, _05469_, \oc8051_golden_model_1.TH1 [7]);
  nor (_05471_, _05470_, _05466_);
  not (_05472_, _05467_);
  nor (_05473_, _05459_, _05472_);
  not (_05474_, _05473_);
  nor (_05475_, _05474_, _05445_);
  and (_05476_, _05475_, \oc8051_golden_model_1.TMOD [7]);
  nor (_05477_, _04563_, _03716_);
  not (_05478_, _05477_);
  or (_05479_, _05478_, _05459_);
  nor (_05480_, _05479_, _05445_);
  and (_05481_, _05480_, \oc8051_golden_model_1.TL0 [7]);
  nor (_05482_, _05481_, _05476_);
  and (_05483_, _05482_, _05471_);
  and (_05484_, _05483_, _05464_);
  and (_05485_, _05484_, _05443_);
  and (_05486_, _05457_, _05243_);
  nand (_05487_, _05486_, _03678_);
  nor (_05488_, _05487_, _05445_);
  and (_05489_, _05488_, \oc8051_golden_model_1.PCON [7]);
  not (_05490_, _05489_);
  and (_05491_, _05454_, _05473_);
  and (_05492_, _05491_, \oc8051_golden_model_1.SBUF [7]);
  and (_05493_, _05427_, _05434_);
  and (_05494_, _05493_, _05433_);
  and (_05495_, _05494_, \oc8051_golden_model_1.IE [7]);
  nor (_05496_, _05495_, _05492_);
  and (_05497_, _05496_, _05490_);
  and (_05498_, _05418_, _05493_);
  and (_05499_, _05498_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05500_, _05436_, _05418_);
  and (_05501_, _05500_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05502_, _05501_, _05499_);
  and (_05503_, _05502_, _05497_);
  not (_05504_, _05418_);
  nor (_05505_, _05504_, _05445_);
  and (_05506_, _05505_, \oc8051_golden_model_1.P0INREG [7]);
  not (_05507_, _05506_);
  nand (_05508_, _05457_, _05416_);
  nor (_05509_, _05508_, _05445_);
  and (_05510_, _05509_, \oc8051_golden_model_1.DPH [7]);
  not (_05511_, _05510_);
  nand (_05512_, _05477_, _05416_);
  nor (_05513_, _05512_, _05445_);
  and (_05514_, _05513_, \oc8051_golden_model_1.DPL [7]);
  nand (_05515_, _05467_, _05416_);
  nor (_05516_, _05515_, _05445_);
  and (_05517_, _05516_, \oc8051_golden_model_1.SP [7]);
  nor (_05518_, _05517_, _05514_);
  and (_05519_, _05518_, _05511_);
  and (_05520_, _05519_, _05507_);
  and (_05521_, _05520_, _05503_);
  and (_05522_, _05521_, _05485_);
  not (_05523_, _05522_);
  and (_05524_, _04646_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_05525_, _04494_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_05526_, _05525_, _05524_);
  and (_05527_, _05526_, _04644_);
  and (_05528_, _04494_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_05529_, _04646_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_05530_, _05529_, _05528_);
  and (_05531_, _05530_, _04652_);
  or (_05532_, _05531_, _05527_);
  nor (_05533_, _05532_, _04659_);
  and (_05534_, _04646_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_05535_, _04494_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_05536_, _05535_, _05534_);
  and (_05537_, _05536_, _04644_);
  and (_05538_, _04494_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_05539_, _04646_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_05540_, _05539_, _05538_);
  and (_05541_, _05540_, _04652_);
  or (_05542_, _05541_, _05537_);
  nor (_05543_, _05542_, _04244_);
  nor (_05544_, _05543_, _05533_);
  nor (_05545_, _05544_, _04676_);
  and (_05546_, _04646_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_05547_, _04494_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_05548_, _05547_, _05546_);
  and (_05549_, _05548_, _04644_);
  and (_05550_, _04494_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_05551_, _04646_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_05552_, _05551_, _05550_);
  and (_05553_, _05552_, _04652_);
  or (_05554_, _05553_, _05549_);
  nor (_05555_, _05554_, _04659_);
  and (_05556_, _04646_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_05557_, _04494_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_05558_, _05557_, _05556_);
  and (_05559_, _05558_, _04644_);
  and (_05560_, _04494_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_05561_, _04646_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_05562_, _05561_, _05560_);
  and (_05563_, _05562_, _04652_);
  or (_05564_, _05563_, _05559_);
  nor (_05565_, _05564_, _04244_);
  nor (_05566_, _05565_, _05555_);
  nor (_05567_, _05566_, _04062_);
  nor (_05568_, _05567_, _05545_);
  and (_05569_, _05568_, _05421_);
  nor (_05570_, _05569_, _05523_);
  not (_05571_, _05570_);
  and (_05572_, _05509_, \oc8051_golden_model_1.DPH [3]);
  and (_05573_, _05475_, \oc8051_golden_model_1.TMOD [3]);
  nor (_05574_, _05573_, _05572_);
  and (_05575_, _05447_, \oc8051_golden_model_1.TCON [3]);
  and (_05576_, _05465_, \oc8051_golden_model_1.SCON [3]);
  nor (_05577_, _05576_, _05575_);
  and (_05578_, _05577_, _05574_);
  and (_05579_, _05513_, \oc8051_golden_model_1.DPL [3]);
  and (_05580_, _05451_, \oc8051_golden_model_1.TH0 [3]);
  nor (_05581_, _05580_, _05579_);
  and (_05582_, _05516_, \oc8051_golden_model_1.SP [3]);
  and (_05583_, _05469_, \oc8051_golden_model_1.TH1 [3]);
  nor (_05584_, _05583_, _05582_);
  and (_05585_, _05584_, _05581_);
  nor (_05586_, _05459_, _05445_);
  and (_05587_, _05586_, _05457_);
  and (_05588_, _05587_, \oc8051_golden_model_1.TL1 [3]);
  and (_05589_, _05586_, _05477_);
  and (_05590_, _05589_, \oc8051_golden_model_1.TL0 [3]);
  nor (_05591_, _05590_, _05588_);
  and (_05592_, _05591_, _05585_);
  and (_05593_, _05592_, _05578_);
  and (_05594_, _05488_, \oc8051_golden_model_1.PCON [3]);
  not (_05595_, _05594_);
  and (_05596_, _05491_, \oc8051_golden_model_1.SBUF [3]);
  and (_05597_, _05494_, \oc8051_golden_model_1.IE [3]);
  nor (_05598_, _05597_, _05596_);
  and (_05599_, _05598_, _05595_);
  and (_05600_, _05424_, \oc8051_golden_model_1.PSW [3]);
  and (_05601_, _05440_, \oc8051_golden_model_1.B [3]);
  nor (_05602_, _05601_, _05600_);
  and (_05603_, _05437_, \oc8051_golden_model_1.IP [3]);
  and (_05604_, _05429_, \oc8051_golden_model_1.ACC [3]);
  nor (_05605_, _05604_, _05603_);
  and (_05606_, _05605_, _05602_);
  and (_05607_, _05505_, \oc8051_golden_model_1.P0INREG [3]);
  not (_05608_, _05607_);
  and (_05609_, _05455_, \oc8051_golden_model_1.P1INREG [3]);
  not (_05610_, _05609_);
  and (_05611_, _05498_, \oc8051_golden_model_1.P2INREG [3]);
  and (_05612_, _05500_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_05613_, _05612_, _05611_);
  and (_05614_, _05613_, _05610_);
  and (_05615_, _05614_, _05608_);
  and (_05616_, _05615_, _05606_);
  and (_05617_, _05616_, _05599_);
  and (_05618_, _05617_, _05593_);
  not (_05619_, _05618_);
  and (_05620_, _05119_, _05421_);
  nor (_05621_, _05620_, _05619_);
  not (_05622_, _05621_);
  and (_05623_, _05475_, \oc8051_golden_model_1.TMOD [1]);
  not (_05624_, _05623_);
  and (_05625_, _05465_, \oc8051_golden_model_1.SCON [1]);
  and (_05626_, _05491_, \oc8051_golden_model_1.SBUF [1]);
  nor (_05627_, _05626_, _05625_);
  and (_05628_, _05627_, _05624_);
  and (_05629_, _05451_, \oc8051_golden_model_1.TH0 [1]);
  and (_05630_, _05494_, \oc8051_golden_model_1.IE [1]);
  nor (_05631_, _05630_, _05629_);
  and (_05632_, _05509_, \oc8051_golden_model_1.DPH [1]);
  and (_05633_, _05469_, \oc8051_golden_model_1.TH1 [1]);
  nor (_05634_, _05633_, _05632_);
  and (_05635_, _05634_, _05631_);
  and (_05636_, _05589_, \oc8051_golden_model_1.TL0 [1]);
  and (_05637_, _05587_, \oc8051_golden_model_1.TL1 [1]);
  nor (_05638_, _05637_, _05636_);
  and (_05639_, _05638_, _05635_);
  and (_05640_, _05639_, _05628_);
  and (_05641_, _05513_, \oc8051_golden_model_1.DPL [1]);
  not (_05642_, _05641_);
  and (_05643_, _05516_, \oc8051_golden_model_1.SP [1]);
  and (_05644_, _05447_, \oc8051_golden_model_1.TCON [1]);
  nor (_05645_, _05644_, _05643_);
  and (_05646_, _05645_, _05642_);
  and (_05647_, _05424_, \oc8051_golden_model_1.PSW [1]);
  and (_05648_, _05440_, \oc8051_golden_model_1.B [1]);
  nor (_05649_, _05648_, _05647_);
  and (_05650_, _05437_, \oc8051_golden_model_1.IP [1]);
  and (_05651_, _05429_, \oc8051_golden_model_1.ACC [1]);
  nor (_05652_, _05651_, _05650_);
  and (_05653_, _05652_, _05649_);
  and (_05654_, _05488_, \oc8051_golden_model_1.PCON [1]);
  not (_05655_, _05654_);
  and (_05656_, _05498_, \oc8051_golden_model_1.P2INREG [1]);
  and (_05657_, _05500_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_05658_, _05657_, _05656_);
  and (_05659_, _05658_, _05655_);
  and (_05660_, _05505_, \oc8051_golden_model_1.P0INREG [1]);
  and (_05661_, _05455_, \oc8051_golden_model_1.P1INREG [1]);
  nor (_05662_, _05661_, _05660_);
  and (_05663_, _05662_, _05659_);
  and (_05664_, _05663_, _05653_);
  and (_05665_, _05664_, _05646_);
  and (_05666_, _05665_, _05640_);
  not (_05667_, _05666_);
  and (_05668_, _04900_, _05421_);
  nor (_05669_, _05668_, _05667_);
  and (_05670_, _05509_, \oc8051_golden_model_1.DPH [0]);
  and (_05671_, _05475_, \oc8051_golden_model_1.TMOD [0]);
  nor (_05672_, _05671_, _05670_);
  and (_05673_, _05447_, \oc8051_golden_model_1.TCON [0]);
  and (_05674_, _05465_, \oc8051_golden_model_1.SCON [0]);
  nor (_05675_, _05674_, _05673_);
  and (_05676_, _05675_, _05672_);
  and (_05677_, _05513_, \oc8051_golden_model_1.DPL [0]);
  and (_05678_, _05451_, \oc8051_golden_model_1.TH0 [0]);
  nor (_05679_, _05678_, _05677_);
  and (_05680_, _05516_, \oc8051_golden_model_1.SP [0]);
  and (_05681_, _05469_, \oc8051_golden_model_1.TH1 [0]);
  nor (_05682_, _05681_, _05680_);
  and (_05683_, _05682_, _05679_);
  and (_05684_, _05587_, \oc8051_golden_model_1.TL1 [0]);
  and (_05685_, _05589_, \oc8051_golden_model_1.TL0 [0]);
  nor (_05686_, _05685_, _05684_);
  and (_05687_, _05686_, _05683_);
  and (_05688_, _05687_, _05676_);
  and (_05689_, _05488_, \oc8051_golden_model_1.PCON [0]);
  not (_05690_, _05689_);
  and (_05691_, _05491_, \oc8051_golden_model_1.SBUF [0]);
  and (_05692_, _05494_, \oc8051_golden_model_1.IE [0]);
  nor (_05693_, _05692_, _05691_);
  and (_05694_, _05693_, _05690_);
  and (_05695_, _05437_, \oc8051_golden_model_1.IP [0]);
  and (_05696_, _05429_, \oc8051_golden_model_1.ACC [0]);
  nor (_05697_, _05696_, _05695_);
  and (_05698_, _05424_, \oc8051_golden_model_1.PSW [0]);
  and (_05699_, _05440_, \oc8051_golden_model_1.B [0]);
  nor (_05700_, _05699_, _05698_);
  and (_05701_, _05700_, _05697_);
  and (_05702_, _05505_, \oc8051_golden_model_1.P0INREG [0]);
  not (_05703_, _05702_);
  and (_05704_, _05455_, \oc8051_golden_model_1.P1INREG [0]);
  not (_05705_, _05704_);
  and (_05706_, _05498_, \oc8051_golden_model_1.P2INREG [0]);
  and (_05707_, _05500_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_05708_, _05707_, _05706_);
  and (_05709_, _05708_, _05705_);
  and (_05710_, _05709_, _05703_);
  and (_05711_, _05710_, _05701_);
  and (_05712_, _05711_, _05694_);
  and (_05713_, _05712_, _05688_);
  not (_05714_, _05713_);
  and (_05715_, _04700_, _05421_);
  nor (_05716_, _05715_, _05714_);
  nor (_05717_, _05716_, _05669_);
  and (_05718_, _05424_, \oc8051_golden_model_1.PSW [2]);
  and (_05719_, _05440_, \oc8051_golden_model_1.B [2]);
  nor (_05720_, _05719_, _05718_);
  and (_05721_, _05437_, \oc8051_golden_model_1.IP [2]);
  and (_05722_, _05429_, \oc8051_golden_model_1.ACC [2]);
  nor (_05723_, _05722_, _05721_);
  and (_05724_, _05723_, _05720_);
  and (_05725_, _05447_, \oc8051_golden_model_1.TCON [2]);
  and (_05726_, _05451_, \oc8051_golden_model_1.TH0 [2]);
  nor (_05727_, _05726_, _05725_);
  and (_05728_, _05455_, \oc8051_golden_model_1.P1INREG [2]);
  and (_05729_, _05461_, \oc8051_golden_model_1.TL1 [2]);
  nor (_05730_, _05729_, _05728_);
  and (_05731_, _05730_, _05727_);
  and (_05732_, _05465_, \oc8051_golden_model_1.SCON [2]);
  and (_05733_, _05469_, \oc8051_golden_model_1.TH1 [2]);
  nor (_05734_, _05733_, _05732_);
  and (_05735_, _05475_, \oc8051_golden_model_1.TMOD [2]);
  and (_05736_, _05480_, \oc8051_golden_model_1.TL0 [2]);
  nor (_05737_, _05736_, _05735_);
  and (_05738_, _05737_, _05734_);
  and (_05739_, _05738_, _05731_);
  and (_05740_, _05739_, _05724_);
  and (_05741_, _05488_, \oc8051_golden_model_1.PCON [2]);
  not (_05742_, _05741_);
  and (_05743_, _05491_, \oc8051_golden_model_1.SBUF [2]);
  and (_05744_, _05494_, \oc8051_golden_model_1.IE [2]);
  nor (_05745_, _05744_, _05743_);
  and (_05746_, _05745_, _05742_);
  and (_05747_, _05498_, \oc8051_golden_model_1.P2INREG [2]);
  and (_05748_, _05500_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_05749_, _05748_, _05747_);
  and (_05750_, _05749_, _05746_);
  and (_05751_, _05505_, \oc8051_golden_model_1.P0INREG [2]);
  not (_05752_, _05751_);
  and (_05753_, _05509_, \oc8051_golden_model_1.DPH [2]);
  not (_05754_, _05753_);
  and (_05755_, _05513_, \oc8051_golden_model_1.DPL [2]);
  and (_05756_, _05516_, \oc8051_golden_model_1.SP [2]);
  nor (_05757_, _05756_, _05755_);
  and (_05758_, _05757_, _05754_);
  and (_05759_, _05758_, _05752_);
  and (_05760_, _05759_, _05750_);
  and (_05761_, _05760_, _05740_);
  not (_05762_, _05761_);
  and (_05763_, _05307_, _05421_);
  nor (_05764_, _05763_, _05762_);
  not (_05765_, _05764_);
  and (_05766_, _05765_, _05717_);
  and (_05767_, _05766_, _05622_);
  and (_05768_, _05424_, \oc8051_golden_model_1.PSW [5]);
  and (_05769_, _05429_, \oc8051_golden_model_1.ACC [5]);
  nor (_05770_, _05769_, _05768_);
  and (_05771_, _05437_, \oc8051_golden_model_1.IP [5]);
  and (_05772_, _05440_, \oc8051_golden_model_1.B [5]);
  nor (_05773_, _05772_, _05771_);
  and (_05774_, _05773_, _05770_);
  and (_05775_, _05447_, \oc8051_golden_model_1.TCON [5]);
  and (_05776_, _05451_, \oc8051_golden_model_1.TH0 [5]);
  nor (_05777_, _05776_, _05775_);
  and (_05778_, _05455_, \oc8051_golden_model_1.P1INREG [5]);
  and (_05779_, _05461_, \oc8051_golden_model_1.TL1 [5]);
  nor (_05780_, _05779_, _05778_);
  and (_05781_, _05780_, _05777_);
  and (_05782_, _05465_, \oc8051_golden_model_1.SCON [5]);
  and (_05783_, _05469_, \oc8051_golden_model_1.TH1 [5]);
  nor (_05784_, _05783_, _05782_);
  and (_05785_, _05475_, \oc8051_golden_model_1.TMOD [5]);
  and (_05786_, _05480_, \oc8051_golden_model_1.TL0 [5]);
  nor (_05787_, _05786_, _05785_);
  and (_05788_, _05787_, _05784_);
  and (_05789_, _05788_, _05781_);
  and (_05790_, _05789_, _05774_);
  and (_05791_, _05488_, \oc8051_golden_model_1.PCON [5]);
  not (_05792_, _05791_);
  and (_05793_, _05491_, \oc8051_golden_model_1.SBUF [5]);
  and (_05794_, _05494_, \oc8051_golden_model_1.IE [5]);
  nor (_05795_, _05794_, _05793_);
  and (_05796_, _05795_, _05792_);
  and (_05797_, _05498_, \oc8051_golden_model_1.P2INREG [5]);
  and (_05798_, _05500_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_05799_, _05798_, _05797_);
  and (_05800_, _05799_, _05796_);
  and (_05801_, _05505_, \oc8051_golden_model_1.P0INREG [5]);
  not (_05802_, _05801_);
  and (_05803_, _05509_, \oc8051_golden_model_1.DPH [5]);
  not (_05804_, _05803_);
  and (_05805_, _05513_, \oc8051_golden_model_1.DPL [5]);
  and (_05806_, _05516_, \oc8051_golden_model_1.SP [5]);
  nor (_05807_, _05806_, _05805_);
  and (_05808_, _05807_, _05804_);
  and (_05809_, _05808_, _05802_);
  and (_05810_, _05809_, _05800_);
  and (_05811_, _05810_, _05790_);
  not (_05812_, _05811_);
  and (_05813_, _04646_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_05814_, _04494_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_05815_, _05814_, _05813_);
  and (_05816_, _05815_, _04644_);
  and (_05817_, _04494_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_05818_, _04646_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_05819_, _05818_, _05817_);
  and (_05820_, _05819_, _04652_);
  or (_05821_, _05820_, _05816_);
  nor (_05822_, _05821_, _04659_);
  and (_05823_, _04646_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_05824_, _04494_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_05825_, _05824_, _05823_);
  and (_05826_, _05825_, _04644_);
  and (_05827_, _04494_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_05828_, _04646_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_05829_, _05828_, _05827_);
  and (_05830_, _05829_, _04652_);
  or (_05831_, _05830_, _05826_);
  nor (_05832_, _05831_, _04244_);
  nor (_05833_, _05832_, _05822_);
  nor (_05834_, _05833_, _04676_);
  and (_05835_, _04646_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_05836_, _04494_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_05837_, _05836_, _05835_);
  and (_05838_, _05837_, _04644_);
  and (_05839_, _04494_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_05840_, _04646_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_05841_, _05840_, _05839_);
  and (_05842_, _05841_, _04652_);
  or (_05843_, _05842_, _05838_);
  nor (_05844_, _05843_, _04659_);
  and (_05845_, _04646_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_05846_, _04494_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_05847_, _05846_, _05845_);
  and (_05848_, _05847_, _04644_);
  and (_05849_, _04494_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_05850_, _04646_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_05851_, _05850_, _05849_);
  and (_05852_, _05851_, _04652_);
  or (_05853_, _05852_, _05848_);
  nor (_05854_, _05853_, _04244_);
  nor (_05855_, _05854_, _05844_);
  nor (_05856_, _05855_, _04062_);
  nor (_05857_, _05856_, _05834_);
  and (_05858_, _05857_, _05421_);
  nor (_05859_, _05858_, _05812_);
  and (_05860_, _05424_, \oc8051_golden_model_1.PSW [4]);
  and (_05861_, _05440_, \oc8051_golden_model_1.B [4]);
  nor (_05862_, _05861_, _05860_);
  and (_05863_, _05437_, \oc8051_golden_model_1.IP [4]);
  and (_05864_, _05429_, \oc8051_golden_model_1.ACC [4]);
  nor (_05865_, _05864_, _05863_);
  and (_05866_, _05865_, _05862_);
  and (_05867_, _05447_, \oc8051_golden_model_1.TCON [4]);
  and (_05868_, _05451_, \oc8051_golden_model_1.TH0 [4]);
  nor (_05869_, _05868_, _05867_);
  and (_05870_, _05455_, \oc8051_golden_model_1.P1INREG [4]);
  and (_05871_, _05461_, \oc8051_golden_model_1.TL1 [4]);
  nor (_05872_, _05871_, _05870_);
  and (_05873_, _05872_, _05869_);
  and (_05874_, _05465_, \oc8051_golden_model_1.SCON [4]);
  and (_05875_, _05469_, \oc8051_golden_model_1.TH1 [4]);
  nor (_05876_, _05875_, _05874_);
  and (_05877_, _05475_, \oc8051_golden_model_1.TMOD [4]);
  and (_05878_, _05480_, \oc8051_golden_model_1.TL0 [4]);
  nor (_05879_, _05878_, _05877_);
  and (_05880_, _05879_, _05876_);
  and (_05881_, _05880_, _05873_);
  and (_05882_, _05881_, _05866_);
  and (_05883_, _05488_, \oc8051_golden_model_1.PCON [4]);
  not (_05884_, _05883_);
  and (_05885_, _05491_, \oc8051_golden_model_1.SBUF [4]);
  and (_05886_, _05494_, \oc8051_golden_model_1.IE [4]);
  nor (_05887_, _05886_, _05885_);
  and (_05888_, _05887_, _05884_);
  and (_05889_, _05498_, \oc8051_golden_model_1.P2INREG [4]);
  and (_05890_, _05500_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_05891_, _05890_, _05889_);
  and (_05892_, _05891_, _05888_);
  and (_05893_, _05505_, \oc8051_golden_model_1.P0INREG [4]);
  not (_05894_, _05893_);
  and (_05895_, _05509_, \oc8051_golden_model_1.DPH [4]);
  not (_05896_, _05895_);
  and (_05897_, _05513_, \oc8051_golden_model_1.DPL [4]);
  and (_05898_, _05516_, \oc8051_golden_model_1.SP [4]);
  nor (_05899_, _05898_, _05897_);
  and (_05900_, _05899_, _05896_);
  and (_05901_, _05900_, _05894_);
  and (_05902_, _05901_, _05892_);
  and (_05903_, _05902_, _05882_);
  not (_05904_, _05903_);
  and (_05905_, _04646_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_05906_, _04494_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_05907_, _05906_, _05905_);
  and (_05908_, _05907_, _04644_);
  and (_05909_, _04494_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_05910_, _04646_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05911_, _05910_, _05909_);
  and (_05912_, _05911_, _04652_);
  or (_05913_, _05912_, _05908_);
  nor (_05914_, _05913_, _04659_);
  and (_05915_, _04646_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_05916_, _04494_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_05917_, _05916_, _05915_);
  and (_05918_, _05917_, _04644_);
  and (_05919_, _04494_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_05920_, _04646_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05921_, _05920_, _05919_);
  and (_05922_, _05921_, _04652_);
  or (_05923_, _05922_, _05918_);
  nor (_05924_, _05923_, _04244_);
  nor (_05925_, _05924_, _05914_);
  nor (_05926_, _05925_, _04676_);
  and (_05927_, _04646_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_05928_, _04494_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_05929_, _05928_, _05927_);
  and (_05930_, _05929_, _04644_);
  and (_05931_, _04494_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_05932_, _04646_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_05933_, _05932_, _05931_);
  and (_05934_, _05933_, _04652_);
  or (_05935_, _05934_, _05930_);
  nor (_05936_, _05935_, _04659_);
  and (_05937_, _04646_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_05938_, _04494_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_05939_, _05938_, _05937_);
  and (_05940_, _05939_, _04644_);
  and (_05941_, _04494_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_05942_, _04646_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_05943_, _05942_, _05941_);
  and (_05944_, _05943_, _04652_);
  or (_05945_, _05944_, _05940_);
  nor (_05946_, _05945_, _04244_);
  nor (_05947_, _05946_, _05936_);
  nor (_05949_, _05947_, _04062_);
  nor (_05950_, _05949_, _05926_);
  and (_05952_, _05950_, _05421_);
  nor (_05953_, _05952_, _05904_);
  nor (_05955_, _05953_, _05859_);
  and (_05956_, _05955_, _05767_);
  nor (_05958_, _05956_, _05571_);
  and (_05959_, _05437_, \oc8051_golden_model_1.IP [6]);
  and (_05961_, _05440_, \oc8051_golden_model_1.B [6]);
  nor (_05962_, _05961_, _05959_);
  and (_05964_, _05424_, \oc8051_golden_model_1.PSW [6]);
  and (_05965_, _05429_, \oc8051_golden_model_1.ACC [6]);
  nor (_05967_, _05965_, _05964_);
  and (_05968_, _05967_, _05962_);
  and (_05970_, _05447_, \oc8051_golden_model_1.TCON [6]);
  and (_05971_, _05451_, \oc8051_golden_model_1.TH0 [6]);
  nor (_05973_, _05971_, _05970_);
  and (_05974_, _05455_, \oc8051_golden_model_1.P1INREG [6]);
  and (_05976_, _05461_, \oc8051_golden_model_1.TL1 [6]);
  nor (_05977_, _05976_, _05974_);
  and (_05979_, _05977_, _05973_);
  and (_05980_, _05465_, \oc8051_golden_model_1.SCON [6]);
  and (_05982_, _05469_, \oc8051_golden_model_1.TH1 [6]);
  nor (_05983_, _05982_, _05980_);
  and (_05985_, _05475_, \oc8051_golden_model_1.TMOD [6]);
  and (_05986_, _05480_, \oc8051_golden_model_1.TL0 [6]);
  nor (_05987_, _05986_, _05985_);
  and (_05988_, _05987_, _05983_);
  and (_05989_, _05988_, _05979_);
  and (_05990_, _05989_, _05968_);
  and (_05991_, _05488_, \oc8051_golden_model_1.PCON [6]);
  not (_05992_, _05991_);
  and (_05993_, _05491_, \oc8051_golden_model_1.SBUF [6]);
  and (_05994_, _05494_, \oc8051_golden_model_1.IE [6]);
  nor (_05995_, _05994_, _05993_);
  and (_05996_, _05995_, _05992_);
  and (_05997_, _05498_, \oc8051_golden_model_1.P2INREG [6]);
  and (_05998_, _05500_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_05999_, _05998_, _05997_);
  and (_06000_, _05999_, _05996_);
  and (_06001_, _05505_, \oc8051_golden_model_1.P0INREG [6]);
  not (_06002_, _06001_);
  and (_06003_, _05509_, \oc8051_golden_model_1.DPH [6]);
  not (_06004_, _06003_);
  and (_06005_, _05513_, \oc8051_golden_model_1.DPL [6]);
  and (_06006_, _05516_, \oc8051_golden_model_1.SP [6]);
  nor (_06007_, _06006_, _06005_);
  and (_06008_, _06007_, _06004_);
  and (_06009_, _06008_, _06002_);
  and (_06010_, _06009_, _06000_);
  and (_06011_, _06010_, _05990_);
  not (_06012_, _06011_);
  and (_06013_, _04646_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_06014_, _04494_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_06015_, _06014_, _06013_);
  and (_06016_, _06015_, _04644_);
  nor (_06017_, _04646_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor (_06018_, _04494_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor (_06019_, _06018_, _06017_);
  and (_06020_, _06019_, _04652_);
  nor (_06021_, _06020_, _06016_);
  nor (_06022_, _06021_, _04659_);
  and (_06023_, _04646_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_06024_, _04494_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_06025_, _06024_, _06023_);
  and (_06026_, _06025_, _04644_);
  nor (_06027_, _04646_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_06028_, _04494_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_06029_, _06028_, _06027_);
  and (_06030_, _06029_, _04652_);
  nor (_06031_, _06030_, _06026_);
  nor (_06032_, _06031_, _04244_);
  or (_06033_, _06032_, _06022_);
  nor (_06034_, _06033_, _04062_);
  and (_06035_, _04646_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_06036_, _04494_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_06037_, _06036_, _06035_);
  and (_06038_, _06037_, _04644_);
  and (_06039_, _04494_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_06040_, _04646_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_06041_, _06040_, _06039_);
  and (_06042_, _06041_, _04652_);
  or (_06044_, _06042_, _06038_);
  nor (_06046_, _06044_, _04659_);
  and (_06047_, _04646_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_06049_, _04494_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_06050_, _06049_, _06047_);
  and (_06052_, _06050_, _04644_);
  and (_06053_, _04494_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_06055_, _04646_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_06056_, _06055_, _06053_);
  and (_06058_, _06056_, _04652_);
  or (_06059_, _06058_, _06052_);
  nor (_06061_, _06059_, _04244_);
  nor (_06062_, _06061_, _06046_);
  nor (_06064_, _06062_, _04676_);
  nor (_06065_, _06064_, _06034_);
  and (_06067_, _06065_, _05421_);
  nor (_06068_, _06067_, _06012_);
  and (_06070_, _06068_, _05570_);
  nor (_06071_, _06068_, _05570_);
  nor (_06073_, _06071_, _06070_);
  not (_06074_, _06073_);
  and (_06076_, _06074_, _05956_);
  nor (_06077_, _06076_, _05958_);
  and (_06078_, _06077_, _04831_);
  not (_06079_, _05569_);
  not (_06080_, _03814_);
  nor (_06081_, _04527_, _04094_);
  and (_06082_, _06081_, _03679_);
  and (_06083_, _06082_, _06080_);
  not (_06084_, _06083_);
  nor (_06085_, _06084_, _05445_);
  and (_06086_, _06085_, \oc8051_golden_model_1.TCON [7]);
  and (_06087_, _06082_, _03814_);
  and (_06088_, _06087_, _05439_);
  and (_06089_, _06088_, \oc8051_golden_model_1.B [7]);
  nor (_06090_, _06089_, _06086_);
  and (_06091_, _06083_, _05436_);
  and (_06092_, _06091_, \oc8051_golden_model_1.IP [7]);
  not (_06093_, _06092_);
  and (_06094_, _06087_, _05423_);
  and (_06095_, _06094_, \oc8051_golden_model_1.PSW [7]);
  and (_06096_, _06087_, _05428_);
  and (_06097_, _06096_, \oc8051_golden_model_1.ACC [7]);
  nor (_06098_, _06097_, _06095_);
  and (_06099_, _06098_, _06093_);
  and (_06100_, _06099_, _06090_);
  and (_06101_, _06083_, _05454_);
  and (_06102_, _06101_, \oc8051_golden_model_1.SCON [7]);
  and (_06103_, _06083_, _05493_);
  and (_06104_, _06103_, \oc8051_golden_model_1.IE [7]);
  nor (_06105_, _06104_, _06102_);
  and (_06106_, _06087_, _05493_);
  and (_06107_, _06106_, \oc8051_golden_model_1.P2INREG [7]);
  and (_06108_, _06087_, _05436_);
  and (_06109_, _06108_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06110_, _06109_, _06107_);
  not (_06111_, _06087_);
  nor (_06112_, _06111_, _05445_);
  and (_06113_, _06112_, \oc8051_golden_model_1.P0INREG [7]);
  and (_06114_, _06087_, _05454_);
  and (_06115_, _06114_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_06116_, _06115_, _06113_);
  and (_06117_, _06116_, _06110_);
  and (_06118_, _06117_, _06105_);
  and (_06119_, _06118_, _06100_);
  and (_06120_, _06119_, _06079_);
  nor (_06121_, _06120_, _05486_);
  and (_06122_, _06121_, _03681_);
  not (_06123_, _06065_);
  nor (_06124_, _05950_, _05857_);
  nor (_06125_, _04900_, _04700_);
  nor (_06126_, _05307_, _05119_);
  and (_06127_, _06126_, _06125_);
  and (_06128_, _06127_, _06124_);
  and (_06129_, _06128_, _06123_);
  or (_06130_, _06129_, _05568_);
  nand (_06131_, _06129_, _05568_);
  and (_06132_, _06131_, _06130_);
  and (_06133_, _06132_, _05053_);
  or (_06134_, _06133_, _04812_);
  not (_06135_, _05016_);
  nor (_06136_, _05031_, _04773_);
  and (_06137_, _06136_, _06135_);
  and (_06138_, _06137_, _05042_);
  and (_06139_, _06138_, _04778_);
  or (_06140_, _06139_, _03647_);
  not (_06141_, _03456_);
  and (_06142_, _05486_, \oc8051_golden_model_1.PSW [7]);
  nor (_06143_, _06142_, _06121_);
  nor (_06144_, _06143_, _05183_);
  not (_06145_, _05486_);
  nor (_06146_, _06120_, _06145_);
  not (_06147_, _06146_);
  nand (_06148_, _06120_, _06145_);
  and (_06149_, _06148_, _06147_);
  and (_06150_, _06149_, _03755_);
  or (_06151_, _06121_, _05005_);
  and (_06152_, _05953_, _05859_);
  and (_06153_, _05716_, _05669_);
  and (_06154_, _05764_, _05621_);
  and (_06155_, _06154_, _06153_);
  and (_06156_, _06155_, _06152_);
  and (_06157_, _06156_, _06068_);
  nor (_06158_, _06157_, _05571_);
  and (_06159_, _06157_, _05571_);
  nor (_06160_, _06159_, _06158_);
  and (_06161_, _06160_, _04723_);
  nor (_06162_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_06163_, _06162_, _04182_);
  nor (_06164_, _06163_, _03847_);
  nor (_06165_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_06166_, _06165_, _03847_);
  and (_06167_, _06166_, _03683_);
  nor (_06168_, _06167_, _06164_);
  nor (_06169_, _06168_, _04183_);
  not (_06170_, _06169_);
  nor (_06171_, _05119_, _04939_);
  not (_06172_, _04183_);
  and (_06173_, _04939_, _03678_);
  or (_06174_, _06173_, _06172_);
  or (_06175_, _06174_, _06171_);
  and (_06176_, _06175_, _06170_);
  nor (_06177_, _06162_, _04182_);
  nor (_06178_, _06177_, _06163_);
  nor (_06179_, _06178_, _04183_);
  not (_06180_, _06179_);
  or (_06181_, _05307_, _05131_);
  nand (_06182_, _04939_, _04139_);
  and (_06183_, _06182_, _04183_);
  nand (_06184_, _06183_, _06181_);
  and (_06185_, _06184_, _06180_);
  not (_06186_, _06185_);
  nor (_06187_, _04839_, _04183_);
  not (_06188_, _06187_);
  and (_06189_, _04900_, _04940_);
  nor (_06190_, _04940_, _04563_);
  or (_06191_, _06190_, _06172_);
  or (_06192_, _06191_, _06189_);
  nand (_06193_, _06192_, _06188_);
  or (_06194_, _05131_, _04700_);
  and (_06195_, _04939_, _03715_);
  nor (_06196_, _06195_, _06172_);
  nand (_06197_, _06196_, _06194_);
  nor (_06198_, _04183_, \oc8051_golden_model_1.SP [0]);
  not (_06199_, _06198_);
  and (_06200_, _06199_, _06197_);
  and (_06201_, _06200_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_06202_, _06199_, _06197_);
  and (_06203_, _06202_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_06204_, _06203_, _06201_);
  and (_06205_, _06204_, _06193_);
  and (_06206_, _06192_, _06188_);
  and (_06207_, _06200_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_06208_, _06202_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_06209_, _06208_, _06207_);
  and (_06210_, _06209_, _06206_);
  or (_06211_, _06210_, _06205_);
  nor (_06212_, _06211_, _06186_);
  and (_06213_, _06200_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_06214_, _06202_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_06215_, _06214_, _06213_);
  and (_06216_, _06215_, _06193_);
  and (_06217_, _06200_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_06218_, _06202_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_06219_, _06218_, _06217_);
  and (_06220_, _06219_, _06206_);
  or (_06221_, _06220_, _06216_);
  nor (_06222_, _06221_, _06185_);
  nor (_06223_, _06222_, _06212_);
  nor (_06224_, _06223_, _06176_);
  not (_06225_, _06176_);
  and (_06226_, _06202_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_06227_, _06200_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_06228_, _06227_, _06226_);
  and (_06229_, _06228_, _06193_);
  and (_06230_, _06200_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_06231_, _06202_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_06232_, _06231_, _06230_);
  and (_06233_, _06232_, _06206_);
  or (_06234_, _06233_, _06229_);
  nor (_06235_, _06234_, _06186_);
  and (_06236_, _06200_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_06237_, _06202_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_06238_, _06237_, _06236_);
  and (_06239_, _06238_, _06193_);
  and (_06240_, _06200_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_06241_, _06202_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_06242_, _06241_, _06240_);
  and (_06243_, _06242_, _06206_);
  or (_06244_, _06243_, _06239_);
  nor (_06245_, _06244_, _06185_);
  nor (_06246_, _06245_, _06235_);
  nor (_06247_, _06246_, _06225_);
  nor (_06248_, _06247_, _06224_);
  or (_06249_, _06248_, _04717_);
  not (_06250_, _04723_);
  and (_06251_, _06132_, _04267_);
  and (_06252_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_06253_, _06252_, \oc8051_golden_model_1.PC [6]);
  and (_06254_, _06253_, _03550_);
  and (_06255_, _06254_, \oc8051_golden_model_1.PC [7]);
  nor (_06256_, _06254_, \oc8051_golden_model_1.PC [7]);
  nor (_06257_, _06256_, _06255_);
  not (_06258_, _06257_);
  nand (_06259_, _06258_, _03768_);
  or (_06260_, _03768_, \oc8051_golden_model_1.ACC [7]);
  and (_06261_, _06260_, _06259_);
  and (_06262_, _06261_, _04266_);
  or (_06263_, _06262_, _04716_);
  or (_06264_, _06263_, _06251_);
  and (_06265_, _06264_, _06250_);
  and (_06266_, _06265_, _06249_);
  or (_06267_, _06266_, _06161_);
  and (_06268_, _06267_, _05152_);
  and (_06269_, _06148_, _04721_);
  or (_06270_, _06269_, _05045_);
  or (_06271_, _06270_, _06268_);
  nor (_06272_, _06257_, _03431_);
  nor (_06273_, _06272_, _04734_);
  and (_06274_, _06273_, _06271_);
  and (_06275_, _05568_, _04734_);
  or (_06276_, _06275_, _04743_);
  or (_06277_, _06276_, _06274_);
  and (_06278_, _06277_, _06151_);
  or (_06279_, _06278_, _03758_);
  nand (_06280_, _05570_, _03758_);
  and (_06281_, _06280_, _03756_);
  and (_06282_, _06281_, _06279_);
  or (_06283_, _06282_, _06150_);
  and (_06284_, _06283_, _03428_);
  or (_06285_, _06258_, _03428_);
  nand (_06286_, _06285_, _03840_);
  or (_06287_, _06286_, _06284_);
  nand (_06288_, _05570_, _03841_);
  and (_06289_, _06288_, _06287_);
  or (_06290_, _06289_, _05131_);
  and (_06291_, _06248_, _05421_);
  nand (_06292_, _05522_, _05131_);
  or (_06293_, _06292_, _06291_);
  and (_06294_, _06293_, _05183_);
  and (_06295_, _06294_, _06290_);
  or (_06296_, _06295_, _06144_);
  and (_06297_, _06296_, _06141_);
  nand (_06298_, _06257_, _03456_);
  nand (_06299_, _06298_, _03735_);
  or (_06300_, _06299_, _06297_);
  or (_06301_, _05568_, _03735_);
  and (_06302_, _06301_, _06300_);
  or (_06303_, _06302_, _03739_);
  not (_06304_, _03740_);
  not (_06305_, _03739_);
  or (_06306_, _06248_, _06305_);
  and (_06307_, _06306_, _06304_);
  and (_06308_, _06307_, _06303_);
  not (_06309_, _06138_);
  nor (_06310_, _03647_, _03820_);
  not (_06311_, _06310_);
  and (_06312_, _03993_, _01924_);
  and (_06313_, _03974_, _01911_);
  nor (_06314_, _06313_, _06312_);
  and (_06315_, _03971_, _01980_);
  and (_06316_, _03987_, _01976_);
  nor (_06317_, _06316_, _06315_);
  and (_06318_, _06317_, _06314_);
  and (_06319_, _04000_, _01991_);
  and (_06320_, _03989_, _01988_);
  nor (_06321_, _06320_, _06319_);
  and (_06322_, _03969_, _01958_);
  and (_06323_, _03961_, _01967_);
  nor (_06324_, _06323_, _06322_);
  and (_06325_, _06324_, _06321_);
  and (_06326_, _06325_, _06318_);
  and (_06327_, _03982_, _01938_);
  and (_06328_, _03984_, _01954_);
  nor (_06329_, _06328_, _06327_);
  and (_06330_, _03952_, _42427_);
  and (_06331_, _03976_, _01929_);
  nor (_06332_, _06331_, _06330_);
  and (_06333_, _06332_, _06329_);
  and (_06334_, _03995_, _01971_);
  and (_06335_, _03965_, _01985_);
  nor (_06336_, _06335_, _06334_);
  and (_06337_, _03998_, _01933_);
  and (_06338_, _03957_, _01948_);
  nor (_06339_, _06338_, _06337_);
  and (_06340_, _06339_, _06336_);
  and (_06341_, _06340_, _06333_);
  and (_06342_, _06341_, _06326_);
  and (_06343_, _06342_, _05568_);
  and (_06344_, _04595_, _04382_);
  not (_06345_, _04005_);
  and (_06346_, _04180_, _06345_);
  and (_06347_, _06346_, _06344_);
  not (_06348_, _06342_);
  and (_06349_, _03952_, _42462_);
  and (_06350_, _03989_, _02417_);
  nor (_06351_, _06350_, _06349_);
  and (_06352_, _03998_, _02396_);
  and (_06353_, _03965_, _02424_);
  nor (_06354_, _06353_, _06352_);
  and (_06355_, _06354_, _06351_);
  and (_06356_, _03984_, _02402_);
  and (_06357_, _04000_, _02427_);
  nor (_06358_, _06357_, _06356_);
  and (_06359_, _03969_, _02430_);
  and (_06360_, _03971_, _02411_);
  nor (_06361_, _06360_, _06359_);
  and (_06362_, _06361_, _06358_);
  and (_06363_, _06362_, _06355_);
  and (_06364_, _03961_, _02407_);
  and (_06365_, _03987_, _02409_);
  nor (_06366_, _06365_, _06364_);
  and (_06367_, _03993_, _02394_);
  and (_06368_, _03982_, _02432_);
  nor (_06369_, _06368_, _06367_);
  and (_06370_, _06369_, _06366_);
  and (_06371_, _03976_, _02398_);
  and (_06372_, _03957_, _02434_);
  nor (_06373_, _06372_, _06371_);
  and (_06374_, _03974_, _02422_);
  and (_06375_, _03995_, _02415_);
  nor (_06376_, _06375_, _06374_);
  and (_06377_, _06376_, _06373_);
  and (_06378_, _06377_, _06370_);
  and (_06379_, _06378_, _06363_);
  and (_06380_, _06379_, _06348_);
  and (_06381_, _03952_, _42457_);
  and (_06382_, _03965_, _02379_);
  nor (_06383_, _06382_, _06381_);
  and (_06384_, _03998_, _02351_);
  and (_06385_, _03987_, _02364_);
  nor (_06386_, _06385_, _06384_);
  and (_06387_, _06386_, _06383_);
  and (_06388_, _03984_, _02357_);
  and (_06389_, _04000_, _02381_);
  nor (_06390_, _06389_, _06388_);
  and (_06391_, _03969_, _02384_);
  and (_06392_, _03971_, _02366_);
  nor (_06393_, _06392_, _06391_);
  and (_06394_, _06393_, _06390_);
  and (_06395_, _06394_, _06387_);
  and (_06396_, _03961_, _02362_);
  and (_06397_, _03989_, _02372_);
  nor (_06398_, _06397_, _06396_);
  and (_06399_, _03993_, _02349_);
  and (_06400_, _03982_, _02386_);
  nor (_06401_, _06400_, _06399_);
  and (_06402_, _06401_, _06398_);
  and (_06403_, _03976_, _02353_);
  and (_06404_, _03957_, _02388_);
  nor (_06405_, _06404_, _06403_);
  and (_06406_, _03974_, _02377_);
  and (_06407_, _03995_, _02370_);
  nor (_06408_, _06407_, _06406_);
  and (_06409_, _06408_, _06405_);
  and (_06410_, _06409_, _06402_);
  and (_06411_, _06410_, _06395_);
  and (_06412_, _03952_, _42452_);
  and (_06413_, _03957_, _02343_);
  nor (_06414_, _06413_, _06412_);
  and (_06415_, _03982_, _02341_);
  and (_06416_, _03987_, _02319_);
  nor (_06417_, _06416_, _06415_);
  and (_06418_, _06417_, _06414_);
  and (_06419_, _03993_, _02304_);
  and (_06420_, _03974_, _02332_);
  nor (_06421_, _06420_, _06419_);
  and (_06422_, _03969_, _02312_);
  and (_06423_, _03961_, _02317_);
  nor (_06424_, _06423_, _06422_);
  and (_06425_, _06424_, _06421_);
  and (_06426_, _06425_, _06418_);
  and (_06427_, _03971_, _02321_);
  and (_06428_, _04000_, _02336_);
  nor (_06429_, _06428_, _06427_);
  and (_06430_, _03965_, _02334_);
  and (_06431_, _03989_, _02327_);
  nor (_06432_, _06431_, _06430_);
  and (_06433_, _06432_, _06429_);
  and (_06434_, _03976_, _02308_);
  and (_06435_, _03995_, _02325_);
  nor (_06436_, _06435_, _06434_);
  and (_06437_, _03998_, _02306_);
  and (_06438_, _03984_, _02339_);
  nor (_06439_, _06438_, _06437_);
  and (_06440_, _06439_, _06436_);
  and (_06441_, _06440_, _06433_);
  and (_06442_, _06441_, _06426_);
  nor (_06443_, _06442_, _06411_);
  and (_06444_, _06443_, _06380_);
  and (_06445_, _06444_, _06347_);
  and (_06446_, _06445_, \oc8051_golden_model_1.IP [7]);
  not (_06447_, _06411_);
  and (_06448_, _06442_, _06447_);
  and (_06449_, _04180_, _04005_);
  and (_06450_, _06449_, _06344_);
  nor (_06451_, _06379_, _06342_);
  and (_06452_, _06451_, _06450_);
  and (_06453_, _06452_, _06448_);
  and (_06454_, _06453_, \oc8051_golden_model_1.ACC [7]);
  nor (_06455_, _06454_, _06446_);
  not (_06456_, _06442_);
  and (_06457_, _06456_, _06411_);
  and (_06458_, _06457_, _06452_);
  and (_06459_, _06458_, \oc8051_golden_model_1.PSW [7]);
  and (_06460_, _06452_, _06443_);
  and (_06461_, _06460_, \oc8051_golden_model_1.B [7]);
  nor (_06462_, _06461_, _06459_);
  and (_06463_, _06462_, _06455_);
  and (_06464_, _06442_, _06380_);
  and (_06465_, _06464_, _06411_);
  and (_06466_, _06465_, _06449_);
  not (_06467_, _04595_);
  and (_06468_, _06467_, _04382_);
  and (_06469_, _06468_, _06466_);
  and (_06470_, _06469_, \oc8051_golden_model_1.DPL [7]);
  and (_06471_, _06468_, _06346_);
  and (_06472_, _06471_, _06465_);
  and (_06473_, _06472_, \oc8051_golden_model_1.TL0 [7]);
  nor (_06474_, _06473_, _06470_);
  nor (_06475_, _04595_, _04382_);
  and (_06476_, _06475_, _06465_);
  and (_06477_, _06476_, _06449_);
  and (_06478_, _06477_, \oc8051_golden_model_1.DPH [7]);
  not (_06479_, _04382_);
  and (_06480_, _04595_, _06479_);
  nor (_06481_, _04180_, _04005_);
  and (_06482_, _06481_, _06465_);
  and (_06483_, _06482_, _06480_);
  and (_06484_, _06483_, \oc8051_golden_model_1.TH1 [7]);
  nor (_06485_, _06484_, _06478_);
  and (_06486_, _06485_, _06474_);
  and (_06487_, _06486_, _06463_);
  and (_06488_, _06482_, _06344_);
  and (_06489_, _06488_, \oc8051_golden_model_1.TH0 [7]);
  and (_06490_, _06476_, _06346_);
  and (_06491_, _06490_, \oc8051_golden_model_1.TL1 [7]);
  nor (_06492_, _06491_, _06489_);
  and (_06493_, _06465_, _06347_);
  and (_06494_, _06493_, \oc8051_golden_model_1.TCON [7]);
  not (_06495_, _04180_);
  and (_06496_, _06495_, _04005_);
  and (_06497_, _06496_, _06476_);
  and (_06498_, _06497_, \oc8051_golden_model_1.PCON [7]);
  nor (_06499_, _06498_, _06494_);
  and (_06500_, _06499_, _06492_);
  and (_06501_, _06465_, _06450_);
  and (_06502_, _06501_, \oc8051_golden_model_1.P0INREG [7]);
  not (_06503_, _06502_);
  and (_06504_, _06457_, _06380_);
  and (_06505_, _06504_, _06450_);
  and (_06506_, _06505_, \oc8051_golden_model_1.P1INREG [7]);
  and (_06507_, _06450_, _06444_);
  and (_06508_, _06507_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06509_, _06508_, _06506_);
  and (_06510_, _06509_, _06503_);
  and (_06511_, _06480_, _06346_);
  and (_06512_, _06511_, _06465_);
  and (_06513_, _06512_, \oc8051_golden_model_1.TMOD [7]);
  and (_06514_, _06448_, _06380_);
  and (_06515_, _06514_, _06450_);
  and (_06516_, _06515_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_06517_, _06516_, _06513_);
  and (_06518_, _06517_, _06510_);
  and (_06519_, _06480_, _06466_);
  and (_06520_, _06519_, \oc8051_golden_model_1.SP [7]);
  not (_06521_, _06520_);
  and (_06522_, _06514_, _06347_);
  and (_06523_, _06522_, \oc8051_golden_model_1.IE [7]);
  not (_06524_, _06523_);
  and (_06525_, _06504_, _06347_);
  and (_06526_, _06525_, \oc8051_golden_model_1.SCON [7]);
  and (_06527_, _06511_, _06504_);
  and (_06528_, _06527_, \oc8051_golden_model_1.SBUF [7]);
  nor (_06529_, _06528_, _06526_);
  and (_06530_, _06529_, _06524_);
  and (_06531_, _06530_, _06521_);
  and (_06532_, _06531_, _06518_);
  and (_06533_, _06532_, _06500_);
  and (_06534_, _06533_, _06487_);
  not (_06535_, _06534_);
  nor (_06536_, _06535_, _06343_);
  nor (_06537_, _06536_, _06311_);
  or (_06538_, _06537_, _06309_);
  or (_06539_, _06538_, _06308_);
  and (_06540_, _06539_, _06140_);
  and (_06541_, _06348_, _04779_);
  or (_06542_, _06541_, _03401_);
  or (_06543_, _06542_, _06540_);
  and (_06544_, _06258_, _03401_);
  nor (_06545_, _06544_, _04791_);
  and (_06546_, _06545_, _06543_);
  and (_06547_, _06342_, _05570_);
  nor (_06548_, _06342_, _05570_);
  nor (_06549_, _06548_, _06547_);
  and (_06550_, _06549_, _04791_);
  or (_06551_, _06550_, _04793_);
  or (_06552_, _06551_, _06546_);
  not (_06553_, _04793_);
  not (_06554_, \oc8051_golden_model_1.ACC [7]);
  nor (_06555_, _05570_, _06554_);
  and (_06556_, _05570_, _06554_);
  nor (_06557_, _06556_, _06555_);
  or (_06558_, _06557_, _06553_);
  and (_06559_, _06558_, _04789_);
  and (_06560_, _06559_, _06552_);
  and (_06561_, _06548_, _04788_);
  or (_06562_, _06561_, _06560_);
  and (_06563_, _06562_, _04787_);
  and (_06564_, _06555_, _04786_);
  or (_06565_, _06564_, _03388_);
  or (_06566_, _06565_, _06563_);
  not (_06567_, _03914_);
  nor (_06568_, _06567_, _03647_);
  and (_06569_, _06258_, _03388_);
  nor (_06570_, _06569_, _06568_);
  and (_06571_, _06570_, _06566_);
  not (_06572_, _04011_);
  nor (_06573_, _06572_, _03647_);
  not (_06574_, _06568_);
  nor (_06575_, _06547_, _06574_);
  or (_06576_, _06575_, _06573_);
  or (_06577_, _06576_, _06571_);
  nand (_06578_, _06556_, _06573_);
  and (_06579_, _06578_, _03384_);
  and (_06580_, _06579_, _06577_);
  nand (_06581_, _06257_, _03383_);
  and (_06582_, _03730_, _03244_);
  or (_06583_, _04632_, _06582_);
  and (_06584_, _03767_, _03244_);
  nor (_06585_, _06584_, _04200_);
  not (_06586_, _06585_);
  nor (_06587_, _06586_, _06583_);
  nand (_06588_, _06587_, _06581_);
  or (_06589_, _06588_, _06580_);
  not (_06590_, _05053_);
  or (_06591_, _06587_, _06132_);
  and (_06592_, _06591_, _06590_);
  and (_06593_, _06592_, _06589_);
  or (_06594_, _06593_, _06134_);
  not (_06595_, _04811_);
  not (_06596_, _06248_);
  or (_06597_, _06200_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_06598_, _06202_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_06599_, _06598_, _06193_);
  and (_06600_, _06599_, _06597_);
  or (_06601_, _06202_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_06602_, _06200_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_06603_, _06602_, _06206_);
  and (_06604_, _06603_, _06601_);
  nor (_06605_, _06604_, _06600_);
  nand (_06606_, _06605_, _06185_);
  or (_06607_, _06200_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_06608_, _06202_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_06609_, _06608_, _06193_);
  and (_06610_, _06609_, _06607_);
  or (_06611_, _06202_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_06612_, _06200_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_06613_, _06612_, _06206_);
  and (_06614_, _06613_, _06611_);
  nor (_06615_, _06614_, _06610_);
  nand (_06616_, _06615_, _06186_);
  nand (_06617_, _06616_, _06606_);
  nand (_06618_, _06617_, _06225_);
  nand (_06619_, _06202_, \oc8051_golden_model_1.IRAM[1] [6]);
  nand (_06620_, _06200_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_06621_, _06620_, _06193_);
  nand (_06622_, _06621_, _06619_);
  nand (_06623_, _06200_, \oc8051_golden_model_1.IRAM[2] [6]);
  nand (_06624_, _06202_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_06625_, _06624_, _06206_);
  nand (_06626_, _06625_, _06623_);
  nand (_06627_, _06626_, _06622_);
  nand (_06628_, _06627_, _06185_);
  nand (_06629_, _06200_, \oc8051_golden_model_1.IRAM[4] [6]);
  nand (_06630_, _06202_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_06631_, _06630_, _06193_);
  nand (_06632_, _06631_, _06629_);
  nand (_06633_, _06200_, \oc8051_golden_model_1.IRAM[6] [6]);
  nand (_06634_, _06202_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_06635_, _06634_, _06206_);
  nand (_06636_, _06635_, _06633_);
  nand (_06637_, _06636_, _06632_);
  nand (_06638_, _06637_, _06186_);
  nand (_06639_, _06638_, _06628_);
  nand (_06640_, _06639_, _06176_);
  and (_06641_, _06640_, _06618_);
  not (_06642_, _06641_);
  or (_06643_, _06200_, \oc8051_golden_model_1.IRAM[9] [1]);
  or (_06644_, _06202_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_06645_, _06644_, _06193_);
  and (_06646_, _06645_, _06643_);
  or (_06648_, _06202_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_06649_, _06200_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_06650_, _06649_, _06206_);
  and (_06651_, _06650_, _06648_);
  nor (_06652_, _06651_, _06646_);
  nand (_06653_, _06652_, _06185_);
  or (_06654_, _06200_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_06655_, _06202_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_06656_, _06655_, _06193_);
  and (_06657_, _06656_, _06654_);
  or (_06658_, _06202_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_06659_, _06200_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_06660_, _06659_, _06206_);
  and (_06661_, _06660_, _06658_);
  nor (_06662_, _06661_, _06657_);
  nand (_06663_, _06662_, _06186_);
  nand (_06664_, _06663_, _06653_);
  nand (_06665_, _06664_, _06225_);
  or (_06666_, _06200_, _04850_);
  or (_06667_, _06202_, _04848_);
  and (_06668_, _06667_, _06193_);
  nand (_06669_, _06668_, _06666_);
  or (_06670_, _06202_, _04856_);
  or (_06671_, _06200_, _04854_);
  and (_06672_, _06671_, _06206_);
  nand (_06673_, _06672_, _06670_);
  nand (_06674_, _06673_, _06669_);
  nand (_06675_, _06674_, _06185_);
  or (_06676_, _06202_, _04868_);
  or (_06677_, _06200_, _04870_);
  and (_06678_, _06677_, _06193_);
  nand (_06679_, _06678_, _06676_);
  or (_06680_, _06202_, _04864_);
  or (_06681_, _06200_, _04862_);
  and (_06682_, _06681_, _06206_);
  nand (_06683_, _06682_, _06680_);
  nand (_06684_, _06683_, _06679_);
  nand (_06685_, _06684_, _06186_);
  nand (_06686_, _06685_, _06675_);
  nand (_06687_, _06686_, _06176_);
  nand (_06688_, _06687_, _06665_);
  or (_06689_, _06200_, \oc8051_golden_model_1.IRAM[9] [0]);
  or (_06690_, _06202_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_06691_, _06690_, _06193_);
  and (_06692_, _06691_, _06689_);
  or (_06693_, _06202_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_06694_, _06200_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_06695_, _06694_, _06206_);
  and (_06696_, _06695_, _06693_);
  nor (_06697_, _06696_, _06692_);
  nand (_06698_, _06697_, _06185_);
  or (_06699_, _06200_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_06700_, _06202_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_06701_, _06700_, _06193_);
  and (_06702_, _06701_, _06699_);
  or (_06703_, _06202_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_06704_, _06200_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_06705_, _06704_, _06206_);
  and (_06706_, _06705_, _06703_);
  nor (_06707_, _06706_, _06702_);
  nand (_06708_, _06707_, _06186_);
  nand (_06709_, _06708_, _06698_);
  nand (_06710_, _06709_, _06225_);
  or (_06711_, _06200_, _04645_);
  or (_06712_, _06202_, _04245_);
  and (_06713_, _06712_, _06193_);
  nand (_06714_, _06713_, _06711_);
  or (_06715_, _06202_, _04653_);
  or (_06716_, _06200_, _04650_);
  and (_06717_, _06716_, _06206_);
  nand (_06718_, _06717_, _06715_);
  nand (_06719_, _06718_, _06714_);
  nand (_06720_, _06719_, _06185_);
  or (_06721_, _06202_, _04666_);
  or (_06722_, _06200_, _04668_);
  and (_06723_, _06722_, _06193_);
  nand (_06724_, _06723_, _06721_);
  or (_06725_, _06202_, _04662_);
  or (_06726_, _06200_, _04660_);
  and (_06727_, _06726_, _06206_);
  nand (_06728_, _06727_, _06725_);
  nand (_06729_, _06728_, _06724_);
  nand (_06730_, _06729_, _06186_);
  nand (_06731_, _06730_, _06720_);
  nand (_06732_, _06731_, _06176_);
  nand (_06733_, _06732_, _06710_);
  and (_06734_, _06733_, _06688_);
  or (_06735_, _06200_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_06736_, _06202_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_06737_, _06736_, _06193_);
  and (_06738_, _06737_, _06735_);
  or (_06739_, _06202_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_06740_, _06200_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_06741_, _06740_, _06206_);
  and (_06742_, _06741_, _06739_);
  nor (_06743_, _06742_, _06738_);
  nand (_06744_, _06743_, _06185_);
  or (_06745_, _06200_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_06746_, _06202_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_06747_, _06746_, _06193_);
  and (_06748_, _06747_, _06745_);
  or (_06749_, _06202_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_06750_, _06200_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_06751_, _06750_, _06206_);
  and (_06752_, _06751_, _06749_);
  nor (_06753_, _06752_, _06748_);
  nand (_06754_, _06753_, _06186_);
  nand (_06755_, _06754_, _06744_);
  nand (_06756_, _06755_, _06225_);
  nand (_06757_, _06202_, \oc8051_golden_model_1.IRAM[1] [3]);
  nand (_06758_, _06200_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_06759_, _06758_, _06193_);
  nand (_06760_, _06759_, _06757_);
  nand (_06761_, _06200_, \oc8051_golden_model_1.IRAM[2] [3]);
  nand (_06762_, _06202_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_06763_, _06762_, _06206_);
  nand (_06764_, _06763_, _06761_);
  nand (_06765_, _06764_, _06760_);
  nand (_06766_, _06765_, _06185_);
  nand (_06767_, _06200_, \oc8051_golden_model_1.IRAM[4] [3]);
  nand (_06768_, _06202_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_06769_, _06768_, _06193_);
  nand (_06770_, _06769_, _06767_);
  nand (_06771_, _06200_, \oc8051_golden_model_1.IRAM[6] [3]);
  nand (_06772_, _06202_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_06773_, _06772_, _06206_);
  nand (_06774_, _06773_, _06771_);
  nand (_06775_, _06774_, _06770_);
  nand (_06776_, _06775_, _06186_);
  nand (_06777_, _06776_, _06766_);
  nand (_06778_, _06777_, _06176_);
  nand (_06779_, _06778_, _06756_);
  or (_06780_, _06200_, \oc8051_golden_model_1.IRAM[9] [2]);
  or (_06781_, _06202_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_06782_, _06781_, _06193_);
  and (_06783_, _06782_, _06780_);
  or (_06784_, _06202_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_06785_, _06200_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_06786_, _06785_, _06206_);
  and (_06787_, _06786_, _06784_);
  nor (_06788_, _06787_, _06783_);
  nand (_06789_, _06788_, _06185_);
  or (_06790_, _06200_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_06791_, _06202_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_06792_, _06791_, _06193_);
  and (_06793_, _06792_, _06790_);
  or (_06794_, _06202_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_06795_, _06200_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_06796_, _06795_, _06206_);
  and (_06797_, _06796_, _06794_);
  nor (_06798_, _06797_, _06793_);
  nand (_06799_, _06798_, _06186_);
  nand (_06800_, _06799_, _06789_);
  nand (_06801_, _06800_, _06225_);
  or (_06802_, _06200_, _05257_);
  or (_06803_, _06202_, _05255_);
  and (_06804_, _06803_, _06193_);
  nand (_06805_, _06804_, _06802_);
  or (_06806_, _06202_, _05263_);
  or (_06807_, _06200_, _05261_);
  and (_06808_, _06807_, _06206_);
  nand (_06809_, _06808_, _06806_);
  nand (_06810_, _06809_, _06805_);
  nand (_06811_, _06810_, _06185_);
  or (_06812_, _06202_, _05275_);
  or (_06813_, _06200_, _05277_);
  and (_06814_, _06813_, _06193_);
  nand (_06815_, _06814_, _06812_);
  or (_06816_, _06202_, _05271_);
  or (_06817_, _06200_, _05269_);
  and (_06818_, _06817_, _06206_);
  nand (_06819_, _06818_, _06816_);
  nand (_06820_, _06819_, _06815_);
  nand (_06821_, _06820_, _06186_);
  nand (_06822_, _06821_, _06811_);
  nand (_06823_, _06822_, _06176_);
  nand (_06824_, _06823_, _06801_);
  and (_06825_, _06824_, _06779_);
  and (_06826_, _06825_, _06734_);
  or (_06827_, _06200_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_06828_, _06202_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_06829_, _06828_, _06193_);
  and (_06830_, _06829_, _06827_);
  or (_06831_, _06202_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_06832_, _06200_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_06833_, _06832_, _06206_);
  and (_06834_, _06833_, _06831_);
  nor (_06835_, _06834_, _06830_);
  nand (_06836_, _06835_, _06185_);
  or (_06837_, _06200_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_06838_, _06202_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_06839_, _06838_, _06193_);
  and (_06840_, _06839_, _06837_);
  or (_06841_, _06202_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_06842_, _06200_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_06843_, _06842_, _06206_);
  and (_06844_, _06843_, _06841_);
  nor (_06845_, _06844_, _06840_);
  nand (_06846_, _06845_, _06186_);
  nand (_06847_, _06846_, _06836_);
  nand (_06848_, _06847_, _06225_);
  nand (_06849_, _06202_, \oc8051_golden_model_1.IRAM[1] [5]);
  nand (_06850_, _06200_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_06851_, _06850_, _06193_);
  nand (_06852_, _06851_, _06849_);
  nand (_06853_, _06200_, \oc8051_golden_model_1.IRAM[2] [5]);
  nand (_06854_, _06202_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_06855_, _06854_, _06206_);
  nand (_06856_, _06855_, _06853_);
  nand (_06857_, _06856_, _06852_);
  nand (_06858_, _06857_, _06185_);
  not (_06859_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_06860_, _06202_, _06859_);
  not (_06861_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_06862_, _06200_, _06861_);
  and (_06863_, _06862_, _06193_);
  nand (_06864_, _06863_, _06860_);
  nand (_06865_, _06200_, \oc8051_golden_model_1.IRAM[6] [5]);
  nand (_06866_, _06202_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_06867_, _06866_, _06206_);
  nand (_06868_, _06867_, _06865_);
  nand (_06869_, _06868_, _06864_);
  nand (_06870_, _06869_, _06186_);
  nand (_06871_, _06870_, _06858_);
  nand (_06872_, _06871_, _06176_);
  nand (_06873_, _06872_, _06848_);
  or (_06874_, _06200_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_06875_, _06202_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_06876_, _06875_, _06193_);
  and (_06877_, _06876_, _06874_);
  or (_06878_, _06202_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_06879_, _06200_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_06880_, _06879_, _06206_);
  and (_06881_, _06880_, _06878_);
  nor (_06882_, _06881_, _06877_);
  nand (_06883_, _06882_, _06185_);
  or (_06884_, _06200_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_06885_, _06202_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_06886_, _06885_, _06193_);
  and (_06887_, _06886_, _06884_);
  or (_06888_, _06202_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_06889_, _06200_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_06890_, _06889_, _06206_);
  and (_06891_, _06890_, _06888_);
  nor (_06892_, _06891_, _06887_);
  nand (_06893_, _06892_, _06186_);
  nand (_06894_, _06893_, _06883_);
  nand (_06895_, _06894_, _06225_);
  nand (_06896_, _06202_, \oc8051_golden_model_1.IRAM[1] [4]);
  nand (_06897_, _06200_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_06898_, _06897_, _06193_);
  nand (_06899_, _06898_, _06896_);
  nand (_06900_, _06200_, \oc8051_golden_model_1.IRAM[2] [4]);
  nand (_06901_, _06202_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_06902_, _06901_, _06206_);
  nand (_06903_, _06902_, _06900_);
  nand (_06904_, _06903_, _06899_);
  nand (_06905_, _06904_, _06185_);
  nand (_06906_, _06200_, \oc8051_golden_model_1.IRAM[4] [4]);
  nand (_06907_, _06202_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_06908_, _06907_, _06193_);
  nand (_06909_, _06908_, _06906_);
  nand (_06910_, _06200_, \oc8051_golden_model_1.IRAM[6] [4]);
  nand (_06911_, _06202_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_06912_, _06911_, _06206_);
  nand (_06913_, _06912_, _06910_);
  nand (_06914_, _06913_, _06909_);
  nand (_06915_, _06914_, _06186_);
  nand (_06916_, _06915_, _06905_);
  nand (_06917_, _06916_, _06176_);
  nand (_06918_, _06917_, _06895_);
  and (_06919_, _06918_, _06873_);
  and (_06920_, _06919_, _06826_);
  and (_06921_, _06920_, _06642_);
  nor (_06922_, _06921_, _06596_);
  and (_06923_, _06921_, _06596_);
  or (_06924_, _06923_, _06922_);
  or (_06925_, _06924_, _04813_);
  and (_06926_, _06925_, _06595_);
  and (_06927_, _06926_, _06594_);
  and (_06928_, _06160_, _04811_);
  or (_06929_, _06928_, _03899_);
  or (_06930_, _06929_, _06927_);
  and (_06931_, _03123_, _03102_);
  and (_06932_, _06931_, _06253_);
  and (_06933_, _06932_, \oc8051_golden_model_1.PC [7]);
  nor (_06934_, _06932_, \oc8051_golden_model_1.PC [7]);
  nor (_06935_, _06934_, _06933_);
  not (_06936_, _06935_);
  nand (_06937_, _06936_, _03899_);
  and (_06938_, _06937_, _06930_);
  or (_06939_, _06938_, _03414_);
  and (_06940_, _06258_, _03414_);
  nor (_06941_, _06940_, _03681_);
  and (_06942_, _06941_, _06939_);
  or (_06943_, _06942_, _06122_);
  and (_06944_, _06943_, _04482_);
  and (_06945_, _04900_, _04700_);
  and (_06946_, _05307_, _05119_);
  and (_06947_, _06946_, _06945_);
  and (_06948_, _05950_, _05857_);
  and (_06949_, _06948_, _06947_);
  or (_06950_, _06949_, _05568_);
  nor (_06951_, _06065_, _05568_);
  and (_06952_, _06065_, _05568_);
  nor (_06953_, _06952_, _06951_);
  not (_06954_, _06953_);
  nand (_06955_, _06954_, _06949_);
  and (_06956_, _06955_, _04483_);
  and (_06957_, _06956_, _06950_);
  or (_06958_, _06957_, _04826_);
  or (_06959_, _06958_, _06944_);
  not (_06960_, _04831_);
  and (_06961_, _06687_, _06665_);
  and (_06962_, _06732_, _06710_);
  and (_06963_, _06962_, _06961_);
  and (_06964_, _06778_, _06756_);
  and (_06965_, _06823_, _06801_);
  and (_06966_, _06965_, _06964_);
  and (_06967_, _06966_, _06963_);
  and (_06968_, _06872_, _06848_);
  and (_06969_, _06917_, _06895_);
  and (_06970_, _06969_, _06968_);
  and (_06971_, _06970_, _06967_);
  and (_06972_, _06971_, _06641_);
  nor (_06973_, _06972_, _06596_);
  and (_06974_, _06972_, _06596_);
  or (_06975_, _06974_, _06973_);
  or (_06976_, _06975_, _04827_);
  and (_06977_, _06976_, _06960_);
  and (_06978_, _06977_, _06959_);
  or (_06979_, _06978_, _06078_);
  and (_06980_, _06979_, _05407_);
  or (_06981_, _06980_, _05415_);
  and (_06982_, _06981_, _05405_);
  not (_06983_, \oc8051_golden_model_1.PC [15]);
  and (_06984_, _06933_, \oc8051_golden_model_1.PC [8]);
  and (_06985_, _06984_, \oc8051_golden_model_1.PC [9]);
  and (_06986_, _06985_, \oc8051_golden_model_1.PC [10]);
  and (_06987_, _06986_, \oc8051_golden_model_1.PC [11]);
  and (_06988_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and (_06989_, _06988_, _06987_);
  and (_06990_, _06989_, \oc8051_golden_model_1.PC [14]);
  and (_06991_, _06990_, _06983_);
  nor (_06992_, _06990_, _06983_);
  or (_06993_, _06992_, _06991_);
  or (_06994_, _06993_, _03900_);
  and (_06995_, _06255_, \oc8051_golden_model_1.PC [8]);
  and (_06996_, _06995_, \oc8051_golden_model_1.PC [9]);
  and (_06997_, _06996_, \oc8051_golden_model_1.PC [10]);
  and (_06998_, _06997_, \oc8051_golden_model_1.PC [11]);
  and (_06999_, _06998_, _06988_);
  and (_07000_, _06999_, \oc8051_golden_model_1.PC [14]);
  and (_07001_, _07000_, _06983_);
  nor (_07002_, _07000_, _06983_);
  or (_07003_, _07002_, _07001_);
  or (_07004_, _07003_, _03899_);
  and (_07005_, _07004_, _06994_);
  and (_07006_, _07005_, _05400_);
  and (_07007_, _07006_, _05403_);
  or (_40679_, _07007_, _06982_);
  not (_07008_, \oc8051_golden_model_1.B [7]);
  nor (_07009_, _43152_, _07008_);
  and (_07010_, _03919_, _03397_);
  not (_07011_, _07010_);
  and (_07012_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_07013_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_07014_, _07013_, _07012_);
  not (_07015_, \oc8051_golden_model_1.B [1]);
  nor (_07016_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_07017_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_07018_, _07017_, _07016_);
  and (_07019_, _07018_, _07015_);
  nor (_07020_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not (_07021_, _07020_);
  and (_07022_, \oc8051_golden_model_1.B [0], _06554_);
  nor (_07023_, _07022_, _07021_);
  and (_07024_, _07023_, _07019_);
  and (_07025_, _07024_, _07014_);
  or (_07026_, _07024_, _06554_);
  not (_07027_, \oc8051_golden_model_1.B [2]);
  not (_07028_, \oc8051_golden_model_1.B [3]);
  not (_07029_, \oc8051_golden_model_1.B [4]);
  not (_07030_, \oc8051_golden_model_1.B [5]);
  nor (_07031_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_07032_, _07031_, _07030_);
  and (_07033_, _07032_, _07029_);
  and (_07034_, _07033_, _07028_);
  and (_07035_, _07034_, _07027_);
  not (_07036_, \oc8051_golden_model_1.ACC [6]);
  and (_07037_, \oc8051_golden_model_1.B [0], _07036_);
  nor (_07038_, _07037_, _06554_);
  nor (_07039_, _07038_, _07015_);
  not (_07040_, _07039_);
  and (_07041_, _07040_, _07035_);
  nor (_07042_, _07041_, _07026_);
  nor (_07043_, _07042_, _07025_);
  and (_07044_, _07041_, \oc8051_golden_model_1.B [0]);
  nor (_07045_, _07044_, _07036_);
  and (_07046_, _07045_, _07015_);
  nor (_07047_, _07045_, _07015_);
  nor (_07048_, _07047_, _07046_);
  and (_07049_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_07050_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_07051_, _07050_, _07049_);
  nor (_07052_, _07051_, \oc8051_golden_model_1.ACC [4]);
  nor (_07053_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  not (_07054_, \oc8051_golden_model_1.B [0]);
  and (_07055_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_07056_, _07055_, _07054_);
  nor (_07057_, _07056_, _07053_);
  nor (_07058_, _07057_, _07052_);
  not (_07059_, _07058_);
  and (_07060_, _07059_, _07048_);
  nor (_07061_, _07043_, \oc8051_golden_model_1.B [2]);
  nor (_07062_, _07061_, _07046_);
  not (_07063_, _07062_);
  nor (_07064_, _07063_, _07060_);
  and (_07065_, \oc8051_golden_model_1.B [2], _06554_);
  nor (_07066_, _07065_, \oc8051_golden_model_1.B [7]);
  and (_07067_, _07066_, _07018_);
  not (_07068_, _07067_);
  nor (_07069_, _07068_, _07064_);
  nor (_07070_, _07069_, _07043_);
  nor (_07071_, _07070_, _07025_);
  and (_07072_, _07033_, \oc8051_golden_model_1.ACC [7]);
  nor (_07073_, _07072_, _07034_);
  nor (_07074_, _07059_, _07048_);
  nor (_07075_, _07074_, _07060_);
  not (_07076_, _07075_);
  and (_07077_, _07076_, _07069_);
  nor (_07078_, _07069_, _07045_);
  nor (_07079_, _07078_, _07077_);
  and (_07080_, _07079_, _07027_);
  nor (_07081_, _07079_, _07027_);
  nor (_07082_, _07081_, _07080_);
  not (_07083_, _07082_);
  not (_07084_, \oc8051_golden_model_1.ACC [5]);
  nor (_07085_, _07069_, _07084_);
  and (_07086_, _07069_, _07051_);
  or (_07087_, _07086_, _07085_);
  and (_07088_, _07087_, _07015_);
  nor (_07089_, _07087_, _07015_);
  not (_07090_, \oc8051_golden_model_1.ACC [4]);
  and (_07091_, \oc8051_golden_model_1.B [0], _07090_);
  nor (_07092_, _07091_, _07089_);
  nor (_07093_, _07092_, _07088_);
  nor (_07094_, _07093_, _07083_);
  nor (_07095_, _07071_, \oc8051_golden_model_1.B [3]);
  nor (_07096_, _07095_, _07080_);
  not (_07097_, _07096_);
  nor (_07098_, _07097_, _07094_);
  nor (_07099_, _07098_, _07073_);
  nor (_07100_, _07099_, _07071_);
  nor (_07101_, _07100_, _07025_);
  nor (_07102_, _07101_, \oc8051_golden_model_1.B [4]);
  not (_07103_, _07099_);
  and (_07104_, _07093_, _07083_);
  nor (_07105_, _07104_, _07094_);
  nor (_07106_, _07105_, _07103_);
  nor (_07107_, _07099_, _07079_);
  nor (_07108_, _07107_, _07106_);
  and (_07109_, _07108_, _07028_);
  nor (_07110_, _07108_, _07028_);
  nor (_07111_, _07110_, _07109_);
  not (_07112_, _07111_);
  nor (_07113_, _07099_, _07087_);
  nor (_07114_, _07089_, _07088_);
  and (_07115_, _07114_, _07091_);
  nor (_07116_, _07114_, _07091_);
  nor (_07117_, _07116_, _07115_);
  and (_07118_, _07117_, _07099_);
  or (_07119_, _07118_, _07113_);
  nor (_07120_, _07119_, \oc8051_golden_model_1.B [2]);
  and (_07121_, _07119_, \oc8051_golden_model_1.B [2]);
  nor (_07122_, _07099_, _07090_);
  and (_07123_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_07124_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_07125_, _07124_, _07123_);
  and (_07126_, _07099_, _07125_);
  or (_07127_, _07126_, _07122_);
  and (_07128_, _07127_, _07015_);
  and (_07129_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_07130_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_07131_, _07130_, _07129_);
  nor (_07132_, _07131_, \oc8051_golden_model_1.ACC [2]);
  nor (_07133_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_07134_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_07135_, _07134_, _07054_);
  nor (_07136_, _07135_, _07133_);
  nor (_07137_, _07136_, _07132_);
  not (_07138_, _07137_);
  nor (_07139_, _07127_, _07015_);
  nor (_07140_, _07139_, _07128_);
  and (_07141_, _07140_, _07138_);
  nor (_07142_, _07141_, _07128_);
  nor (_07143_, _07142_, _07121_);
  nor (_07144_, _07143_, _07120_);
  nor (_07145_, _07144_, _07112_);
  or (_07146_, _07145_, _07109_);
  nor (_07147_, _07146_, _07102_);
  and (_07148_, _07032_, \oc8051_golden_model_1.ACC [7]);
  or (_07149_, _07148_, _07033_);
  not (_07150_, _07149_);
  nor (_07151_, _07150_, _07147_);
  nor (_07152_, _07151_, _07101_);
  nor (_07153_, _07152_, _07025_);
  and (_07154_, _07031_, \oc8051_golden_model_1.ACC [7]);
  nor (_07155_, _07154_, _07032_);
  nor (_07156_, _07153_, \oc8051_golden_model_1.B [5]);
  and (_07157_, _07144_, _07112_);
  nor (_07158_, _07157_, _07145_);
  not (_07159_, _07158_);
  and (_07160_, _07159_, _07151_);
  nor (_07161_, _07151_, _07108_);
  nor (_07162_, _07161_, _07160_);
  and (_07163_, _07162_, _07029_);
  nor (_07164_, _07162_, _07029_);
  nor (_07165_, _07164_, _07163_);
  not (_07166_, _07165_);
  nor (_07167_, _07151_, _07119_);
  nor (_07168_, _07121_, _07120_);
  and (_07169_, _07168_, _07142_);
  nor (_07170_, _07168_, _07142_);
  nor (_07171_, _07170_, _07169_);
  not (_07172_, _07171_);
  and (_07173_, _07172_, _07151_);
  nor (_07174_, _07173_, _07167_);
  nor (_07175_, _07174_, \oc8051_golden_model_1.B [3]);
  and (_07176_, _07174_, \oc8051_golden_model_1.B [3]);
  nor (_07177_, _07140_, _07138_);
  nor (_07178_, _07177_, _07141_);
  not (_07179_, _07178_);
  and (_07180_, _07179_, _07151_);
  nor (_07181_, _07151_, _07127_);
  nor (_07182_, _07181_, _07180_);
  and (_07183_, _07182_, _07027_);
  not (_07184_, \oc8051_golden_model_1.ACC [3]);
  nor (_07185_, _07151_, _07184_);
  and (_07186_, _07151_, _07131_);
  or (_07187_, _07186_, _07185_);
  and (_07188_, _07187_, _07015_);
  nor (_07189_, _07187_, _07015_);
  not (_07190_, \oc8051_golden_model_1.ACC [2]);
  and (_07191_, \oc8051_golden_model_1.B [0], _07190_);
  nor (_07192_, _07191_, _07189_);
  nor (_07193_, _07192_, _07188_);
  nor (_07194_, _07182_, _07027_);
  nor (_07195_, _07194_, _07183_);
  not (_07196_, _07195_);
  nor (_07197_, _07196_, _07193_);
  nor (_07198_, _07197_, _07183_);
  nor (_07199_, _07198_, _07176_);
  nor (_07200_, _07199_, _07175_);
  nor (_07201_, _07200_, _07166_);
  or (_07202_, _07201_, _07163_);
  nor (_07203_, _07202_, _07156_);
  nor (_07204_, _07203_, _07155_);
  nor (_07205_, _07204_, _07153_);
  nor (_07206_, _07205_, _07025_);
  not (_07207_, _07204_);
  and (_07208_, _07200_, _07166_);
  nor (_07209_, _07208_, _07201_);
  nor (_07210_, _07209_, _07207_);
  nor (_07211_, _07204_, _07162_);
  nor (_07212_, _07211_, _07210_);
  and (_07213_, _07212_, _07030_);
  nor (_07214_, _07212_, _07030_);
  nor (_07215_, _07214_, _07213_);
  not (_07216_, _07215_);
  nor (_07217_, _07176_, _07175_);
  nor (_07218_, _07217_, _07198_);
  and (_07219_, _07217_, _07198_);
  or (_07220_, _07219_, _07218_);
  nor (_07221_, _07220_, _07207_);
  and (_07222_, _07207_, _07174_);
  nor (_07223_, _07222_, _07221_);
  and (_07224_, _07223_, _07029_);
  nor (_07225_, _07223_, _07029_);
  and (_07226_, _07196_, _07193_);
  nor (_07227_, _07226_, _07197_);
  nor (_07228_, _07227_, _07207_);
  nor (_07229_, _07204_, _07182_);
  nor (_07230_, _07229_, _07228_);
  and (_07231_, _07230_, _07028_);
  nor (_07232_, _07189_, _07188_);
  nor (_07233_, _07232_, _07191_);
  and (_07234_, _07232_, _07191_);
  or (_07235_, _07234_, _07233_);
  nor (_07236_, _07235_, _07207_);
  nor (_07237_, _07204_, _07187_);
  nor (_07238_, _07237_, _07236_);
  and (_07239_, _07238_, _07027_);
  nor (_07240_, _07238_, _07027_);
  nor (_07241_, _07204_, \oc8051_golden_model_1.ACC [2]);
  and (_07242_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07243_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07244_, _07243_, _07242_);
  nor (_07245_, _07207_, _07244_);
  nor (_07246_, _07245_, _07241_);
  and (_07247_, _07246_, _07015_);
  and (_07248_, \oc8051_golden_model_1.B [0], _03474_);
  not (_07249_, _07248_);
  nor (_07250_, _07246_, _07015_);
  nor (_07251_, _07250_, _07247_);
  and (_07252_, _07251_, _07249_);
  nor (_07253_, _07252_, _07247_);
  nor (_07254_, _07253_, _07240_);
  nor (_07255_, _07254_, _07239_);
  not (_07256_, _07255_);
  nor (_07257_, _07230_, _07028_);
  nor (_07258_, _07257_, _07231_);
  and (_07259_, _07258_, _07256_);
  nor (_07260_, _07259_, _07231_);
  nor (_07261_, _07260_, _07225_);
  nor (_07262_, _07261_, _07224_);
  nor (_07263_, _07262_, _07216_);
  nor (_07264_, _07206_, \oc8051_golden_model_1.B [6]);
  or (_07265_, _07264_, _07213_);
  or (_07266_, _07265_, _07263_);
  and (_07267_, \oc8051_golden_model_1.B [6], _06554_);
  nor (_07268_, _07267_, \oc8051_golden_model_1.B [7]);
  and (_07269_, _07268_, _07266_);
  nor (_07270_, _07269_, _07206_);
  or (_07271_, _07270_, _07025_);
  and (_07272_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  nor (_07273_, _07271_, \oc8051_golden_model_1.B [7]);
  nor (_07274_, _07273_, _07272_);
  not (_07275_, \oc8051_golden_model_1.B [6]);
  and (_07276_, _07262_, _07216_);
  nor (_07277_, _07276_, _07263_);
  not (_07278_, _07277_);
  and (_07279_, _07278_, _07269_);
  nor (_07280_, _07269_, _07212_);
  nor (_07281_, _07280_, _07279_);
  nor (_07282_, _07281_, _07275_);
  not (_07283_, _07282_);
  nor (_07284_, _07283_, _07274_);
  nor (_07285_, _07240_, _07239_);
  nor (_07286_, _07285_, _07253_);
  and (_07287_, _07285_, _07253_);
  nor (_07288_, _07287_, _07286_);
  and (_07289_, _07288_, _07269_);
  nor (_07290_, _07269_, _07238_);
  or (_07291_, _07290_, _07289_);
  nor (_07292_, _07291_, \oc8051_golden_model_1.B [3]);
  and (_07293_, _07291_, \oc8051_golden_model_1.B [3]);
  nor (_07294_, _07293_, _07292_);
  nor (_07295_, _07251_, _07249_);
  nor (_07296_, _07295_, _07252_);
  and (_07297_, _07296_, _07269_);
  not (_07298_, _07246_);
  nor (_07299_, _07269_, _07298_);
  nor (_07300_, _07299_, _07297_);
  and (_07301_, _07300_, \oc8051_golden_model_1.B [2]);
  nor (_07302_, _07300_, \oc8051_golden_model_1.B [2]);
  nor (_07303_, _07302_, _07301_);
  and (_07304_, _07303_, _07294_);
  nor (_07305_, _07269_, \oc8051_golden_model_1.ACC [1]);
  and (_07306_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07307_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  or (_07308_, _07307_, _07306_);
  and (_07309_, _07269_, _07308_);
  nor (_07310_, _07309_, _07305_);
  and (_07311_, _07310_, _07015_);
  nor (_07312_, _07310_, _07015_);
  and (_07313_, _07054_, \oc8051_golden_model_1.ACC [0]);
  not (_07314_, _07313_);
  nor (_07315_, _07314_, _07312_);
  nor (_07316_, _07315_, _07311_);
  and (_07317_, _07316_, _07304_);
  not (_07318_, _07317_);
  and (_07319_, _07301_, _07294_);
  nor (_07320_, _07319_, _07293_);
  and (_07321_, _07320_, _07318_);
  and (_07322_, _07281_, _07275_);
  nor (_07323_, _07322_, _07282_);
  not (_07324_, _07323_);
  nor (_07325_, _07324_, _07274_);
  nor (_07326_, _07258_, _07256_);
  nor (_07327_, _07326_, _07259_);
  and (_07328_, _07327_, _07269_);
  not (_07329_, _07230_);
  nor (_07330_, _07269_, _07329_);
  nor (_07331_, _07330_, _07328_);
  and (_07332_, _07331_, \oc8051_golden_model_1.B [4]);
  nor (_07333_, _07331_, \oc8051_golden_model_1.B [4]);
  nor (_07334_, _07333_, _07332_);
  nor (_07335_, _07225_, _07224_);
  nor (_07336_, _07335_, _07260_);
  and (_07337_, _07335_, _07260_);
  nor (_07338_, _07337_, _07336_);
  and (_07339_, _07338_, _07269_);
  nor (_07340_, _07269_, _07223_);
  or (_07341_, _07340_, _07339_);
  and (_07342_, _07341_, \oc8051_golden_model_1.B [5]);
  nor (_07343_, _07341_, \oc8051_golden_model_1.B [5]);
  nor (_07344_, _07343_, _07342_);
  and (_07345_, _07344_, _07334_);
  and (_07346_, _07345_, _07325_);
  not (_07347_, _07346_);
  nor (_07348_, _07347_, _07321_);
  and (_07349_, _07206_, \oc8051_golden_model_1.B [7]);
  and (_07350_, _07344_, _07332_);
  nor (_07351_, _07350_, _07342_);
  not (_07352_, _07351_);
  and (_07353_, _07352_, _07325_);
  or (_07354_, _07353_, _07349_);
  or (_07355_, _07354_, _07348_);
  nor (_07356_, _07355_, _07284_);
  and (_07357_, \oc8051_golden_model_1.B [0], _03498_);
  not (_07358_, _07357_);
  nor (_07359_, _07312_, _07311_);
  and (_07360_, _07359_, _07358_);
  and (_07361_, _07360_, _07314_);
  and (_07362_, _07361_, _07304_);
  and (_07363_, _07362_, _07346_);
  nor (_07364_, _07363_, _07356_);
  and (_07365_, _07364_, _07271_);
  or (_07366_, _07365_, _07025_);
  or (_07367_, _07366_, _07011_);
  nor (_07368_, _06088_, _07008_);
  and (_07369_, _06121_, _06088_);
  or (_07370_, _07369_, _07368_);
  and (_07371_, _07370_, _03759_);
  nor (_07372_, _05440_, _07008_);
  and (_07373_, _06160_, _05440_);
  or (_07374_, _07373_, _07372_);
  or (_07375_, _07374_, _04722_);
  and (_07376_, _05440_, \oc8051_golden_model_1.ACC [7]);
  or (_07377_, _07376_, _07372_);
  and (_07378_, _07377_, _04707_);
  nor (_07379_, _04707_, _07008_);
  or (_07380_, _07379_, _03850_);
  or (_07381_, _07380_, _07378_);
  and (_07382_, _07381_, _03764_);
  and (_07383_, _07382_, _07375_);
  and (_07384_, _06148_, _06088_);
  or (_07385_, _07384_, _07368_);
  and (_07386_, _07385_, _03763_);
  or (_07387_, _07386_, _03848_);
  or (_07388_, _07387_, _07383_);
  and (_07389_, _05568_, _05440_);
  or (_07390_, _07389_, _07372_);
  or (_07391_, _07390_, _04733_);
  and (_07392_, _07391_, _07388_);
  or (_07393_, _07392_, _03854_);
  or (_07394_, _07377_, _03855_);
  and (_07395_, _07394_, _03760_);
  and (_07396_, _07395_, _07393_);
  or (_07397_, _07396_, _07371_);
  and (_07398_, _07397_, _03753_);
  and (_07399_, _03919_, _03821_);
  or (_07400_, _07368_, _06147_);
  and (_07401_, _07400_, _03752_);
  and (_07402_, _07401_, _07385_);
  or (_07403_, _07402_, _07399_);
  or (_07404_, _07403_, _07398_);
  not (_07405_, _07399_);
  and (_07406_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_07407_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_07408_, _07407_, _07406_);
  and (_07409_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_07410_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_07411_, _07410_, _07012_);
  nor (_07412_, _07411_, _07408_);
  and (_07413_, _07412_, _07409_);
  nor (_07414_, _07413_, _07408_);
  and (_07415_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_07416_, _07410_, _07415_);
  and (_07417_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_07418_, _07417_, _07406_);
  nor (_07419_, _07418_, _07416_);
  not (_07420_, _07419_);
  nor (_07421_, _07420_, _07414_);
  and (_07422_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_07423_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_07424_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_07425_, _07424_, _07423_);
  nor (_07426_, _07424_, _07423_);
  nor (_07427_, _07426_, _07425_);
  and (_07428_, _07427_, _07422_);
  nor (_07429_, _07427_, _07422_);
  nor (_07430_, _07429_, _07428_);
  and (_07431_, _07420_, _07414_);
  nor (_07432_, _07431_, _07421_);
  and (_07433_, _07432_, _07430_);
  nor (_07434_, _07433_, _07421_);
  not (_07435_, _07410_);
  and (_07436_, _07435_, _07415_);
  and (_07437_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_07438_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_07439_, _07438_, _07423_);
  and (_07440_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_07441_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_07442_, _07441_, _07440_);
  nor (_07443_, _07442_, _07439_);
  and (_07444_, _07443_, _07437_);
  nor (_07445_, _07443_, _07437_);
  nor (_07446_, _07445_, _07444_);
  and (_07447_, _07446_, _07436_);
  nor (_07448_, _07446_, _07436_);
  nor (_07449_, _07448_, _07447_);
  not (_07450_, _07449_);
  nor (_07451_, _07450_, _07434_);
  and (_07452_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_07453_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_07454_, _07453_, _07452_);
  nor (_07455_, _07428_, _07425_);
  and (_07456_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_07457_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_07458_, _07457_, _07456_);
  nor (_07459_, _07457_, _07456_);
  nor (_07460_, _07459_, _07458_);
  not (_07461_, _07460_);
  nor (_07462_, _07461_, _07455_);
  and (_07463_, _07461_, _07455_);
  nor (_07464_, _07463_, _07462_);
  and (_07465_, _07464_, _07454_);
  nor (_07466_, _07464_, _07454_);
  nor (_07467_, _07466_, _07465_);
  and (_07468_, _07450_, _07434_);
  nor (_07469_, _07468_, _07451_);
  and (_07470_, _07469_, _07467_);
  nor (_07471_, _07470_, _07451_);
  nor (_07472_, _07444_, _07439_);
  and (_07473_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_07474_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_07475_, _07474_, _07473_);
  nor (_07476_, _07474_, _07473_);
  nor (_07477_, _07476_, _07475_);
  not (_07478_, _07477_);
  nor (_07479_, _07478_, _07472_);
  and (_07480_, _07478_, _07472_);
  nor (_07481_, _07480_, _07479_);
  and (_07482_, _07481_, _07458_);
  nor (_07483_, _07481_, _07458_);
  nor (_07484_, _07483_, _07482_);
  nor (_07485_, _07447_, _07416_);
  and (_07486_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_07487_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_07488_, _07438_, _07487_);
  nor (_07489_, _07438_, _07487_);
  nor (_07490_, _07489_, _07488_);
  and (_07491_, _07490_, _07486_);
  nor (_07492_, _07490_, _07486_);
  nor (_07493_, _07492_, _07491_);
  not (_07494_, _07493_);
  nor (_07495_, _07494_, _07485_);
  and (_07496_, _07494_, _07485_);
  nor (_07497_, _07496_, _07495_);
  and (_07498_, _07497_, _07484_);
  nor (_07499_, _07497_, _07484_);
  nor (_07500_, _07499_, _07498_);
  not (_07501_, _07500_);
  nor (_07502_, _07501_, _07471_);
  nor (_07503_, _07465_, _07462_);
  not (_07504_, _07503_);
  and (_07505_, _07501_, _07471_);
  nor (_07506_, _07505_, _07502_);
  and (_07507_, _07506_, _07504_);
  nor (_07508_, _07507_, _07502_);
  nor (_07509_, _07482_, _07479_);
  not (_07510_, _07509_);
  nor (_07511_, _07498_, _07495_);
  not (_07512_, _07511_);
  and (_07513_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_07514_, _07438_, _07513_);
  and (_07515_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_07516_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_07517_, _07516_, _07515_);
  nor (_07518_, _07517_, _07514_);
  nor (_07519_, _07491_, _07488_);
  and (_07520_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_07521_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_07522_, _07521_, _07520_);
  nor (_07523_, _07521_, _07520_);
  nor (_07524_, _07523_, _07522_);
  not (_07525_, _07524_);
  nor (_07526_, _07525_, _07519_);
  and (_07527_, _07525_, _07519_);
  nor (_07528_, _07527_, _07526_);
  and (_07529_, _07528_, _07475_);
  nor (_07530_, _07528_, _07475_);
  nor (_07531_, _07530_, _07529_);
  and (_07532_, _07531_, _07518_);
  nor (_07533_, _07531_, _07518_);
  nor (_07534_, _07533_, _07532_);
  and (_07535_, _07534_, _07512_);
  nor (_07536_, _07534_, _07512_);
  nor (_07537_, _07536_, _07535_);
  and (_07538_, _07537_, _07510_);
  nor (_07539_, _07537_, _07510_);
  nor (_07540_, _07539_, _07538_);
  not (_07541_, _07540_);
  nor (_07542_, _07541_, _07508_);
  nor (_07543_, _07538_, _07535_);
  nor (_07544_, _07529_, _07526_);
  not (_07545_, _07544_);
  and (_07546_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_07547_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_07548_, _07547_, _07546_);
  nor (_07549_, _07547_, _07546_);
  nor (_07550_, _07549_, _07548_);
  and (_07551_, _07550_, _07514_);
  nor (_07552_, _07550_, _07514_);
  nor (_07553_, _07552_, _07551_);
  and (_07554_, _07553_, _07522_);
  nor (_07555_, _07553_, _07522_);
  nor (_07556_, _07555_, _07554_);
  and (_07557_, _07556_, _07513_);
  nor (_07558_, _07556_, _07513_);
  nor (_07559_, _07558_, _07557_);
  and (_07560_, _07559_, _07532_);
  nor (_07561_, _07559_, _07532_);
  nor (_07562_, _07561_, _07560_);
  and (_07563_, _07562_, _07545_);
  nor (_07564_, _07562_, _07545_);
  nor (_07565_, _07564_, _07563_);
  not (_07566_, _07565_);
  nor (_07567_, _07566_, _07543_);
  and (_07568_, _07566_, _07543_);
  nor (_07569_, _07568_, _07567_);
  and (_07570_, _07569_, _07542_);
  nor (_07571_, _07563_, _07560_);
  nor (_07572_, _07554_, _07551_);
  not (_07573_, _07572_);
  and (_07574_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_07575_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_07576_, _07575_, _07574_);
  nor (_07577_, _07575_, _07574_);
  nor (_07578_, _07577_, _07576_);
  and (_07579_, _07578_, _07548_);
  nor (_07580_, _07578_, _07548_);
  nor (_07581_, _07580_, _07579_);
  and (_07582_, _07581_, _07557_);
  nor (_07583_, _07581_, _07557_);
  nor (_07584_, _07583_, _07582_);
  and (_07585_, _07584_, _07573_);
  nor (_07586_, _07584_, _07573_);
  nor (_07587_, _07586_, _07585_);
  not (_07588_, _07587_);
  nor (_07589_, _07588_, _07571_);
  and (_07590_, _07588_, _07571_);
  nor (_07591_, _07590_, _07589_);
  and (_07592_, _07591_, _07567_);
  nor (_07593_, _07591_, _07567_);
  nor (_07594_, _07593_, _07592_);
  and (_07595_, _07594_, _07570_);
  nor (_07596_, _07594_, _07570_);
  nor (_07597_, _07596_, _07595_);
  and (_07598_, _07410_, _07049_);
  and (_07599_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_07600_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_07601_, _07600_, _07407_);
  nor (_07602_, _07601_, _07598_);
  and (_07603_, _07602_, _07599_);
  nor (_07604_, _07603_, _07598_);
  not (_07605_, _07604_);
  nor (_07606_, _07412_, _07409_);
  nor (_07607_, _07606_, _07413_);
  and (_07608_, _07607_, _07605_);
  and (_07609_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_07610_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_07611_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_07612_, _07611_, _07610_);
  nor (_07613_, _07611_, _07610_);
  nor (_07614_, _07613_, _07612_);
  and (_07615_, _07614_, _07609_);
  nor (_07616_, _07614_, _07609_);
  nor (_07617_, _07616_, _07615_);
  nor (_07618_, _07607_, _07605_);
  nor (_07619_, _07618_, _07608_);
  and (_07620_, _07619_, _07617_);
  nor (_07621_, _07620_, _07608_);
  nor (_07622_, _07432_, _07430_);
  nor (_07623_, _07622_, _07433_);
  not (_07624_, _07623_);
  nor (_07625_, _07624_, _07621_);
  and (_07626_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_07627_, _07626_, _07453_);
  nor (_07628_, _07615_, _07612_);
  nor (_07629_, _07453_, _07452_);
  nor (_07630_, _07629_, _07454_);
  not (_07631_, _07630_);
  nor (_07632_, _07631_, _07628_);
  and (_07633_, _07631_, _07628_);
  nor (_07634_, _07633_, _07632_);
  and (_07635_, _07634_, _07627_);
  nor (_07636_, _07634_, _07627_);
  nor (_07637_, _07636_, _07635_);
  and (_07638_, _07624_, _07621_);
  nor (_07639_, _07638_, _07625_);
  and (_07640_, _07639_, _07637_);
  nor (_07641_, _07640_, _07625_);
  nor (_07642_, _07469_, _07467_);
  nor (_07643_, _07642_, _07470_);
  not (_07644_, _07643_);
  nor (_07645_, _07644_, _07641_);
  nor (_07646_, _07635_, _07632_);
  not (_07647_, _07646_);
  and (_07648_, _07644_, _07641_);
  nor (_07649_, _07648_, _07645_);
  and (_07650_, _07649_, _07647_);
  nor (_07651_, _07650_, _07645_);
  nor (_07652_, _07506_, _07504_);
  nor (_07653_, _07652_, _07507_);
  not (_07654_, _07653_);
  nor (_07655_, _07654_, _07651_);
  and (_07656_, _07541_, _07508_);
  nor (_07657_, _07656_, _07542_);
  and (_07658_, _07657_, _07655_);
  nor (_07659_, _07569_, _07542_);
  nor (_07660_, _07659_, _07570_);
  nand (_07661_, _07660_, _07658_);
  and (_07662_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_07663_, _07662_, _07049_);
  and (_07664_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_07665_, _07662_, _07049_);
  nor (_07666_, _07665_, _07663_);
  and (_07667_, _07666_, _07664_);
  nor (_07668_, _07667_, _07663_);
  not (_07669_, _07668_);
  nor (_07670_, _07602_, _07599_);
  nor (_07671_, _07670_, _07603_);
  and (_07672_, _07671_, _07669_);
  and (_07673_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_07674_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_07675_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_07676_, _07675_, _07674_);
  nor (_07677_, _07675_, _07674_);
  nor (_07678_, _07677_, _07676_);
  and (_07679_, _07678_, _07673_);
  nor (_07680_, _07678_, _07673_);
  nor (_07681_, _07680_, _07679_);
  nor (_07682_, _07671_, _07669_);
  nor (_07683_, _07682_, _07672_);
  and (_07684_, _07683_, _07681_);
  nor (_07685_, _07684_, _07672_);
  not (_07686_, _07685_);
  nor (_07687_, _07619_, _07617_);
  nor (_07688_, _07687_, _07620_);
  and (_07689_, _07688_, _07686_);
  nor (_07690_, _07679_, _07676_);
  and (_07691_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_07692_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_07693_, _07692_, _07691_);
  nor (_07694_, _07693_, _07627_);
  not (_07695_, _07694_);
  nor (_07696_, _07695_, _07690_);
  and (_07697_, _07695_, _07690_);
  nor (_07698_, _07697_, _07696_);
  nor (_07699_, _07688_, _07686_);
  nor (_07700_, _07699_, _07689_);
  and (_07701_, _07700_, _07698_);
  nor (_07702_, _07701_, _07689_);
  nor (_07703_, _07639_, _07637_);
  nor (_07704_, _07703_, _07640_);
  not (_07705_, _07704_);
  nor (_07706_, _07705_, _07702_);
  and (_07707_, _07705_, _07702_);
  nor (_07708_, _07707_, _07706_);
  and (_07709_, _07708_, _07696_);
  nor (_07710_, _07709_, _07706_);
  nor (_07711_, _07649_, _07647_);
  nor (_07712_, _07711_, _07650_);
  not (_07713_, _07712_);
  nor (_07714_, _07713_, _07710_);
  and (_07715_, _07654_, _07651_);
  nor (_07716_, _07715_, _07655_);
  and (_07717_, _07716_, _07714_);
  nor (_07718_, _07657_, _07655_);
  nor (_07719_, _07718_, _07658_);
  and (_07720_, _07719_, _07717_);
  nor (_07721_, _07719_, _07717_);
  nor (_07722_, _07721_, _07720_);
  and (_07723_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_07724_, _07723_, _07123_);
  and (_07725_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_07726_, _07723_, _07123_);
  nor (_07727_, _07726_, _07724_);
  and (_07728_, _07727_, _07725_);
  nor (_07729_, _07728_, _07724_);
  not (_07730_, _07729_);
  nor (_07731_, _07666_, _07664_);
  nor (_07732_, _07731_, _07667_);
  and (_07733_, _07732_, _07730_);
  and (_07734_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_07735_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_07736_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_07737_, _07736_, _07735_);
  nor (_07738_, _07736_, _07735_);
  nor (_07739_, _07738_, _07737_);
  and (_07740_, _07739_, _07734_);
  nor (_07741_, _07739_, _07734_);
  nor (_07742_, _07741_, _07740_);
  nor (_07743_, _07732_, _07730_);
  nor (_07744_, _07743_, _07733_);
  and (_07745_, _07744_, _07742_);
  nor (_07746_, _07745_, _07733_);
  not (_07747_, _07746_);
  nor (_07748_, _07683_, _07681_);
  nor (_07749_, _07748_, _07684_);
  and (_07750_, _07749_, _07747_);
  not (_07751_, _07626_);
  nor (_07752_, _07740_, _07737_);
  nor (_07753_, _07752_, _07751_);
  and (_07754_, _07752_, _07751_);
  nor (_07755_, _07754_, _07753_);
  nor (_07756_, _07749_, _07747_);
  nor (_07757_, _07756_, _07750_);
  and (_07758_, _07757_, _07755_);
  nor (_07759_, _07758_, _07750_);
  not (_07760_, _07759_);
  nor (_07761_, _07700_, _07698_);
  nor (_07762_, _07761_, _07701_);
  and (_07763_, _07762_, _07760_);
  nor (_07764_, _07762_, _07760_);
  nor (_07765_, _07764_, _07763_);
  and (_07766_, _07765_, _07753_);
  nor (_07767_, _07766_, _07763_);
  nor (_07768_, _07708_, _07696_);
  nor (_07769_, _07768_, _07709_);
  not (_07770_, _07769_);
  nor (_07771_, _07770_, _07767_);
  and (_07772_, _07713_, _07710_);
  nor (_07773_, _07772_, _07714_);
  and (_07774_, _07773_, _07771_);
  nor (_07775_, _07716_, _07714_);
  nor (_07776_, _07775_, _07717_);
  nand (_07777_, _07776_, _07774_);
  or (_07778_, _07776_, _07774_);
  and (_07779_, _07778_, _07777_);
  and (_07780_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_07781_, _07780_, _07129_);
  and (_07782_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07783_, _07780_, _07129_);
  nor (_07784_, _07783_, _07781_);
  and (_07785_, _07784_, _07782_);
  nor (_07786_, _07785_, _07781_);
  not (_07787_, _07786_);
  nor (_07788_, _07727_, _07725_);
  nor (_07789_, _07788_, _07728_);
  and (_07790_, _07789_, _07787_);
  and (_07791_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_07792_, _07791_, _07736_);
  and (_07793_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_07794_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_07795_, _07794_, _07793_);
  nor (_07796_, _07795_, _07792_);
  nor (_07797_, _07789_, _07787_);
  nor (_07798_, _07797_, _07790_);
  and (_07799_, _07798_, _07796_);
  nor (_07800_, _07799_, _07790_);
  not (_07801_, _07800_);
  nor (_07802_, _07744_, _07742_);
  nor (_07803_, _07802_, _07745_);
  and (_07804_, _07803_, _07801_);
  nor (_07805_, _07803_, _07801_);
  nor (_07806_, _07805_, _07804_);
  and (_07807_, _07806_, _07792_);
  nor (_07808_, _07807_, _07804_);
  not (_07809_, _07808_);
  nor (_07810_, _07757_, _07755_);
  nor (_07811_, _07810_, _07758_);
  and (_07812_, _07811_, _07809_);
  nor (_07813_, _07765_, _07753_);
  nor (_07814_, _07813_, _07766_);
  and (_07815_, _07814_, _07812_);
  and (_07816_, _07770_, _07767_);
  nor (_07817_, _07816_, _07771_);
  and (_07818_, _07817_, _07815_);
  nor (_07819_, _07773_, _07771_);
  nor (_07820_, _07819_, _07774_);
  and (_07821_, _07820_, _07818_);
  nor (_07822_, _07820_, _07818_);
  nor (_07823_, _07822_, _07821_);
  and (_07824_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_07825_, _07824_, _07242_);
  and (_07826_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_07827_, _07824_, _07242_);
  nor (_07828_, _07827_, _07825_);
  and (_07829_, _07828_, _07826_);
  nor (_07830_, _07829_, _07825_);
  not (_07831_, _07830_);
  nor (_07832_, _07784_, _07782_);
  nor (_07833_, _07832_, _07785_);
  and (_07834_, _07833_, _07831_);
  nor (_07835_, _07833_, _07831_);
  nor (_07836_, _07835_, _07834_);
  and (_07837_, _07836_, _07791_);
  nor (_07838_, _07837_, _07834_);
  not (_07839_, _07838_);
  nor (_07840_, _07798_, _07796_);
  nor (_07841_, _07840_, _07799_);
  and (_07842_, _07841_, _07839_);
  nor (_07843_, _07806_, _07792_);
  nor (_07844_, _07843_, _07807_);
  and (_07845_, _07844_, _07842_);
  nor (_07846_, _07811_, _07809_);
  nor (_07847_, _07846_, _07812_);
  and (_07848_, _07847_, _07845_);
  nor (_07849_, _07814_, _07812_);
  nor (_07850_, _07849_, _07815_);
  and (_07851_, _07850_, _07848_);
  nor (_07852_, _07817_, _07815_);
  nor (_07853_, _07852_, _07818_);
  and (_07854_, _07853_, _07851_);
  and (_07855_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_07856_, _07824_, _07855_);
  nor (_07857_, _07828_, _07826_);
  nor (_07858_, _07857_, _07829_);
  and (_07859_, _07858_, _07856_);
  nor (_07860_, _07836_, _07791_);
  nor (_07861_, _07860_, _07837_);
  and (_07862_, _07861_, _07859_);
  nor (_07863_, _07841_, _07839_);
  nor (_07864_, _07863_, _07842_);
  and (_07865_, _07864_, _07862_);
  nor (_07866_, _07844_, _07842_);
  nor (_07867_, _07866_, _07845_);
  and (_07868_, _07867_, _07865_);
  nor (_07869_, _07847_, _07845_);
  nor (_07870_, _07869_, _07848_);
  and (_07871_, _07870_, _07868_);
  nor (_07872_, _07850_, _07848_);
  nor (_07873_, _07872_, _07851_);
  and (_07874_, _07873_, _07871_);
  nor (_07875_, _07853_, _07851_);
  nor (_07876_, _07875_, _07854_);
  and (_07877_, _07876_, _07874_);
  nor (_07878_, _07877_, _07854_);
  not (_07879_, _07878_);
  and (_07880_, _07879_, _07823_);
  or (_07881_, _07880_, _07821_);
  nand (_07882_, _07881_, _07779_);
  and (_07883_, _07882_, _07777_);
  not (_07884_, _07883_);
  and (_07885_, _07884_, _07722_);
  or (_07886_, _07885_, _07720_);
  or (_07887_, _07660_, _07658_);
  and (_07888_, _07887_, _07661_);
  nand (_07889_, _07888_, _07886_);
  and (_07890_, _07889_, _07661_);
  not (_07891_, _07890_);
  and (_07892_, _07891_, _07597_);
  or (_07893_, _07892_, _07595_);
  not (_07894_, _07547_);
  and (_07895_, _07894_, _07272_);
  nor (_07896_, _07895_, _07579_);
  nor (_07897_, _07585_, _07582_);
  nor (_07898_, _07897_, _07896_);
  and (_07899_, _07897_, _07896_);
  nor (_07900_, _07899_, _07898_);
  nor (_07901_, _07592_, _07589_);
  and (_07902_, _07901_, _07900_);
  nor (_07903_, _07901_, _07900_);
  or (_07904_, _07903_, _07902_);
  and (_07905_, _07904_, _07893_);
  and (_07906_, _07900_, _07589_);
  or (_07907_, _07898_, _07576_);
  or (_07908_, _07907_, _07906_);
  and (_07909_, _07900_, _07592_);
  or (_07910_, _07909_, _07908_);
  or (_07911_, _07910_, _07905_);
  or (_07912_, _07911_, _07405_);
  and (_07913_, _07912_, _03747_);
  and (_07914_, _07913_, _07404_);
  not (_07915_, _06088_);
  nor (_07916_, _06143_, _07915_);
  or (_07917_, _07916_, _07368_);
  and (_07918_, _07917_, _03746_);
  nor (_07919_, _03834_, _03724_);
  or (_07920_, _07919_, _03720_);
  not (_07921_, _03422_);
  and (_07922_, _03728_, _07921_);
  and (_07923_, _07922_, _03397_);
  not (_07924_, _07923_);
  and (_07925_, _07924_, _07920_);
  and (_07926_, _07925_, _03738_);
  not (_07927_, _07926_);
  or (_07928_, _07927_, _07918_);
  or (_07929_, _07928_, _07914_);
  and (_07930_, _06248_, _05440_);
  or (_07931_, _07372_, _03738_);
  or (_07932_, _07931_, _07930_);
  or (_07933_, _07925_, _07390_);
  and (_07934_, _07933_, _03820_);
  and (_07935_, _07934_, _07932_);
  and (_07936_, _07935_, _07929_);
  not (_07937_, _05440_);
  nor (_07938_, _06536_, _07937_);
  or (_07939_, _07938_, _07372_);
  and (_07940_, _07939_, _03455_);
  or (_07941_, _07940_, _07010_);
  or (_07942_, _07941_, _07936_);
  and (_07943_, _07942_, _07367_);
  or (_07944_, _07943_, _03903_);
  and (_07945_, _06348_, _05440_);
  or (_07946_, _07945_, _07372_);
  or (_07947_, _07946_, _04778_);
  and (_07948_, _07947_, _04790_);
  and (_07949_, _07948_, _07944_);
  and (_07950_, _06549_, _05440_);
  or (_07951_, _07950_, _07372_);
  and (_07952_, _07951_, _03897_);
  or (_07953_, _07952_, _04018_);
  or (_07954_, _07953_, _07949_);
  and (_07955_, _06557_, _05440_);
  or (_07956_, _07955_, _07372_);
  or (_07957_, _07956_, _04792_);
  and (_07958_, _07957_, _03909_);
  and (_07959_, _07958_, _07954_);
  or (_07960_, _07372_, _05571_);
  and (_07961_, _07946_, _03908_);
  and (_07962_, _07961_, _07960_);
  or (_07963_, _07962_, _07959_);
  and (_07964_, _07963_, _04785_);
  and (_07965_, _07377_, _04027_);
  and (_07966_, _07965_, _07960_);
  or (_07967_, _07966_, _03914_);
  or (_07968_, _07967_, _07964_);
  nor (_07969_, _06547_, _07937_);
  or (_07970_, _07372_, _06567_);
  or (_07971_, _07970_, _07969_);
  and (_07972_, _07971_, _06572_);
  and (_07973_, _07972_, _07968_);
  nor (_07974_, _06556_, _07937_);
  or (_07975_, _07974_, _07372_);
  and (_07976_, _07975_, _04011_);
  or (_07977_, _07976_, _03773_);
  or (_07978_, _07977_, _07973_);
  or (_07979_, _07374_, _03774_);
  and (_07980_, _07979_, _03375_);
  and (_07981_, _07980_, _07978_);
  and (_07982_, _07370_, _03374_);
  or (_07983_, _07982_, _03772_);
  or (_07984_, _07983_, _07981_);
  and (_07985_, _06077_, _05440_);
  or (_07986_, _07372_, _04060_);
  or (_07987_, _07986_, _07985_);
  and (_07988_, _07987_, _43152_);
  and (_07989_, _07988_, _07984_);
  or (_07990_, _07989_, _07009_);
  and (_40680_, _07990_, _41894_);
  nor (_07991_, _43152_, _06554_);
  and (_07992_, _03719_, _03409_);
  not (_07993_, _07992_);
  and (_07994_, _03726_, _03409_);
  nor (_07995_, _03730_, _03834_);
  nor (_07996_, _07995_, _04452_);
  nor (_07997_, _07996_, _07994_);
  and (_07998_, _07997_, _04451_);
  and (_07999_, _07998_, _07993_);
  nor (_08000_, _05568_, \oc8051_golden_model_1.ACC [7]);
  and (_08001_, _05568_, \oc8051_golden_model_1.ACC [7]);
  nor (_08002_, _08001_, _08000_);
  and (_08003_, _06065_, \oc8051_golden_model_1.ACC [6]);
  nor (_08004_, _06065_, \oc8051_golden_model_1.ACC [6]);
  nor (_08005_, _08004_, _08003_);
  and (_08006_, _05857_, \oc8051_golden_model_1.ACC [5]);
  nor (_08007_, _05857_, \oc8051_golden_model_1.ACC [5]);
  nor (_08008_, _08007_, _08006_);
  not (_08009_, _08008_);
  and (_08010_, _05950_, \oc8051_golden_model_1.ACC [4]);
  nor (_08011_, _05950_, \oc8051_golden_model_1.ACC [4]);
  nor (_08012_, _08011_, _08010_);
  and (_08013_, _05119_, \oc8051_golden_model_1.ACC [3]);
  nor (_08014_, _05119_, \oc8051_golden_model_1.ACC [3]);
  and (_08015_, _05307_, \oc8051_golden_model_1.ACC [2]);
  nor (_08016_, _05307_, \oc8051_golden_model_1.ACC [2]);
  nor (_08017_, _08016_, _08015_);
  not (_08018_, _08017_);
  and (_08019_, _04900_, \oc8051_golden_model_1.ACC [1]);
  nor (_08020_, _04900_, \oc8051_golden_model_1.ACC [1]);
  nor (_08021_, _08020_, _08019_);
  and (_08022_, _04700_, \oc8051_golden_model_1.ACC [0]);
  and (_08023_, _08022_, _08021_);
  nor (_08024_, _08023_, _08019_);
  nor (_08025_, _08024_, _08018_);
  nor (_08026_, _08025_, _08015_);
  nor (_08027_, _08026_, _08014_);
  or (_08028_, _08027_, _08013_);
  and (_08029_, _08028_, _08012_);
  nor (_08030_, _08029_, _08010_);
  nor (_08031_, _08030_, _08009_);
  or (_08032_, _08031_, _08006_);
  and (_08033_, _08032_, _08005_);
  nor (_08034_, _08033_, _08003_);
  nor (_08035_, _08034_, _08002_);
  and (_08036_, _08034_, _08002_);
  or (_08037_, _08036_, _08035_);
  and (_08038_, _08037_, _07993_);
  or (_08039_, _08038_, _07999_);
  and (_08040_, _06949_, \oc8051_golden_model_1.PSW [7]);
  and (_08041_, _08040_, _06952_);
  and (_08042_, _08040_, _06065_);
  nor (_08043_, _08042_, _05568_);
  nor (_08044_, _08043_, _08041_);
  nor (_08045_, _08044_, _06554_);
  and (_08046_, _08044_, _06554_);
  nor (_08047_, _08046_, _08045_);
  nor (_08048_, _08040_, _06065_);
  nor (_08049_, _08048_, _08042_);
  and (_08050_, _08049_, \oc8051_golden_model_1.ACC [6]);
  nor (_08051_, _08049_, _07036_);
  and (_08052_, _08049_, _07036_);
  nor (_08053_, _08052_, _08051_);
  not (_08054_, _08053_);
  and (_08055_, _06947_, _05950_);
  and (_08056_, _08055_, \oc8051_golden_model_1.PSW [7]);
  nor (_08057_, _08056_, _05857_);
  nor (_08058_, _08057_, _08040_);
  and (_08059_, _08058_, \oc8051_golden_model_1.ACC [5]);
  nor (_08060_, _08058_, _07084_);
  and (_08061_, _08058_, _07084_);
  nor (_08062_, _08061_, _08060_);
  and (_08063_, _06945_, \oc8051_golden_model_1.PSW [7]);
  and (_08064_, _08063_, _06946_);
  nor (_08065_, _08064_, _05950_);
  nor (_08066_, _08065_, _08056_);
  and (_08067_, _08066_, \oc8051_golden_model_1.ACC [4]);
  nor (_08068_, _08066_, _07090_);
  and (_08069_, _08066_, _07090_);
  nor (_08070_, _08069_, _08068_);
  not (_08071_, _08070_);
  and (_08072_, _06945_, _05307_);
  and (_08073_, _08072_, \oc8051_golden_model_1.PSW [7]);
  nor (_08074_, _08073_, _05119_);
  nor (_08075_, _08074_, _08064_);
  and (_08076_, _08075_, \oc8051_golden_model_1.ACC [3]);
  nor (_08077_, _08075_, _07184_);
  and (_08078_, _08075_, _07184_);
  nor (_08079_, _08078_, _08077_);
  nor (_08080_, _08063_, _05307_);
  nor (_08081_, _08080_, _08073_);
  and (_08082_, _08081_, \oc8051_golden_model_1.ACC [2]);
  nor (_08083_, _08081_, _07190_);
  and (_08084_, _08081_, _07190_);
  nor (_08085_, _08084_, _08083_);
  and (_08086_, _04700_, \oc8051_golden_model_1.PSW [7]);
  nor (_08087_, _08086_, _04900_);
  nor (_08088_, _08087_, _08063_);
  and (_08089_, _08088_, \oc8051_golden_model_1.ACC [1]);
  and (_08090_, _08088_, _03474_);
  nor (_08091_, _08088_, _03474_);
  nor (_08092_, _08091_, _08090_);
  nor (_08093_, _04700_, \oc8051_golden_model_1.PSW [7]);
  nor (_08094_, _08093_, _08086_);
  and (_08095_, _08094_, \oc8051_golden_model_1.ACC [0]);
  not (_08096_, _08095_);
  nor (_08097_, _08096_, _08092_);
  nor (_08098_, _08097_, _08089_);
  nor (_08099_, _08098_, _08085_);
  nor (_08100_, _08099_, _08082_);
  nor (_08101_, _08100_, _08079_);
  or (_08102_, _08101_, _08076_);
  and (_08103_, _08102_, _08071_);
  nor (_08104_, _08103_, _08067_);
  nor (_08105_, _08104_, _08062_);
  or (_08106_, _08105_, _08059_);
  and (_08107_, _08106_, _08054_);
  nor (_08108_, _08107_, _08050_);
  nor (_08109_, _08108_, _08047_);
  and (_08110_, _08108_, _08047_);
  nor (_08111_, _08110_, _08109_);
  not (_08112_, _04434_);
  nor (_08113_, _04233_, _04203_);
  and (_08114_, _08113_, _04221_);
  or (_08115_, _03825_, _03822_);
  and (_08116_, _08115_, _03382_);
  nor (_08117_, _08116_, _04616_);
  and (_08118_, _08117_, _08114_);
  and (_08119_, _08118_, _08112_);
  or (_08120_, _08119_, _08111_);
  nand (_08121_, _03387_, _03370_);
  not (_08122_, _08121_);
  and (_08123_, _08122_, _08001_);
  nor (_08124_, _05429_, _06554_);
  and (_08125_, _06549_, _05429_);
  nor (_08126_, _08125_, _08124_);
  nand (_08127_, _08126_, _03897_);
  not (_08128_, _08047_);
  nor (_08129_, _08068_, _08060_);
  nor (_08130_, _08129_, _08061_);
  and (_08131_, _08070_, _08062_);
  not (_08132_, _08131_);
  and (_08133_, _08085_, _08079_);
  and (_08134_, _08094_, _03498_);
  nor (_08135_, _08134_, _08090_);
  or (_08136_, _08135_, _08091_);
  and (_08137_, _08136_, _08133_);
  and (_08138_, _08083_, _08079_);
  or (_08139_, _08138_, _08077_);
  nor (_08140_, _08139_, _08137_);
  nor (_08141_, _08140_, _08132_);
  nor (_08142_, _08141_, _08130_);
  nor (_08143_, _08142_, _08054_);
  or (_08144_, _08143_, _08051_);
  and (_08145_, _08144_, _08128_);
  nor (_08146_, _08144_, _08128_);
  nor (_08147_, _08146_, _08145_);
  and (_08148_, _03719_, _03424_);
  nor (_08149_, _08148_, _04333_);
  and (_08150_, _03726_, _03424_);
  nor (_08151_, _07995_, _04609_);
  nor (_08152_, _08151_, _08150_);
  and (_08153_, _08152_, _08149_);
  nor (_08154_, _08153_, _08147_);
  not (_08155_, _04227_);
  nor (_08156_, _04282_, _04188_);
  and (_08157_, _08156_, _08155_);
  or (_08158_, _08157_, _05568_);
  and (_08159_, _03919_, _03766_);
  not (_08160_, _08159_);
  or (_08161_, _08160_, _06248_);
  not (_08162_, _03436_);
  nor (_08163_, _03850_, _08162_);
  not (_08164_, _08115_);
  and (_08165_, _04291_, _08164_);
  nor (_08166_, _04760_, _03831_);
  and (_08167_, _08166_, _07995_);
  and (_08168_, _08167_, _08165_);
  nor (_08169_, _08168_, _03435_);
  and (_08170_, _08169_, _05568_);
  or (_08171_, _04263_, \oc8051_golden_model_1.ACC [7]);
  nand (_08172_, _04263_, \oc8051_golden_model_1.ACC [7]);
  nand (_08173_, _08172_, _08171_);
  nor (_08174_, _08173_, _08169_);
  or (_08175_, _08174_, _08159_);
  or (_08176_, _08175_, _08170_);
  and (_08177_, _08176_, _08163_);
  and (_08178_, _08177_, _08161_);
  and (_08179_, _03919_, _03762_);
  and (_08180_, _06160_, _05429_);
  nor (_08181_, _08180_, _08124_);
  nor (_08182_, _08181_, _04722_);
  or (_08183_, _08182_, _08179_);
  or (_08184_, _08183_, _08178_);
  nor (_08185_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_08186_, _08185_, _07184_);
  and (_08187_, _08186_, _07055_);
  and (_08188_, _08187_, \oc8051_golden_model_1.ACC [6]);
  and (_08189_, _08188_, \oc8051_golden_model_1.ACC [7]);
  nor (_08190_, _08188_, \oc8051_golden_model_1.ACC [7]);
  nor (_08191_, _08190_, _08189_);
  and (_08192_, _08186_, \oc8051_golden_model_1.ACC [4]);
  nor (_08193_, _08192_, \oc8051_golden_model_1.ACC [5]);
  nor (_08194_, _08193_, _08187_);
  nor (_08195_, _08187_, \oc8051_golden_model_1.ACC [6]);
  nor (_08196_, _08195_, _08188_);
  nor (_08197_, _08196_, _08194_);
  not (_08198_, _08197_);
  and (_08199_, _08198_, _08191_);
  nor (_08200_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_08201_, _08200_, _08197_);
  nor (_08202_, _08201_, _08191_);
  nor (_08203_, _08202_, _08199_);
  not (_08204_, _08203_);
  nand (_08205_, _08204_, _08179_);
  and (_08206_, _08205_, _03856_);
  and (_08207_, _08206_, _08184_);
  nor (_08208_, _06096_, _06554_);
  and (_08209_, _06148_, _06096_);
  nor (_08210_, _08209_, _08208_);
  nor (_08211_, _08210_, _03764_);
  not (_08212_, _08157_);
  and (_08213_, _05568_, _05429_);
  nor (_08214_, _08213_, _08124_);
  nor (_08215_, _08214_, _04733_);
  or (_08216_, _08215_, _08212_);
  or (_08217_, _08216_, _08211_);
  or (_08218_, _08217_, _08207_);
  and (_08219_, _08218_, _08158_);
  or (_08220_, _08219_, _04738_);
  or (_08221_, _06248_, _04739_);
  and (_08222_, _08221_, _03855_);
  and (_08223_, _08222_, _08220_);
  and (_08224_, _03919_, _03757_);
  nor (_08225_, _05570_, _03855_);
  or (_08226_, _08225_, _08224_);
  or (_08227_, _08226_, _08223_);
  nand (_08228_, _08224_, _07184_);
  and (_08229_, _08228_, _08227_);
  or (_08230_, _08229_, _03759_);
  and (_08231_, _06121_, _06096_);
  nor (_08232_, _08231_, _08208_);
  nand (_08233_, _08232_, _03759_);
  and (_08234_, _08233_, _03753_);
  and (_08235_, _08234_, _08230_);
  and (_08236_, _08209_, _06147_);
  nor (_08237_, _08236_, _08208_);
  nor (_08238_, _08237_, _03753_);
  or (_08239_, _08238_, _07399_);
  or (_08240_, _08239_, _08235_);
  nor (_08241_, _07873_, _07871_);
  nor (_08242_, _08241_, _07874_);
  or (_08243_, _08242_, _07405_);
  and (_08244_, _08243_, _08240_);
  and (_08245_, _08244_, _08153_);
  or (_08246_, _08245_, _08154_);
  or (_08247_, _08246_, _04330_);
  not (_08248_, _04330_);
  and (_08249_, _06972_, \oc8051_golden_model_1.PSW [7]);
  nor (_08250_, _08249_, _06596_);
  and (_08251_, _08249_, _06596_);
  nor (_08252_, _08251_, _08250_);
  and (_08253_, _08252_, \oc8051_golden_model_1.ACC [7]);
  nor (_08254_, _08252_, \oc8051_golden_model_1.ACC [7]);
  nor (_08255_, _08254_, _08253_);
  not (_08256_, _08255_);
  and (_08257_, _06971_, \oc8051_golden_model_1.PSW [7]);
  nor (_08258_, _08257_, _06641_);
  nor (_08259_, _08258_, _08249_);
  nor (_08260_, _08259_, _07036_);
  and (_08261_, _06967_, _06969_);
  and (_08262_, _08261_, \oc8051_golden_model_1.PSW [7]);
  nor (_08263_, _08262_, _06968_);
  nor (_08264_, _08263_, _08257_);
  and (_08265_, _08264_, _07084_);
  nor (_08266_, _08264_, _07084_);
  and (_08267_, _06963_, \oc8051_golden_model_1.PSW [7]);
  and (_08268_, _08267_, _06966_);
  nor (_08269_, _08268_, _06969_);
  nor (_08270_, _08269_, _08262_);
  nor (_08271_, _08270_, _07090_);
  nor (_08272_, _08271_, _08266_);
  nor (_08273_, _08272_, _08265_);
  nor (_08274_, _08266_, _08265_);
  not (_08275_, _08274_);
  and (_08276_, _08270_, _07090_);
  or (_08277_, _08276_, _08271_);
  or (_08278_, _08277_, _08275_);
  and (_08279_, _06963_, _06965_);
  and (_08280_, _08279_, \oc8051_golden_model_1.PSW [7]);
  nor (_08281_, _08280_, _06964_);
  nor (_08282_, _08281_, _08268_);
  nor (_08283_, _08282_, _07184_);
  and (_08284_, _08282_, _07184_);
  nor (_08285_, _08284_, _08283_);
  nor (_08286_, _08267_, _06965_);
  nor (_08287_, _08286_, _08280_);
  nor (_08288_, _08287_, _07190_);
  and (_08289_, _08287_, _07190_);
  nor (_08290_, _08289_, _08288_);
  and (_08291_, _08290_, _08285_);
  and (_08292_, _06962_, \oc8051_golden_model_1.PSW [7]);
  nor (_08293_, _08292_, _06961_);
  nor (_08294_, _08293_, _08267_);
  nor (_08295_, _08294_, _03474_);
  and (_08296_, _08294_, _03474_);
  not (_08297_, \oc8051_golden_model_1.PSW [7]);
  and (_08298_, _06733_, _08297_);
  nor (_08299_, _08298_, _08292_);
  and (_08300_, _08299_, _03498_);
  nor (_08301_, _08300_, _08296_);
  or (_08302_, _08301_, _08295_);
  nand (_08303_, _08302_, _08291_);
  and (_08304_, _08288_, _08285_);
  nor (_08305_, _08304_, _08283_);
  and (_08306_, _08305_, _08303_);
  nor (_08307_, _08306_, _08278_);
  nor (_08308_, _08307_, _08273_);
  and (_08309_, _08259_, _07036_);
  nor (_08310_, _08260_, _08309_);
  not (_08311_, _08310_);
  nor (_08312_, _08311_, _08308_);
  or (_08313_, _08312_, _08260_);
  and (_08314_, _08313_, _08256_);
  nor (_08315_, _08313_, _08256_);
  or (_08316_, _08315_, _08314_);
  or (_08317_, _08316_, _08248_);
  and (_08318_, _08317_, _08247_);
  or (_08319_, _08318_, _03883_);
  and (_08320_, _03919_, _03424_);
  not (_08321_, _08320_);
  not (_08322_, _06068_);
  and (_08323_, _05956_, \oc8051_golden_model_1.PSW [7]);
  and (_08324_, _08323_, _08322_);
  nor (_08325_, _08324_, _05570_);
  and (_08326_, _08324_, _05570_);
  nor (_08327_, _08326_, _08325_);
  and (_08328_, _08327_, \oc8051_golden_model_1.ACC [7]);
  nor (_08329_, _08327_, \oc8051_golden_model_1.ACC [7]);
  nor (_08330_, _08329_, _08328_);
  not (_08331_, _08330_);
  nor (_08332_, _08323_, _08322_);
  nor (_08333_, _08332_, _08324_);
  nor (_08334_, _08333_, _07036_);
  not (_08335_, _05859_);
  not (_08336_, _05953_);
  and (_08337_, _05767_, \oc8051_golden_model_1.PSW [7]);
  and (_08338_, _08337_, _08336_);
  nor (_08339_, _08338_, _08335_);
  nor (_08340_, _08339_, _08323_);
  and (_08341_, _08340_, _07084_);
  nor (_08342_, _08340_, _07084_);
  nor (_08343_, _08337_, _08336_);
  nor (_08344_, _08343_, _08338_);
  nor (_08345_, _08344_, _07090_);
  nor (_08346_, _08345_, _08342_);
  nor (_08347_, _08346_, _08341_);
  nor (_08348_, _08342_, _08341_);
  not (_08349_, _08348_);
  and (_08350_, _08344_, _07090_);
  or (_08351_, _08350_, _08345_);
  or (_08352_, _08351_, _08349_);
  and (_08353_, _05766_, \oc8051_golden_model_1.PSW [7]);
  nor (_08354_, _08353_, _05622_);
  nor (_08355_, _08354_, _08337_);
  nor (_08356_, _08355_, _07184_);
  and (_08357_, _08355_, _07184_);
  nor (_08358_, _08357_, _08356_);
  and (_08359_, _05717_, \oc8051_golden_model_1.PSW [7]);
  nor (_08360_, _08359_, _05765_);
  nor (_08361_, _08360_, _08353_);
  nor (_08362_, _08361_, _07190_);
  and (_08363_, _08361_, _07190_);
  nor (_08364_, _08363_, _08362_);
  and (_08365_, _08364_, _08358_);
  not (_08366_, _05669_);
  nor (_08367_, _05716_, _08297_);
  nor (_08368_, _08367_, _08366_);
  nor (_08369_, _08368_, _08359_);
  nor (_08370_, _08369_, _03474_);
  and (_08371_, _08369_, _03474_);
  and (_08372_, _05716_, _08297_);
  nor (_08373_, _08372_, _08367_);
  and (_08374_, _08373_, _03498_);
  nor (_08375_, _08374_, _08371_);
  or (_08376_, _08375_, _08370_);
  and (_08377_, _08376_, _08365_);
  and (_08378_, _08362_, _08358_);
  or (_08379_, _08378_, _08356_);
  nor (_08380_, _08379_, _08377_);
  nor (_08381_, _08380_, _08352_);
  nor (_08382_, _08381_, _08347_);
  and (_08383_, _08333_, _07036_);
  nor (_08384_, _08334_, _08383_);
  not (_08385_, _08384_);
  nor (_08386_, _08385_, _08382_);
  or (_08387_, _08386_, _08334_);
  and (_08388_, _08387_, _08331_);
  nor (_08389_, _08387_, _08331_);
  or (_08390_, _08389_, _08388_);
  or (_08391_, _08390_, _03888_);
  and (_08392_, _08391_, _08321_);
  and (_08393_, _08392_, _08319_);
  and (_08394_, _05457_, \oc8051_golden_model_1.PSW [7]);
  and (_08395_, _08394_, _05449_);
  and (_08396_, _08395_, _05435_);
  and (_08397_, _08396_, _05232_);
  nor (_08398_, _08397_, _05421_);
  and (_08399_, _08395_, _05419_);
  and (_08400_, _08399_, _05426_);
  and (_08401_, _08400_, _03811_);
  or (_08402_, _08401_, _08398_);
  nor (_08403_, _08402_, _06554_);
  and (_08404_, _08402_, _06554_);
  nor (_08405_, _08404_, _08403_);
  not (_08406_, _08405_);
  nor (_08407_, _08396_, _05232_);
  nor (_08408_, _08407_, _08397_);
  nor (_08409_, _08408_, _07036_);
  and (_08410_, _08408_, _07036_);
  nor (_08411_, _08409_, _08410_);
  nor (_08412_, _08399_, _05426_);
  nor (_08413_, _08412_, _08396_);
  nor (_08414_, _08413_, _07084_);
  and (_08415_, _08413_, _07084_);
  nor (_08416_, _08415_, _08414_);
  not (_08417_, _08416_);
  nor (_08418_, _08395_, _05419_);
  nor (_08419_, _08418_, _08399_);
  and (_08420_, _08419_, _07090_);
  nor (_08421_, _08419_, _07090_);
  or (_08422_, _08421_, _08420_);
  or (_08423_, _08422_, _08417_);
  nor (_08424_, _06142_, _03812_);
  nor (_08425_, _08424_, _08395_);
  nor (_08426_, _08425_, _07184_);
  and (_08427_, _08425_, _07184_);
  nor (_08428_, _08427_, _08426_);
  nor (_08429_, _08394_, _05243_);
  nor (_08430_, _08429_, _06142_);
  nor (_08431_, _08430_, _07190_);
  and (_08432_, _08430_, _07190_);
  nor (_08433_, _08432_, _08431_);
  and (_08434_, _08433_, _08428_);
  nor (_08435_, _03715_, _08297_);
  nor (_08436_, _08435_, _04835_);
  nor (_08437_, _08436_, _08394_);
  nor (_08438_, _08437_, _03474_);
  and (_08439_, _08437_, _03474_);
  and (_08440_, _03715_, _08297_);
  nor (_08441_, _08440_, _08435_);
  and (_08442_, _08441_, _03498_);
  nor (_08443_, _08442_, _08439_);
  or (_08444_, _08443_, _08438_);
  nand (_08445_, _08444_, _08434_);
  nor (_08446_, _08431_, _08426_);
  or (_08447_, _08446_, _08427_);
  and (_08448_, _08447_, _08445_);
  nor (_08449_, _08448_, _08423_);
  nor (_08450_, _08421_, _08414_);
  nor (_08451_, _08450_, _08415_);
  nor (_08452_, _08451_, _08449_);
  not (_08453_, _08452_);
  and (_08454_, _08453_, _08411_);
  or (_08455_, _08454_, _08409_);
  and (_08456_, _08455_, _08406_);
  nor (_08457_, _08455_, _08406_);
  or (_08458_, _08457_, _08456_);
  and (_08459_, _08458_, _08320_);
  or (_08460_, _08459_, _03425_);
  or (_08461_, _08460_, _08393_);
  or (_08462_, _03647_, _03426_);
  and (_08463_, _08462_, _03747_);
  and (_08464_, _08463_, _08461_);
  not (_08465_, _06096_);
  nor (_08466_, _06143_, _08465_);
  nor (_08467_, _08466_, _08208_);
  nor (_08468_, _08467_, _03747_);
  or (_08469_, _08468_, _07927_);
  or (_08470_, _08469_, _08464_);
  and (_08471_, _06248_, _05429_);
  nor (_08472_, _08471_, _08124_);
  nand (_08473_, _08472_, _03737_);
  not (_08474_, _07925_);
  nand (_08475_, _08214_, _08474_);
  and (_08476_, _08475_, _03820_);
  and (_08477_, _08476_, _08473_);
  and (_08478_, _08477_, _08470_);
  not (_08479_, _05429_);
  nor (_08480_, _06536_, _08479_);
  nor (_08481_, _08480_, _08124_);
  nor (_08482_, _08481_, _03820_);
  or (_08483_, _08482_, _07010_);
  or (_08484_, _08483_, _08478_);
  not (_08485_, _07024_);
  nand (_08486_, _08485_, _07010_);
  and (_08487_, _08486_, _03479_);
  and (_08488_, _08487_, _08484_);
  and (_08489_, _03647_, _03469_);
  or (_08490_, _08489_, _03903_);
  or (_08491_, _08490_, _08488_);
  and (_08492_, _03919_, _03400_);
  not (_08493_, _08492_);
  and (_08494_, _06348_, _05429_);
  nor (_08495_, _08494_, _08124_);
  nand (_08496_, _08495_, _03903_);
  and (_08497_, _08496_, _08493_);
  and (_08498_, _08497_, _08491_);
  and (_08499_, _08492_, _03647_);
  and (_08500_, _03767_, _03404_);
  and (_08501_, _03828_, _03404_);
  nor (_08502_, _08501_, _08500_);
  not (_08503_, _08502_);
  or (_08504_, _08503_, _08499_);
  or (_08505_, _08504_, _08498_);
  and (_08506_, _03834_, _03404_);
  nor (_08507_, _08506_, _04400_);
  and (_08508_, _08507_, _04395_);
  or (_08509_, _08502_, _08002_);
  and (_08510_, _08509_, _08508_);
  and (_08511_, _08510_, _08505_);
  and (_08512_, _03719_, _03404_);
  not (_08513_, _08512_);
  and (_08514_, _08513_, _08508_);
  not (_08515_, _08514_);
  or (_08516_, _08512_, _08002_);
  and (_08517_, _08516_, _08515_);
  or (_08518_, _08517_, _08511_);
  and (_08519_, _03736_, _03404_);
  not (_08520_, _08519_);
  or (_08521_, _08513_, _08002_);
  and (_08522_, _08521_, _08520_);
  and (_08523_, _08522_, _08518_);
  nor (_08524_, _06248_, \oc8051_golden_model_1.ACC [7]);
  and (_08525_, _06248_, \oc8051_golden_model_1.ACC [7]);
  nor (_08526_, _08525_, _08524_);
  and (_08527_, _08526_, _08519_);
  or (_08528_, _08527_, _04016_);
  or (_08529_, _08528_, _08523_);
  and (_08530_, _03919_, _03404_);
  not (_08531_, _08530_);
  or (_08532_, _06557_, _04017_);
  and (_08533_, _08532_, _08531_);
  and (_08534_, _08533_, _08529_);
  nor (_08535_, _03647_, \oc8051_golden_model_1.ACC [7]);
  and (_08536_, _03647_, \oc8051_golden_model_1.ACC [7]);
  nor (_08537_, _08536_, _08535_);
  and (_08538_, _08530_, _08537_);
  or (_08539_, _08538_, _03897_);
  or (_08540_, _08539_, _08534_);
  and (_08541_, _08540_, _08127_);
  or (_08542_, _08541_, _04018_);
  or (_08543_, _08124_, _04792_);
  and (_08544_, _08543_, _08121_);
  and (_08545_, _08544_, _08542_);
  or (_08546_, _08545_, _08123_);
  and (_08547_, _03736_, _03387_);
  not (_08548_, _08547_);
  and (_08549_, _08548_, _08546_);
  and (_08550_, _08547_, _08525_);
  or (_08551_, _08550_, _08549_);
  and (_08552_, _08551_, _04026_);
  and (_08553_, _03919_, _03387_);
  and (_08554_, _06555_, _04025_);
  or (_08555_, _08554_, _08553_);
  or (_08556_, _08555_, _08552_);
  not (_08557_, _08553_);
  or (_08558_, _08557_, _08536_);
  and (_08559_, _08558_, _03909_);
  and (_08560_, _08559_, _08556_);
  or (_08561_, _08495_, _06556_);
  nor (_08562_, _08561_, _03909_);
  and (_08563_, _03724_, _03392_);
  or (_08564_, _08563_, _08562_);
  or (_08565_, _08564_, _08560_);
  nand (_08566_, _08563_, _08000_);
  nand (_08567_, _03729_, _03392_);
  and (_08568_, _03719_, _03392_);
  not (_08569_, _08568_);
  and (_08570_, _08569_, _08567_);
  and (_08571_, _08570_, _08566_);
  and (_08572_, _08571_, _08565_);
  and (_08573_, _03736_, _03392_);
  nor (_08574_, _08570_, _08000_);
  or (_08575_, _08574_, _08573_);
  or (_08576_, _08575_, _08572_);
  nand (_08577_, _08573_, _08524_);
  and (_08578_, _08577_, _04014_);
  and (_08579_, _08578_, _08576_);
  and (_08580_, _03919_, _03392_);
  nor (_08581_, _08580_, _04013_);
  not (_08582_, _08581_);
  not (_08583_, _08580_);
  nand (_08584_, _08583_, _06556_);
  and (_08585_, _08584_, _08582_);
  or (_08586_, _08585_, _08579_);
  nand (_08587_, _08580_, _08535_);
  and (_08588_, _08587_, _06567_);
  and (_08589_, _08588_, _08586_);
  not (_08590_, _08119_);
  nor (_08591_, _06547_, _08479_);
  nor (_08592_, _08591_, _08124_);
  nor (_08593_, _08592_, _06567_);
  or (_08594_, _08593_, _08590_);
  or (_08595_, _08594_, _08589_);
  and (_08596_, _08595_, _08120_);
  and (_08597_, _03736_, _03382_);
  or (_08598_, _08597_, _08596_);
  not (_08599_, _08597_);
  and (_08600_, _08259_, \oc8051_golden_model_1.ACC [6]);
  and (_08601_, _08264_, \oc8051_golden_model_1.ACC [5]);
  and (_08602_, _08270_, \oc8051_golden_model_1.ACC [4]);
  and (_08603_, _08282_, \oc8051_golden_model_1.ACC [3]);
  and (_08604_, _08287_, \oc8051_golden_model_1.ACC [2]);
  and (_08605_, _08294_, \oc8051_golden_model_1.ACC [1]);
  nor (_08606_, _08295_, _08296_);
  and (_08607_, _08299_, \oc8051_golden_model_1.ACC [0]);
  not (_08608_, _08607_);
  nor (_08609_, _08608_, _08606_);
  nor (_08610_, _08609_, _08605_);
  nor (_08611_, _08610_, _08290_);
  nor (_08612_, _08611_, _08604_);
  nor (_08613_, _08612_, _08285_);
  or (_08614_, _08613_, _08603_);
  and (_08615_, _08614_, _08277_);
  nor (_08616_, _08615_, _08602_);
  nor (_08617_, _08616_, _08274_);
  or (_08618_, _08617_, _08601_);
  and (_08619_, _08618_, _08311_);
  nor (_08620_, _08619_, _08600_);
  nor (_08621_, _08620_, _08255_);
  and (_08622_, _08620_, _08255_);
  nor (_08623_, _08622_, _08621_);
  or (_08624_, _08623_, _08599_);
  and (_08625_, _08624_, _04023_);
  and (_08626_, _08625_, _08598_);
  and (_08627_, _03919_, _03382_);
  nor (_08628_, _08627_, _04022_);
  not (_08629_, _08628_);
  and (_08630_, _08333_, \oc8051_golden_model_1.ACC [6]);
  and (_08631_, _08340_, \oc8051_golden_model_1.ACC [5]);
  and (_08632_, _08344_, \oc8051_golden_model_1.ACC [4]);
  and (_08633_, _08355_, \oc8051_golden_model_1.ACC [3]);
  and (_08634_, _08361_, \oc8051_golden_model_1.ACC [2]);
  and (_08635_, _08369_, \oc8051_golden_model_1.ACC [1]);
  nor (_08636_, _08370_, _08371_);
  and (_08637_, _08373_, \oc8051_golden_model_1.ACC [0]);
  not (_08638_, _08637_);
  nor (_08639_, _08638_, _08636_);
  nor (_08640_, _08639_, _08635_);
  nor (_08641_, _08640_, _08364_);
  nor (_08642_, _08641_, _08634_);
  nor (_08643_, _08642_, _08358_);
  or (_08644_, _08643_, _08633_);
  and (_08645_, _08644_, _08351_);
  nor (_08646_, _08645_, _08632_);
  nor (_08647_, _08646_, _08348_);
  or (_08648_, _08647_, _08631_);
  and (_08649_, _08648_, _08385_);
  nor (_08650_, _08649_, _08630_);
  nor (_08651_, _08650_, _08330_);
  and (_08652_, _08650_, _08330_);
  nor (_08653_, _08652_, _08651_);
  or (_08654_, _08653_, _08627_);
  and (_08655_, _08654_, _08629_);
  or (_08656_, _08655_, _08626_);
  and (_08657_, _03423_, _03382_);
  not (_08658_, _08657_);
  not (_08659_, _08627_);
  and (_08660_, _08408_, \oc8051_golden_model_1.ACC [6]);
  and (_08661_, _08413_, \oc8051_golden_model_1.ACC [5]);
  and (_08662_, _08419_, \oc8051_golden_model_1.ACC [4]);
  and (_08663_, _08425_, \oc8051_golden_model_1.ACC [3]);
  and (_08664_, _08430_, \oc8051_golden_model_1.ACC [2]);
  and (_08665_, _08437_, \oc8051_golden_model_1.ACC [1]);
  nor (_08666_, _08439_, _08438_);
  and (_08667_, _08441_, \oc8051_golden_model_1.ACC [0]);
  not (_08668_, _08667_);
  nor (_08669_, _08668_, _08666_);
  nor (_08670_, _08669_, _08665_);
  nor (_08671_, _08670_, _08433_);
  nor (_08672_, _08671_, _08664_);
  nor (_08673_, _08672_, _08428_);
  or (_08674_, _08673_, _08663_);
  and (_08675_, _08674_, _08422_);
  nor (_08676_, _08675_, _08662_);
  nor (_08677_, _08676_, _08416_);
  nor (_08678_, _08677_, _08661_);
  nor (_08679_, _08678_, _08411_);
  nor (_08680_, _08679_, _08660_);
  nor (_08681_, _08680_, _08405_);
  and (_08682_, _08680_, _08405_);
  nor (_08683_, _08682_, _08681_);
  or (_08684_, _08683_, _08659_);
  and (_08685_, _08684_, _08658_);
  and (_08686_, _08685_, _08656_);
  nand (_08687_, _08657_, \oc8051_golden_model_1.ACC [6]);
  nand (_08688_, _08687_, _07998_);
  or (_08689_, _08688_, _08686_);
  and (_08690_, _08689_, _08039_);
  and (_08691_, _03736_, _03409_);
  and (_08692_, _08037_, _07992_);
  or (_08693_, _08692_, _08691_);
  or (_08694_, _08693_, _08690_);
  and (_08695_, _06641_, \oc8051_golden_model_1.ACC [6]);
  nor (_08696_, _06641_, \oc8051_golden_model_1.ACC [6]);
  nor (_08697_, _08696_, _08695_);
  and (_08698_, _06968_, \oc8051_golden_model_1.ACC [5]);
  and (_08699_, _06873_, _07084_);
  nor (_08700_, _08699_, _08698_);
  not (_08701_, _08700_);
  and (_08702_, _06969_, \oc8051_golden_model_1.ACC [4]);
  and (_08703_, _06918_, _07090_);
  nor (_08704_, _08703_, _08702_);
  and (_08705_, _06964_, \oc8051_golden_model_1.ACC [3]);
  and (_08706_, _06779_, _07184_);
  and (_08707_, _06965_, \oc8051_golden_model_1.ACC [2]);
  and (_08708_, _06824_, _07190_);
  nor (_08709_, _08708_, _08707_);
  not (_08710_, _08709_);
  and (_08711_, _06961_, \oc8051_golden_model_1.ACC [1]);
  and (_08712_, _06688_, _03474_);
  nor (_08713_, _08712_, _08711_);
  and (_08714_, _06962_, \oc8051_golden_model_1.ACC [0]);
  and (_08715_, _08714_, _08713_);
  nor (_08716_, _08715_, _08711_);
  nor (_08717_, _08716_, _08710_);
  nor (_08718_, _08717_, _08707_);
  nor (_08719_, _08718_, _08706_);
  or (_08720_, _08719_, _08705_);
  and (_08721_, _08720_, _08704_);
  nor (_08722_, _08721_, _08702_);
  nor (_08723_, _08722_, _08701_);
  or (_08724_, _08723_, _08698_);
  and (_08725_, _08724_, _08697_);
  nor (_08726_, _08725_, _08695_);
  nor (_08727_, _08726_, _08526_);
  and (_08728_, _08726_, _08526_);
  nor (_08729_, _08728_, _08727_);
  nand (_08730_, _08729_, _08691_);
  and (_08731_, _08730_, _04140_);
  and (_08732_, _08731_, _08694_);
  and (_08733_, _03919_, _03409_);
  nor (_08734_, _06068_, _07036_);
  and (_08735_, _06068_, _07036_);
  nor (_08736_, _08735_, _08734_);
  nor (_08737_, _05859_, _07084_);
  and (_08738_, _05859_, _07084_);
  nor (_08739_, _05953_, _07090_);
  and (_08740_, _05953_, _07090_);
  nor (_08741_, _08740_, _08739_);
  and (_08742_, _05621_, _07184_);
  not (_08743_, _08742_);
  nor (_08744_, _05621_, _07184_);
  not (_08745_, _08744_);
  nor (_08746_, _05764_, _07190_);
  and (_08747_, _05764_, _07190_);
  nor (_08748_, _08747_, _08746_);
  not (_08749_, _08748_);
  nor (_08750_, _05669_, _03474_);
  and (_08751_, _05669_, _03474_);
  nor (_08752_, _08751_, _08750_);
  nor (_08753_, _05716_, _03498_);
  and (_08754_, _08753_, _08752_);
  nor (_08755_, _08754_, _08750_);
  nor (_08756_, _08755_, _08749_);
  nor (_08757_, _08756_, _08746_);
  nand (_08758_, _08757_, _08745_);
  and (_08759_, _08758_, _08743_);
  and (_08760_, _08759_, _08741_);
  nor (_08761_, _08760_, _08739_);
  nor (_08762_, _08761_, _08738_);
  or (_08763_, _08762_, _08737_);
  and (_08764_, _08763_, _08736_);
  nor (_08765_, _08764_, _08734_);
  nor (_08766_, _08765_, _06557_);
  and (_08767_, _08765_, _06557_);
  or (_08768_, _08767_, _08766_);
  and (_08769_, _08768_, _03779_);
  or (_08770_, _08769_, _08733_);
  or (_08771_, _08770_, _08732_);
  and (_08772_, _03423_, _03409_);
  not (_08773_, _08772_);
  nor (_08774_, _03810_, _07036_);
  and (_08775_, _03810_, _07036_);
  nor (_08776_, _08774_, _08775_);
  nor (_08777_, _04093_, _07084_);
  and (_08778_, _04093_, _07084_);
  nor (_08779_, _08777_, _08778_);
  not (_08780_, _08779_);
  nor (_08781_, _04526_, _07090_);
  and (_08782_, _04526_, _07090_);
  nor (_08783_, _08781_, _08782_);
  nor (_08784_, _03678_, _07184_);
  and (_08785_, _03678_, _07184_);
  nor (_08786_, _04139_, _07190_);
  and (_08787_, _04139_, _07190_);
  nor (_08788_, _08786_, _08787_);
  not (_08789_, _08788_);
  nor (_08790_, _04563_, _03474_);
  and (_08791_, _04563_, _03474_);
  nor (_08792_, _08790_, _08791_);
  nor (_08793_, _03715_, _03498_);
  and (_08794_, _08793_, _08792_);
  nor (_08795_, _08794_, _08790_);
  nor (_08796_, _08795_, _08789_);
  nor (_08797_, _08796_, _08786_);
  nor (_08798_, _08797_, _08785_);
  or (_08799_, _08798_, _08784_);
  and (_08800_, _08799_, _08783_);
  nor (_08801_, _08800_, _08781_);
  nor (_08802_, _08801_, _08780_);
  or (_08803_, _08802_, _08777_);
  and (_08804_, _08803_, _08776_);
  nor (_08805_, _08804_, _08774_);
  nor (_08806_, _08805_, _08537_);
  and (_08807_, _08805_, _08537_);
  nor (_08808_, _08807_, _08806_);
  nand (_08809_, _08808_, _08733_);
  and (_08810_, _08809_, _08773_);
  and (_08811_, _08810_, _08771_);
  and (_08812_, _08772_, \oc8051_golden_model_1.ACC [6]);
  or (_08813_, _08812_, _03773_);
  or (_08814_, _08813_, _08811_);
  and (_08815_, _03919_, _03244_);
  not (_08816_, _08815_);
  nand (_08817_, _08181_, _03773_);
  and (_08818_, _08817_, _08816_);
  and (_08819_, _08818_, _08814_);
  and (_08820_, _03423_, _03244_);
  nor (_08821_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08822_, _08821_, _07133_);
  and (_08823_, _08822_, _07053_);
  and (_08824_, _08823_, _07036_);
  nor (_08825_, _08824_, _06554_);
  and (_08826_, _08824_, _06554_);
  nor (_08827_, _08826_, _08825_);
  nor (_08828_, _08827_, _08816_);
  or (_08829_, _08828_, _08820_);
  or (_08830_, _08829_, _08819_);
  nand (_08831_, _08820_, _08297_);
  and (_08832_, _08831_, _03375_);
  and (_08833_, _08832_, _08830_);
  nor (_08834_, _08232_, _03375_);
  or (_08835_, _08834_, _03772_);
  or (_08836_, _08835_, _08833_);
  and (_08837_, _03919_, _03412_);
  not (_08838_, _08837_);
  and (_08839_, _06077_, _05429_);
  nor (_08840_, _08839_, _08124_);
  nand (_08841_, _08840_, _03772_);
  and (_08842_, _08841_, _08838_);
  and (_08843_, _08842_, _08836_);
  and (_08844_, _03423_, _03412_);
  and (_08845_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08846_, _08845_, _07134_);
  nor (_08847_, _08846_, _07090_);
  and (_08848_, _08847_, \oc8051_golden_model_1.ACC [5]);
  and (_08849_, _08848_, \oc8051_golden_model_1.ACC [6]);
  nor (_08850_, _08849_, \oc8051_golden_model_1.ACC [7]);
  and (_08851_, _08849_, \oc8051_golden_model_1.ACC [7]);
  nor (_08852_, _08851_, _08850_);
  and (_08853_, _08852_, _08837_);
  or (_08854_, _08853_, _08844_);
  or (_08855_, _08854_, _08843_);
  nand (_08856_, _08844_, _03498_);
  and (_08857_, _08856_, _43152_);
  and (_08858_, _08857_, _08855_);
  or (_08859_, _08858_, _07991_);
  and (_40681_, _08859_, _41894_);
  not (_08860_, \oc8051_golden_model_1.SBUF [7]);
  nor (_08861_, _05491_, _08860_);
  and (_08862_, _06077_, _05491_);
  nor (_08863_, _08862_, _08861_);
  nor (_08864_, _08863_, _04060_);
  and (_08865_, _06557_, _05491_);
  nor (_08866_, _08865_, _08861_);
  nor (_08867_, _08866_, _04792_);
  and (_08868_, _05491_, \oc8051_golden_model_1.ACC [7]);
  nor (_08869_, _08868_, _08861_);
  nor (_08870_, _08869_, _04708_);
  nor (_08871_, _04707_, _08860_);
  or (_08872_, _08871_, _08870_);
  and (_08873_, _08872_, _04722_);
  and (_08874_, _06160_, _05491_);
  nor (_08875_, _08874_, _08861_);
  nor (_08876_, _08875_, _04722_);
  or (_08877_, _08876_, _08873_);
  and (_08878_, _08877_, _04733_);
  and (_08879_, _05568_, _05491_);
  nor (_08880_, _08879_, _08861_);
  nor (_08881_, _08880_, _04733_);
  nor (_08882_, _08881_, _08878_);
  nor (_08883_, _08882_, _03854_);
  nor (_08884_, _08869_, _03855_);
  or (_08886_, _08884_, _07927_);
  or (_08887_, _08886_, _08883_);
  and (_08888_, _06248_, _05491_);
  nor (_08889_, _08861_, _03738_);
  not (_08890_, _08889_);
  nor (_08891_, _08890_, _08888_);
  and (_08892_, _08880_, _08474_);
  or (_08893_, _08892_, _03455_);
  nor (_08894_, _08893_, _08891_);
  and (_08895_, _08894_, _08887_);
  not (_08897_, _05491_);
  nor (_08898_, _06536_, _08897_);
  nor (_08899_, _08898_, _08861_);
  nor (_08900_, _08899_, _03820_);
  or (_08901_, _08900_, _08895_);
  and (_08902_, _08901_, _04778_);
  and (_08903_, _06348_, _05491_);
  nor (_08904_, _08903_, _08861_);
  nor (_08905_, _08904_, _04778_);
  or (_08906_, _08905_, _08902_);
  and (_08908_, _08906_, _04790_);
  and (_08909_, _06549_, _05491_);
  nor (_08910_, _08909_, _08861_);
  nor (_08911_, _08910_, _04790_);
  or (_08912_, _08911_, _08908_);
  and (_08913_, _08912_, _04792_);
  nor (_08914_, _08913_, _08867_);
  nor (_08915_, _08914_, _03908_);
  nor (_08916_, _08861_, _05571_);
  not (_08917_, _08916_);
  nor (_08919_, _08904_, _03909_);
  and (_08920_, _08919_, _08917_);
  nor (_08921_, _08920_, _08915_);
  nor (_08922_, _08921_, _04027_);
  nor (_08923_, _08869_, _04785_);
  and (_08924_, _08923_, _08917_);
  or (_08925_, _08924_, _08922_);
  and (_08926_, _08925_, _06567_);
  nor (_08927_, _06547_, _08897_);
  nor (_08928_, _08927_, _08861_);
  nor (_08930_, _08928_, _06567_);
  or (_08931_, _08930_, _08926_);
  and (_08932_, _08931_, _06572_);
  nor (_08933_, _06556_, _08897_);
  nor (_08934_, _08933_, _08861_);
  nor (_08935_, _08934_, _06572_);
  or (_08936_, _08935_, _08932_);
  and (_08937_, _08936_, _03774_);
  nor (_08938_, _08875_, _03774_);
  or (_08939_, _08938_, _08937_);
  and (_08941_, _08939_, _04060_);
  nor (_08942_, _08941_, _08864_);
  nand (_08943_, _08942_, _43152_);
  or (_08944_, _43152_, \oc8051_golden_model_1.SBUF [7]);
  and (_08945_, _08944_, _41894_);
  and (_40683_, _08945_, _08943_);
  not (_08946_, \oc8051_golden_model_1.SCON [7]);
  nor (_08947_, _05465_, _08946_);
  and (_08948_, _06557_, _05465_);
  nor (_08949_, _08948_, _08947_);
  nor (_08951_, _08949_, _04792_);
  and (_08952_, _05465_, \oc8051_golden_model_1.ACC [7]);
  nor (_08953_, _08952_, _08947_);
  nor (_08954_, _08953_, _04708_);
  nor (_08955_, _04707_, _08946_);
  or (_08956_, _08955_, _08954_);
  and (_08957_, _08956_, _04722_);
  and (_08958_, _06160_, _05465_);
  nor (_08959_, _08958_, _08947_);
  nor (_08960_, _08959_, _04722_);
  or (_08961_, _08960_, _08957_);
  and (_08962_, _08961_, _03764_);
  nor (_08963_, _06101_, _08946_);
  and (_08964_, _06148_, _06101_);
  nor (_08965_, _08964_, _08963_);
  nor (_08966_, _08965_, _03764_);
  or (_08967_, _08966_, _03848_);
  or (_08968_, _08967_, _08962_);
  and (_08969_, _05568_, _05465_);
  nor (_08970_, _08969_, _08947_);
  nand (_08971_, _08970_, _03848_);
  and (_08972_, _08971_, _08968_);
  and (_08973_, _08972_, _03855_);
  nor (_08974_, _08953_, _03855_);
  or (_08975_, _08974_, _08973_);
  and (_08976_, _08975_, _03760_);
  and (_08977_, _06121_, _06101_);
  nor (_08978_, _08977_, _08963_);
  nor (_08979_, _08978_, _03760_);
  or (_08980_, _08979_, _03752_);
  or (_08981_, _08980_, _08976_);
  nor (_08982_, _08963_, _06147_);
  nor (_08983_, _08982_, _08965_);
  or (_08984_, _08983_, _03753_);
  and (_08985_, _08984_, _03747_);
  and (_08986_, _08985_, _08981_);
  not (_08987_, _06101_);
  nor (_08988_, _06143_, _08987_);
  nor (_08989_, _08988_, _08963_);
  nor (_08990_, _08989_, _03747_);
  or (_08991_, _08990_, _07927_);
  or (_08992_, _08991_, _08986_);
  and (_08993_, _06248_, _05465_);
  nor (_08994_, _08947_, _03738_);
  not (_08995_, _08994_);
  nor (_08996_, _08995_, _08993_);
  and (_08997_, _08970_, _08474_);
  or (_08998_, _08997_, _03455_);
  nor (_08999_, _08998_, _08996_);
  and (_09000_, _08999_, _08992_);
  not (_09001_, _05465_);
  nor (_09002_, _06536_, _09001_);
  nor (_09003_, _09002_, _08947_);
  nor (_09004_, _09003_, _03820_);
  or (_09005_, _09004_, _09000_);
  and (_09006_, _09005_, _04778_);
  and (_09007_, _06348_, _05465_);
  nor (_09008_, _09007_, _08947_);
  nor (_09009_, _09008_, _04778_);
  or (_09010_, _09009_, _09006_);
  nor (_09011_, _09010_, _03897_);
  and (_09012_, _06549_, _05465_);
  or (_09013_, _08947_, _04790_);
  nor (_09014_, _09013_, _09012_);
  or (_09015_, _09014_, _04018_);
  nor (_09016_, _09015_, _09011_);
  nor (_09017_, _09016_, _08951_);
  nor (_09018_, _09017_, _03908_);
  nor (_09019_, _08947_, _05571_);
  not (_09020_, _09019_);
  nor (_09021_, _09008_, _03909_);
  and (_09022_, _09021_, _09020_);
  nor (_09023_, _09022_, _09018_);
  nor (_09024_, _09023_, _04027_);
  nor (_09025_, _08953_, _04785_);
  and (_09026_, _09025_, _09020_);
  or (_09027_, _09026_, _09024_);
  and (_09028_, _09027_, _06567_);
  nor (_09029_, _06547_, _09001_);
  nor (_09030_, _09029_, _08947_);
  nor (_09031_, _09030_, _06567_);
  or (_09032_, _09031_, _09028_);
  and (_09033_, _09032_, _06572_);
  nor (_09034_, _06556_, _09001_);
  nor (_09035_, _09034_, _08947_);
  nor (_09036_, _09035_, _06572_);
  or (_09037_, _09036_, _09033_);
  and (_09038_, _09037_, _03774_);
  nor (_09039_, _08959_, _03774_);
  or (_09040_, _09039_, _09038_);
  and (_09041_, _09040_, _03375_);
  nor (_09042_, _08978_, _03375_);
  or (_09043_, _09042_, _09041_);
  and (_09044_, _09043_, _04060_);
  and (_09045_, _06077_, _05465_);
  nor (_09046_, _09045_, _08947_);
  nor (_09047_, _09046_, _04060_);
  or (_09048_, _09047_, _09044_);
  or (_09049_, _09048_, _43156_);
  or (_09050_, _43152_, \oc8051_golden_model_1.SCON [7]);
  and (_09051_, _09050_, _41894_);
  and (_40684_, _09051_, _09049_);
  not (_09052_, \oc8051_golden_model_1.PCON [7]);
  nor (_09053_, _05488_, _09052_);
  and (_09054_, _06077_, _05488_);
  nor (_09055_, _09054_, _09053_);
  nor (_09056_, _09055_, _04060_);
  and (_09057_, _06557_, _05488_);
  nor (_09058_, _09057_, _09053_);
  nor (_09059_, _09058_, _04792_);
  and (_09060_, _05488_, \oc8051_golden_model_1.ACC [7]);
  nor (_09061_, _09060_, _09053_);
  nor (_09062_, _09061_, _04708_);
  nor (_09063_, _04707_, _09052_);
  or (_09064_, _09063_, _09062_);
  and (_09065_, _09064_, _04722_);
  and (_09066_, _06160_, _05488_);
  nor (_09067_, _09066_, _09053_);
  nor (_09068_, _09067_, _04722_);
  or (_09069_, _09068_, _09065_);
  and (_09070_, _09069_, _04733_);
  and (_09071_, _05568_, _05488_);
  nor (_09072_, _09071_, _09053_);
  nor (_09073_, _09072_, _04733_);
  nor (_09074_, _09073_, _09070_);
  nor (_09075_, _09074_, _03854_);
  nor (_09076_, _09061_, _03855_);
  or (_09077_, _09076_, _07927_);
  or (_09078_, _09077_, _09075_);
  and (_09079_, _06248_, _05488_);
  nor (_09080_, _09053_, _03738_);
  not (_09081_, _09080_);
  nor (_09082_, _09081_, _09079_);
  and (_09083_, _09072_, _08474_);
  or (_09084_, _09083_, _03455_);
  nor (_09085_, _09084_, _09082_);
  and (_09086_, _09085_, _09078_);
  not (_09087_, _05488_);
  nor (_09088_, _06536_, _09087_);
  nor (_09089_, _09088_, _09053_);
  nor (_09090_, _09089_, _03820_);
  or (_09091_, _09090_, _09086_);
  and (_09092_, _09091_, _04778_);
  and (_09093_, _06348_, _05488_);
  nor (_09094_, _09093_, _09053_);
  nor (_09095_, _09094_, _04778_);
  or (_09096_, _09095_, _09092_);
  and (_09097_, _09096_, _04790_);
  and (_09098_, _06549_, _05488_);
  nor (_09099_, _09098_, _09053_);
  nor (_09100_, _09099_, _04790_);
  or (_09101_, _09100_, _09097_);
  and (_09102_, _09101_, _04792_);
  nor (_09103_, _09102_, _09059_);
  nor (_09104_, _09103_, _03908_);
  nor (_09105_, _09053_, _05571_);
  not (_09106_, _09105_);
  nor (_09107_, _09094_, _03909_);
  and (_09108_, _09107_, _09106_);
  nor (_09109_, _09108_, _09104_);
  nor (_09110_, _09109_, _04027_);
  nor (_09111_, _09061_, _04785_);
  and (_09112_, _09111_, _09106_);
  or (_09113_, _09112_, _09110_);
  and (_09114_, _09113_, _06567_);
  nor (_09115_, _06547_, _09087_);
  nor (_09116_, _09115_, _09053_);
  nor (_09117_, _09116_, _06567_);
  or (_09118_, _09117_, _09114_);
  and (_09119_, _09118_, _06572_);
  nor (_09120_, _06556_, _09087_);
  nor (_09121_, _09120_, _09053_);
  nor (_09122_, _09121_, _06572_);
  or (_09123_, _09122_, _09119_);
  and (_09124_, _09123_, _03774_);
  nor (_09125_, _09067_, _03774_);
  or (_09126_, _09125_, _09124_);
  and (_09127_, _09126_, _04060_);
  nor (_09128_, _09127_, _09056_);
  nand (_09129_, _09128_, _43152_);
  or (_09130_, _43152_, \oc8051_golden_model_1.PCON [7]);
  and (_09131_, _09130_, _41894_);
  and (_40685_, _09131_, _09129_);
  not (_09132_, \oc8051_golden_model_1.TCON [7]);
  nor (_09133_, _05447_, _09132_);
  and (_09134_, _06557_, _05447_);
  nor (_09135_, _09134_, _09133_);
  nor (_09136_, _09135_, _04792_);
  and (_09137_, _05447_, \oc8051_golden_model_1.ACC [7]);
  nor (_09138_, _09137_, _09133_);
  nor (_09139_, _09138_, _04708_);
  nor (_09140_, _04707_, _09132_);
  or (_09141_, _09140_, _09139_);
  and (_09142_, _09141_, _04722_);
  and (_09143_, _06160_, _05447_);
  nor (_09144_, _09143_, _09133_);
  nor (_09145_, _09144_, _04722_);
  or (_09146_, _09145_, _09142_);
  and (_09147_, _09146_, _03764_);
  nor (_09148_, _06085_, _09132_);
  and (_09149_, _06148_, _06085_);
  nor (_09150_, _09149_, _09148_);
  nor (_09151_, _09150_, _03764_);
  or (_09152_, _09151_, _03848_);
  or (_09153_, _09152_, _09147_);
  and (_09154_, _05568_, _05447_);
  nor (_09155_, _09154_, _09133_);
  nand (_09156_, _09155_, _03848_);
  and (_09157_, _09156_, _09153_);
  and (_09158_, _09157_, _03855_);
  nor (_09159_, _09138_, _03855_);
  or (_09160_, _09159_, _09158_);
  and (_09161_, _09160_, _03760_);
  and (_09162_, _06121_, _06085_);
  nor (_09163_, _09162_, _09148_);
  nor (_09164_, _09163_, _03760_);
  or (_09165_, _09164_, _09161_);
  and (_09166_, _09165_, _03753_);
  nor (_09167_, _09148_, _06147_);
  nor (_09168_, _09167_, _09150_);
  and (_09169_, _09168_, _03752_);
  or (_09170_, _09169_, _09166_);
  and (_09171_, _09170_, _03747_);
  not (_09172_, _06085_);
  nor (_09173_, _06143_, _09172_);
  nor (_09174_, _09173_, _09148_);
  nor (_09175_, _09174_, _03747_);
  or (_09176_, _09175_, _07927_);
  or (_09177_, _09176_, _09171_);
  and (_09178_, _06248_, _05447_);
  nor (_09179_, _09133_, _03738_);
  not (_09180_, _09179_);
  nor (_09181_, _09180_, _09178_);
  and (_09182_, _09155_, _08474_);
  or (_09183_, _09182_, _03455_);
  nor (_09184_, _09183_, _09181_);
  and (_09185_, _09184_, _09177_);
  not (_09186_, _05447_);
  nor (_09187_, _06536_, _09186_);
  nor (_09188_, _09187_, _09133_);
  nor (_09189_, _09188_, _03820_);
  or (_09190_, _09189_, _09185_);
  and (_09191_, _09190_, _04778_);
  and (_09192_, _06348_, _05447_);
  nor (_09193_, _09192_, _09133_);
  nor (_09194_, _09193_, _04778_);
  or (_09195_, _09194_, _09191_);
  and (_09196_, _09195_, _04790_);
  and (_09197_, _06549_, _05447_);
  nor (_09198_, _09197_, _09133_);
  nor (_09199_, _09198_, _04790_);
  or (_09200_, _09199_, _09196_);
  and (_09201_, _09200_, _04792_);
  nor (_09202_, _09201_, _09136_);
  nor (_09203_, _09202_, _03908_);
  nor (_09204_, _09133_, _05571_);
  not (_09205_, _09204_);
  nor (_09206_, _09193_, _03909_);
  and (_09207_, _09206_, _09205_);
  nor (_09208_, _09207_, _09203_);
  nor (_09209_, _09208_, _04027_);
  nor (_09210_, _09138_, _04785_);
  and (_09211_, _09210_, _09205_);
  or (_09212_, _09211_, _09209_);
  and (_09213_, _09212_, _06567_);
  nor (_09214_, _06547_, _09186_);
  nor (_09215_, _09214_, _09133_);
  nor (_09216_, _09215_, _06567_);
  or (_09217_, _09216_, _09213_);
  and (_09218_, _09217_, _06572_);
  nor (_09219_, _06556_, _09186_);
  nor (_09220_, _09219_, _09133_);
  nor (_09221_, _09220_, _06572_);
  or (_09222_, _09221_, _09218_);
  and (_09223_, _09222_, _03774_);
  nor (_09224_, _09144_, _03774_);
  or (_09225_, _09224_, _09223_);
  and (_09226_, _09225_, _03375_);
  nor (_09227_, _09163_, _03375_);
  or (_09228_, _09227_, _09226_);
  and (_09229_, _09228_, _04060_);
  and (_09230_, _06077_, _05447_);
  nor (_09231_, _09230_, _09133_);
  nor (_09232_, _09231_, _04060_);
  or (_09233_, _09232_, _09229_);
  or (_09234_, _09233_, _43156_);
  or (_09235_, _43152_, \oc8051_golden_model_1.TCON [7]);
  and (_09236_, _09235_, _41894_);
  and (_40686_, _09236_, _09234_);
  not (_09237_, \oc8051_golden_model_1.TL0 [7]);
  nor (_09238_, _05589_, _09237_);
  and (_09239_, _06077_, _05589_);
  nor (_09240_, _09239_, _09238_);
  nor (_09241_, _09240_, _04060_);
  and (_09242_, _06557_, _05589_);
  nor (_09243_, _09242_, _09238_);
  nor (_09244_, _09243_, _04792_);
  and (_09245_, _05589_, \oc8051_golden_model_1.ACC [7]);
  nor (_09246_, _09245_, _09238_);
  nor (_09247_, _09246_, _04708_);
  nor (_09248_, _04707_, _09237_);
  or (_09249_, _09248_, _09247_);
  and (_09250_, _09249_, _04722_);
  and (_09251_, _06160_, _05589_);
  nor (_09252_, _09251_, _09238_);
  nor (_09253_, _09252_, _04722_);
  or (_09254_, _09253_, _09250_);
  and (_09255_, _09254_, _04733_);
  and (_09256_, _05568_, _05589_);
  nor (_09257_, _09256_, _09238_);
  nor (_09258_, _09257_, _04733_);
  nor (_09259_, _09258_, _09255_);
  nor (_09260_, _09259_, _03854_);
  nor (_09261_, _09246_, _03855_);
  or (_09262_, _09261_, _07927_);
  nor (_09263_, _09262_, _09260_);
  nor (_09264_, _09238_, _03738_);
  nand (_09265_, _06248_, _05589_);
  and (_09266_, _09265_, _09264_);
  and (_09267_, _09257_, _08474_);
  or (_09268_, _09267_, _03455_);
  or (_09269_, _09268_, _09266_);
  nor (_09270_, _09269_, _09263_);
  not (_09271_, _05589_);
  nor (_09272_, _06536_, _09271_);
  nor (_09273_, _09272_, _09238_);
  nor (_09274_, _09273_, _03820_);
  or (_09275_, _09274_, _09270_);
  and (_09276_, _09275_, _04778_);
  and (_09277_, _06348_, _05589_);
  nor (_09278_, _09277_, _09238_);
  nor (_09279_, _09278_, _04778_);
  or (_09280_, _09279_, _09276_);
  and (_09281_, _09280_, _04790_);
  and (_09282_, _06549_, _05480_);
  nor (_09283_, _09282_, _09238_);
  nor (_09284_, _09283_, _04790_);
  or (_09285_, _09284_, _09281_);
  and (_09286_, _09285_, _04792_);
  nor (_09287_, _09286_, _09244_);
  nor (_09288_, _09287_, _03908_);
  nor (_09289_, _09238_, _05571_);
  not (_09290_, _09289_);
  nor (_09291_, _09278_, _03909_);
  and (_09292_, _09291_, _09290_);
  nor (_09293_, _09292_, _09288_);
  nor (_09294_, _09293_, _04027_);
  nor (_09295_, _09246_, _04785_);
  and (_09296_, _09295_, _09290_);
  nor (_09297_, _09296_, _03914_);
  not (_09298_, _09297_);
  nor (_09299_, _09298_, _09294_);
  or (_09300_, _06547_, _09271_);
  nor (_09301_, _09238_, _06567_);
  and (_09302_, _09301_, _09300_);
  or (_09303_, _09302_, _04011_);
  nor (_09304_, _09303_, _09299_);
  nor (_09305_, _06556_, _09271_);
  nor (_09306_, _09305_, _09238_);
  nor (_09307_, _09306_, _06572_);
  or (_09308_, _09307_, _09304_);
  and (_09309_, _09308_, _03774_);
  nor (_09310_, _09252_, _03774_);
  or (_09311_, _09310_, _09309_);
  and (_09312_, _09311_, _04060_);
  nor (_09313_, _09312_, _09241_);
  nand (_09314_, _09313_, _43152_);
  or (_09315_, _43152_, \oc8051_golden_model_1.TL0 [7]);
  and (_09316_, _09315_, _41894_);
  and (_40687_, _09316_, _09314_);
  not (_09317_, \oc8051_golden_model_1.TL1 [7]);
  nor (_09318_, _05587_, _09317_);
  and (_09319_, _06077_, _05587_);
  nor (_09320_, _09319_, _09318_);
  nor (_09321_, _09320_, _04060_);
  and (_09322_, _06557_, _05587_);
  nor (_09323_, _09322_, _09318_);
  nor (_09324_, _09323_, _04792_);
  and (_09325_, _05461_, \oc8051_golden_model_1.ACC [7]);
  nor (_09326_, _09325_, _09318_);
  nor (_09327_, _09326_, _04708_);
  nor (_09328_, _04707_, _09317_);
  or (_09329_, _09328_, _09327_);
  and (_09330_, _09329_, _04722_);
  and (_09331_, _06160_, _05587_);
  nor (_09332_, _09331_, _09318_);
  nor (_09333_, _09332_, _04722_);
  or (_09334_, _09333_, _09330_);
  and (_09335_, _09334_, _04733_);
  and (_09336_, _05568_, _05587_);
  nor (_09337_, _09336_, _09318_);
  nor (_09338_, _09337_, _04733_);
  nor (_09339_, _09338_, _09335_);
  nor (_09340_, _09339_, _03854_);
  nor (_09341_, _09326_, _03855_);
  or (_09342_, _09341_, _07927_);
  or (_09343_, _09342_, _09340_);
  nor (_09344_, _09318_, _03738_);
  nand (_09345_, _06248_, _05587_);
  and (_09346_, _09345_, _09344_);
  and (_09347_, _09337_, _08474_);
  or (_09348_, _09347_, _03455_);
  nor (_09349_, _09348_, _09346_);
  and (_09350_, _09349_, _09343_);
  not (_09351_, _05587_);
  nor (_09352_, _06536_, _09351_);
  nor (_09353_, _09352_, _09318_);
  nor (_09354_, _09353_, _03820_);
  or (_09355_, _09354_, _09350_);
  and (_09356_, _09355_, _04778_);
  and (_09357_, _06348_, _05461_);
  nor (_09358_, _09357_, _09318_);
  nor (_09359_, _09358_, _04778_);
  or (_09360_, _09359_, _09356_);
  nor (_09361_, _09360_, _03897_);
  nand (_09362_, _06549_, _05587_);
  nor (_09363_, _09318_, _04790_);
  and (_09364_, _09363_, _09362_);
  or (_09365_, _09364_, _04018_);
  nor (_09366_, _09365_, _09361_);
  nor (_09367_, _09366_, _09324_);
  nor (_09368_, _09367_, _03908_);
  nor (_09369_, _09318_, _05571_);
  not (_09370_, _09369_);
  nor (_09371_, _09358_, _03909_);
  and (_09372_, _09371_, _09370_);
  nor (_09373_, _09372_, _09368_);
  nor (_09374_, _09373_, _04027_);
  nor (_09375_, _09326_, _04785_);
  and (_09376_, _09375_, _09370_);
  nor (_09377_, _09376_, _03914_);
  not (_09378_, _09377_);
  nor (_09379_, _09378_, _09374_);
  or (_09380_, _06547_, _09351_);
  nor (_09381_, _09318_, _06567_);
  and (_09382_, _09381_, _09380_);
  or (_09383_, _09382_, _04011_);
  nor (_09384_, _09383_, _09379_);
  nor (_09385_, _06556_, _09351_);
  nor (_09386_, _09385_, _09318_);
  nor (_09387_, _09386_, _06572_);
  or (_09388_, _09387_, _09384_);
  and (_09389_, _09388_, _03774_);
  nor (_09390_, _09332_, _03774_);
  or (_09391_, _09390_, _09389_);
  and (_09392_, _09391_, _04060_);
  nor (_09393_, _09392_, _09321_);
  nand (_09394_, _09393_, _43152_);
  or (_09395_, _43152_, \oc8051_golden_model_1.TL1 [7]);
  and (_09396_, _09395_, _41894_);
  and (_40689_, _09396_, _09394_);
  not (_09397_, \oc8051_golden_model_1.TH0 [7]);
  nor (_09398_, _05451_, _09397_);
  and (_09399_, _06077_, _05451_);
  nor (_09400_, _09399_, _09398_);
  nor (_09401_, _09400_, _04060_);
  and (_09402_, _06557_, _05451_);
  nor (_09403_, _09402_, _09398_);
  nor (_09404_, _09403_, _04792_);
  and (_09405_, _05451_, \oc8051_golden_model_1.ACC [7]);
  nor (_09406_, _09405_, _09398_);
  nor (_09407_, _09406_, _04708_);
  nor (_09408_, _04707_, _09397_);
  or (_09409_, _09408_, _09407_);
  and (_09410_, _09409_, _04722_);
  and (_09411_, _06160_, _05451_);
  nor (_09412_, _09411_, _09398_);
  nor (_09413_, _09412_, _04722_);
  or (_09414_, _09413_, _09410_);
  and (_09415_, _09414_, _04733_);
  and (_09416_, _05568_, _05451_);
  nor (_09417_, _09416_, _09398_);
  nor (_09418_, _09417_, _04733_);
  nor (_09419_, _09418_, _09415_);
  nor (_09420_, _09419_, _03854_);
  nor (_09421_, _09406_, _03855_);
  or (_09422_, _09421_, _07927_);
  or (_09423_, _09422_, _09420_);
  and (_09424_, _06248_, _05451_);
  nor (_09425_, _09398_, _03738_);
  not (_09426_, _09425_);
  nor (_09427_, _09426_, _09424_);
  and (_09428_, _09417_, _08474_);
  or (_09429_, _09428_, _03455_);
  nor (_09430_, _09429_, _09427_);
  and (_09431_, _09430_, _09423_);
  not (_09432_, _05451_);
  nor (_09433_, _06536_, _09432_);
  nor (_09434_, _09433_, _09398_);
  nor (_09435_, _09434_, _03820_);
  or (_09436_, _09435_, _09431_);
  and (_09437_, _09436_, _04778_);
  and (_09438_, _06348_, _05451_);
  nor (_09439_, _09438_, _09398_);
  nor (_09440_, _09439_, _04778_);
  or (_09441_, _09440_, _09437_);
  nor (_09442_, _09441_, _03897_);
  and (_09443_, _06549_, _05451_);
  or (_09444_, _09398_, _04790_);
  nor (_09445_, _09444_, _09443_);
  or (_09446_, _09445_, _04018_);
  nor (_09447_, _09446_, _09442_);
  nor (_09448_, _09447_, _09404_);
  nor (_09449_, _09448_, _03908_);
  nor (_09450_, _09398_, _05571_);
  not (_09451_, _09450_);
  nor (_09452_, _09439_, _03909_);
  and (_09453_, _09452_, _09451_);
  nor (_09454_, _09453_, _09449_);
  nor (_09455_, _09454_, _04027_);
  nor (_09456_, _09406_, _04785_);
  and (_09457_, _09456_, _09451_);
  nor (_09458_, _09457_, _03914_);
  not (_09459_, _09458_);
  nor (_09460_, _09459_, _09455_);
  nor (_09461_, _06547_, _09432_);
  or (_09462_, _09398_, _06567_);
  nor (_09463_, _09462_, _09461_);
  or (_09464_, _09463_, _04011_);
  nor (_09465_, _09464_, _09460_);
  nor (_09466_, _06556_, _09432_);
  nor (_09467_, _09466_, _09398_);
  nor (_09468_, _09467_, _06572_);
  or (_09469_, _09468_, _09465_);
  and (_09470_, _09469_, _03774_);
  nor (_09471_, _09412_, _03774_);
  or (_09472_, _09471_, _09470_);
  and (_09473_, _09472_, _04060_);
  nor (_09474_, _09473_, _09401_);
  nand (_09475_, _09474_, _43152_);
  or (_09476_, _43152_, \oc8051_golden_model_1.TH0 [7]);
  and (_09477_, _09476_, _41894_);
  and (_40690_, _09477_, _09475_);
  not (_09478_, \oc8051_golden_model_1.TH1 [7]);
  nor (_09479_, _05469_, _09478_);
  and (_09480_, _06077_, _05469_);
  nor (_09481_, _09480_, _09479_);
  nor (_09482_, _09481_, _04060_);
  and (_09483_, _06557_, _05469_);
  nor (_09484_, _09483_, _09479_);
  nor (_09485_, _09484_, _04792_);
  and (_09486_, _05469_, \oc8051_golden_model_1.ACC [7]);
  nor (_09487_, _09486_, _09479_);
  nor (_09488_, _09487_, _04708_);
  nor (_09489_, _04707_, _09478_);
  or (_09490_, _09489_, _09488_);
  and (_09491_, _09490_, _04722_);
  and (_09492_, _06160_, _05469_);
  nor (_09493_, _09492_, _09479_);
  nor (_09494_, _09493_, _04722_);
  or (_09496_, _09494_, _09491_);
  and (_09497_, _09496_, _04733_);
  and (_09498_, _05568_, _05469_);
  nor (_09499_, _09498_, _09479_);
  nor (_09500_, _09499_, _04733_);
  nor (_09501_, _09500_, _09497_);
  nor (_09502_, _09501_, _03854_);
  nor (_09503_, _09487_, _03855_);
  or (_09504_, _09503_, _07927_);
  or (_09505_, _09504_, _09502_);
  and (_09506_, _06248_, _05469_);
  nor (_09507_, _09479_, _03738_);
  not (_09508_, _09507_);
  nor (_09509_, _09508_, _09506_);
  and (_09510_, _09499_, _08474_);
  or (_09511_, _09510_, _03455_);
  nor (_09512_, _09511_, _09509_);
  and (_09513_, _09512_, _09505_);
  not (_09514_, _05469_);
  nor (_09515_, _06536_, _09514_);
  nor (_09517_, _09515_, _09479_);
  nor (_09518_, _09517_, _03820_);
  or (_09519_, _09518_, _09513_);
  and (_09520_, _09519_, _04778_);
  and (_09521_, _06348_, _05469_);
  nor (_09522_, _09521_, _09479_);
  nor (_09523_, _09522_, _04778_);
  or (_09524_, _09523_, _09520_);
  nor (_09525_, _09524_, _03897_);
  and (_09526_, _06549_, _05469_);
  or (_09527_, _09479_, _04790_);
  nor (_09528_, _09527_, _09526_);
  or (_09529_, _09528_, _04018_);
  nor (_09530_, _09529_, _09525_);
  nor (_09531_, _09530_, _09485_);
  nor (_09532_, _09531_, _03908_);
  nor (_09533_, _09479_, _05571_);
  not (_09534_, _09533_);
  nor (_09535_, _09522_, _03909_);
  and (_09536_, _09535_, _09534_);
  nor (_09537_, _09536_, _09532_);
  nor (_09538_, _09537_, _04027_);
  nor (_09539_, _09487_, _04785_);
  and (_09540_, _09539_, _09534_);
  or (_09541_, _09540_, _09538_);
  and (_09542_, _09541_, _06567_);
  nor (_09543_, _06547_, _09514_);
  nor (_09544_, _09543_, _09479_);
  nor (_09545_, _09544_, _06567_);
  or (_09546_, _09545_, _09542_);
  and (_09547_, _09546_, _06572_);
  nor (_09548_, _06556_, _09514_);
  nor (_09549_, _09548_, _09479_);
  nor (_09550_, _09549_, _06572_);
  or (_09551_, _09550_, _09547_);
  and (_09552_, _09551_, _03774_);
  nor (_09553_, _09493_, _03774_);
  or (_09554_, _09553_, _09552_);
  and (_09555_, _09554_, _04060_);
  nor (_09556_, _09555_, _09482_);
  nand (_09557_, _09556_, _43152_);
  or (_09558_, _43152_, \oc8051_golden_model_1.TH1 [7]);
  and (_09559_, _09558_, _41894_);
  and (_40691_, _09559_, _09557_);
  not (_09560_, \oc8051_golden_model_1.TMOD [7]);
  nor (_09561_, _05475_, _09560_);
  and (_09562_, _06077_, _05475_);
  nor (_09563_, _09562_, _09561_);
  nor (_09564_, _09563_, _04060_);
  and (_09565_, _06557_, _05475_);
  nor (_09566_, _09565_, _09561_);
  nor (_09567_, _09566_, _04792_);
  and (_09568_, _05475_, \oc8051_golden_model_1.ACC [7]);
  nor (_09569_, _09568_, _09561_);
  nor (_09570_, _09569_, _04708_);
  nor (_09571_, _04707_, _09560_);
  or (_09572_, _09571_, _09570_);
  and (_09573_, _09572_, _04722_);
  and (_09574_, _06160_, _05475_);
  nor (_09575_, _09574_, _09561_);
  nor (_09576_, _09575_, _04722_);
  or (_09577_, _09576_, _09573_);
  and (_09578_, _09577_, _04733_);
  and (_09579_, _05568_, _05475_);
  nor (_09580_, _09579_, _09561_);
  nor (_09581_, _09580_, _04733_);
  nor (_09582_, _09581_, _09578_);
  nor (_09583_, _09582_, _03854_);
  nor (_09584_, _09569_, _03855_);
  or (_09585_, _09584_, _07927_);
  or (_09586_, _09585_, _09583_);
  and (_09587_, _06248_, _05475_);
  nor (_09588_, _09561_, _03738_);
  not (_09589_, _09588_);
  nor (_09590_, _09589_, _09587_);
  and (_09591_, _09580_, _08474_);
  or (_09592_, _09591_, _03455_);
  nor (_09593_, _09592_, _09590_);
  and (_09594_, _09593_, _09586_);
  not (_09595_, _05475_);
  nor (_09596_, _06536_, _09595_);
  nor (_09597_, _09596_, _09561_);
  nor (_09598_, _09597_, _03820_);
  or (_09599_, _09598_, _09594_);
  and (_09600_, _09599_, _04778_);
  and (_09601_, _06348_, _05475_);
  nor (_09602_, _09601_, _09561_);
  nor (_09603_, _09602_, _04778_);
  or (_09604_, _09603_, _09600_);
  and (_09605_, _09604_, _04790_);
  and (_09606_, _06549_, _05475_);
  nor (_09607_, _09606_, _09561_);
  nor (_09608_, _09607_, _04790_);
  or (_09609_, _09608_, _09605_);
  and (_09610_, _09609_, _04792_);
  nor (_09611_, _09610_, _09567_);
  nor (_09612_, _09611_, _03908_);
  nor (_09613_, _09561_, _05571_);
  not (_09614_, _09613_);
  nor (_09615_, _09602_, _03909_);
  and (_09616_, _09615_, _09614_);
  nor (_09617_, _09616_, _09612_);
  nor (_09618_, _09617_, _04027_);
  nor (_09619_, _09569_, _04785_);
  and (_09620_, _09619_, _09614_);
  or (_09621_, _09620_, _09618_);
  and (_09622_, _09621_, _06567_);
  nor (_09623_, _06547_, _09595_);
  nor (_09624_, _09623_, _09561_);
  nor (_09625_, _09624_, _06567_);
  or (_09626_, _09625_, _09622_);
  and (_09627_, _09626_, _06572_);
  nor (_09628_, _06556_, _09595_);
  nor (_09629_, _09628_, _09561_);
  nor (_09630_, _09629_, _06572_);
  or (_09631_, _09630_, _09627_);
  and (_09632_, _09631_, _03774_);
  nor (_09633_, _09575_, _03774_);
  or (_09634_, _09633_, _09632_);
  and (_09635_, _09634_, _04060_);
  nor (_09636_, _09635_, _09564_);
  nand (_09637_, _09636_, _43152_);
  or (_09638_, _43152_, \oc8051_golden_model_1.TMOD [7]);
  and (_09639_, _09638_, _41894_);
  and (_40692_, _09639_, _09637_);
  not (_09640_, \oc8051_golden_model_1.IE [7]);
  nor (_09641_, _05494_, _09640_);
  and (_09642_, _06557_, _05494_);
  nor (_09643_, _09642_, _09641_);
  nor (_09644_, _09643_, _04792_);
  and (_09645_, _05494_, \oc8051_golden_model_1.ACC [7]);
  nor (_09646_, _09645_, _09641_);
  nor (_09647_, _09646_, _04708_);
  nor (_09648_, _04707_, _09640_);
  or (_09649_, _09648_, _09647_);
  and (_09650_, _09649_, _04722_);
  and (_09651_, _06160_, _05494_);
  nor (_09652_, _09651_, _09641_);
  nor (_09653_, _09652_, _04722_);
  or (_09654_, _09653_, _09650_);
  and (_09655_, _09654_, _03764_);
  nor (_09656_, _06103_, _09640_);
  and (_09657_, _06148_, _06103_);
  nor (_09658_, _09657_, _09656_);
  nor (_09659_, _09658_, _03764_);
  or (_09660_, _09659_, _03848_);
  or (_09661_, _09660_, _09655_);
  and (_09662_, _05568_, _05494_);
  nor (_09663_, _09662_, _09641_);
  nand (_09664_, _09663_, _03848_);
  and (_09665_, _09664_, _09661_);
  and (_09666_, _09665_, _03855_);
  nor (_09667_, _09646_, _03855_);
  or (_09668_, _09667_, _09666_);
  and (_09669_, _09668_, _03760_);
  and (_09670_, _06121_, _06103_);
  nor (_09671_, _09670_, _09656_);
  nor (_09672_, _09671_, _03760_);
  or (_09673_, _09672_, _09669_);
  and (_09674_, _09673_, _03753_);
  nor (_09675_, _09656_, _06147_);
  nor (_09676_, _09675_, _09658_);
  and (_09677_, _09676_, _03752_);
  or (_09678_, _09677_, _09674_);
  and (_09679_, _09678_, _03747_);
  not (_09680_, _06103_);
  nor (_09681_, _06143_, _09680_);
  nor (_09682_, _09681_, _09656_);
  nor (_09683_, _09682_, _03747_);
  or (_09684_, _09683_, _07927_);
  or (_09685_, _09684_, _09679_);
  and (_09686_, _06248_, _05494_);
  nor (_09687_, _09641_, _03738_);
  not (_09688_, _09687_);
  nor (_09689_, _09688_, _09686_);
  and (_09690_, _09663_, _08474_);
  or (_09691_, _09690_, _03455_);
  nor (_09692_, _09691_, _09689_);
  and (_09693_, _09692_, _09685_);
  not (_09694_, _05494_);
  nor (_09695_, _06536_, _09694_);
  nor (_09696_, _09695_, _09641_);
  nor (_09697_, _09696_, _03820_);
  or (_09698_, _09697_, _09693_);
  and (_09699_, _09698_, _04778_);
  and (_09700_, _06348_, _05494_);
  nor (_09701_, _09700_, _09641_);
  nor (_09702_, _09701_, _04778_);
  or (_09703_, _09702_, _09699_);
  nor (_09704_, _09703_, _03897_);
  and (_09705_, _06549_, _05494_);
  or (_09706_, _09641_, _04790_);
  nor (_09707_, _09706_, _09705_);
  or (_09708_, _09707_, _04018_);
  nor (_09709_, _09708_, _09704_);
  nor (_09710_, _09709_, _09644_);
  nor (_09711_, _09710_, _03908_);
  nor (_09712_, _09641_, _05571_);
  not (_09713_, _09712_);
  nor (_09714_, _09701_, _03909_);
  and (_09715_, _09714_, _09713_);
  nor (_09716_, _09715_, _09711_);
  nor (_09717_, _09716_, _04027_);
  nor (_09718_, _09646_, _04785_);
  and (_09719_, _09718_, _09713_);
  or (_09720_, _09719_, _09717_);
  and (_09721_, _09720_, _06567_);
  nor (_09722_, _06547_, _09694_);
  nor (_09723_, _09722_, _09641_);
  nor (_09724_, _09723_, _06567_);
  or (_09725_, _09724_, _09721_);
  and (_09726_, _09725_, _06572_);
  nor (_09727_, _06556_, _09694_);
  nor (_09728_, _09727_, _09641_);
  nor (_09729_, _09728_, _06572_);
  or (_09730_, _09729_, _09726_);
  and (_09731_, _09730_, _03774_);
  nor (_09732_, _09652_, _03774_);
  or (_09733_, _09732_, _09731_);
  and (_09734_, _09733_, _03375_);
  nor (_09735_, _09671_, _03375_);
  or (_09736_, _09735_, _09734_);
  and (_09737_, _09736_, _04060_);
  and (_09738_, _06077_, _05494_);
  nor (_09739_, _09738_, _09641_);
  nor (_09740_, _09739_, _04060_);
  or (_09741_, _09740_, _09737_);
  or (_09742_, _09741_, _43156_);
  or (_09743_, _43152_, \oc8051_golden_model_1.IE [7]);
  and (_09744_, _09743_, _41894_);
  and (_40693_, _09744_, _09742_);
  not (_09745_, \oc8051_golden_model_1.IP [7]);
  nor (_09746_, _05437_, _09745_);
  and (_09747_, _06557_, _05437_);
  nor (_09748_, _09747_, _09746_);
  nor (_09749_, _09748_, _04792_);
  and (_09750_, _05437_, \oc8051_golden_model_1.ACC [7]);
  nor (_09751_, _09750_, _09746_);
  nor (_09752_, _09751_, _04708_);
  nor (_09753_, _04707_, _09745_);
  or (_09754_, _09753_, _09752_);
  and (_09755_, _09754_, _04722_);
  and (_09756_, _06160_, _05437_);
  nor (_09757_, _09756_, _09746_);
  nor (_09758_, _09757_, _04722_);
  or (_09759_, _09758_, _09755_);
  and (_09760_, _09759_, _03764_);
  nor (_09761_, _06091_, _09745_);
  and (_09762_, _06148_, _06091_);
  nor (_09763_, _09762_, _09761_);
  nor (_09764_, _09763_, _03764_);
  or (_09765_, _09764_, _03848_);
  or (_09766_, _09765_, _09760_);
  and (_09767_, _05568_, _05437_);
  nor (_09768_, _09767_, _09746_);
  nand (_09769_, _09768_, _03848_);
  and (_09770_, _09769_, _09766_);
  and (_09771_, _09770_, _03855_);
  nor (_09772_, _09751_, _03855_);
  or (_09773_, _09772_, _09771_);
  and (_09774_, _09773_, _03760_);
  and (_09775_, _06121_, _06091_);
  nor (_09776_, _09775_, _09761_);
  nor (_09777_, _09776_, _03760_);
  or (_09778_, _09777_, _03752_);
  or (_09779_, _09778_, _09774_);
  nor (_09780_, _09761_, _06147_);
  nor (_09781_, _09780_, _09763_);
  or (_09782_, _09781_, _03753_);
  and (_09783_, _09782_, _03747_);
  and (_09784_, _09783_, _09779_);
  not (_09785_, _06091_);
  nor (_09786_, _06143_, _09785_);
  nor (_09787_, _09786_, _09761_);
  nor (_09788_, _09787_, _03747_);
  or (_09789_, _09788_, _07927_);
  or (_09790_, _09789_, _09784_);
  and (_09791_, _06248_, _05437_);
  nor (_09792_, _09746_, _03738_);
  not (_09793_, _09792_);
  nor (_09794_, _09793_, _09791_);
  and (_09795_, _09768_, _08474_);
  or (_09796_, _09795_, _03455_);
  nor (_09797_, _09796_, _09794_);
  and (_09798_, _09797_, _09790_);
  not (_09799_, _05437_);
  nor (_09800_, _06536_, _09799_);
  nor (_09801_, _09800_, _09746_);
  nor (_09802_, _09801_, _03820_);
  or (_09803_, _09802_, _09798_);
  and (_09804_, _09803_, _04778_);
  and (_09805_, _06348_, _05437_);
  nor (_09806_, _09805_, _09746_);
  nor (_09807_, _09806_, _04778_);
  or (_09808_, _09807_, _09804_);
  nor (_09809_, _09808_, _03897_);
  and (_09810_, _06549_, _05437_);
  or (_09811_, _09746_, _04790_);
  nor (_09812_, _09811_, _09810_);
  or (_09813_, _09812_, _04018_);
  nor (_09814_, _09813_, _09809_);
  nor (_09815_, _09814_, _09749_);
  nor (_09816_, _09815_, _03908_);
  nor (_09817_, _09746_, _05571_);
  not (_09818_, _09817_);
  nor (_09819_, _09806_, _03909_);
  and (_09820_, _09819_, _09818_);
  nor (_09821_, _09820_, _09816_);
  nor (_09822_, _09821_, _04027_);
  nor (_09823_, _09751_, _04785_);
  and (_09824_, _09823_, _09818_);
  nor (_09825_, _09824_, _03914_);
  not (_09826_, _09825_);
  nor (_09827_, _09826_, _09822_);
  nor (_09828_, _06547_, _09799_);
  or (_09829_, _09746_, _06567_);
  nor (_09830_, _09829_, _09828_);
  or (_09831_, _09830_, _04011_);
  nor (_09832_, _09831_, _09827_);
  nor (_09833_, _06556_, _09799_);
  nor (_09834_, _09833_, _09746_);
  nor (_09835_, _09834_, _06572_);
  or (_09836_, _09835_, _09832_);
  and (_09837_, _09836_, _03774_);
  nor (_09838_, _09757_, _03774_);
  or (_09839_, _09838_, _09837_);
  and (_09840_, _09839_, _03375_);
  nor (_09841_, _09776_, _03375_);
  or (_09842_, _09841_, _09840_);
  and (_09843_, _09842_, _04060_);
  and (_09844_, _06077_, _05437_);
  nor (_09845_, _09844_, _09746_);
  nor (_09846_, _09845_, _04060_);
  or (_09847_, _09846_, _09843_);
  or (_09848_, _09847_, _43156_);
  or (_09849_, _43152_, \oc8051_golden_model_1.IP [7]);
  and (_09850_, _09849_, _41894_);
  and (_40695_, _09850_, _09848_);
  or (_09851_, _43152_, \oc8051_golden_model_1.DPL [7]);
  and (_09852_, _09851_, _41894_);
  not (_09853_, \oc8051_golden_model_1.DPL [7]);
  nor (_09854_, _05513_, _09853_);
  and (_09855_, _06557_, _05513_);
  or (_09856_, _09855_, _09854_);
  and (_09857_, _09856_, _04018_);
  and (_09858_, _06348_, _05513_);
  or (_09859_, _09858_, _09854_);
  or (_09860_, _09859_, _04778_);
  not (_09861_, _03921_);
  and (_09862_, _06160_, _05513_);
  or (_09863_, _09862_, _09854_);
  or (_09864_, _09863_, _04722_);
  and (_09865_, _05513_, \oc8051_golden_model_1.ACC [7]);
  or (_09866_, _09865_, _09854_);
  and (_09867_, _09866_, _04707_);
  nor (_09868_, _04707_, _09853_);
  or (_09869_, _09868_, _03850_);
  or (_09870_, _09869_, _09867_);
  and (_09871_, _09870_, _04733_);
  and (_09872_, _09871_, _09864_);
  and (_09873_, _05568_, _05513_);
  or (_09874_, _09873_, _09854_);
  and (_09875_, _09874_, _03848_);
  or (_09876_, _09875_, _03854_);
  or (_09877_, _09876_, _09872_);
  and (_09878_, _03821_, _03423_);
  not (_09879_, _09878_);
  or (_09880_, _09866_, _03855_);
  and (_09881_, _09880_, _09879_);
  and (_09882_, _09881_, _09877_);
  and (_09883_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_09884_, _09883_, \oc8051_golden_model_1.DPL [2]);
  and (_09885_, _09884_, \oc8051_golden_model_1.DPL [3]);
  and (_09886_, _09885_, \oc8051_golden_model_1.DPL [4]);
  and (_09887_, _09886_, \oc8051_golden_model_1.DPL [5]);
  and (_09888_, _09887_, \oc8051_golden_model_1.DPL [6]);
  nor (_09889_, _09888_, \oc8051_golden_model_1.DPL [7]);
  and (_09890_, _09888_, \oc8051_golden_model_1.DPL [7]);
  nor (_09891_, _09890_, _09889_);
  and (_09892_, _09891_, _09878_);
  or (_09893_, _09892_, _09882_);
  and (_09894_, _09893_, _09861_);
  nor (_09895_, _06342_, _09861_);
  or (_09896_, _09895_, _07927_);
  or (_09897_, _09896_, _09894_);
  and (_09898_, _06248_, _05513_);
  or (_09899_, _09854_, _03738_);
  or (_09900_, _09899_, _09898_);
  or (_09901_, _09874_, _07925_);
  and (_09902_, _09901_, _03820_);
  and (_09903_, _09902_, _09900_);
  and (_09904_, _09903_, _09897_);
  not (_09905_, _05513_);
  nor (_09906_, _06536_, _09905_);
  or (_09907_, _09906_, _09854_);
  and (_09908_, _09907_, _03455_);
  or (_09909_, _09908_, _03903_);
  or (_09910_, _09909_, _09904_);
  and (_09911_, _09910_, _09860_);
  or (_09912_, _09911_, _03897_);
  and (_09913_, _06549_, _05513_);
  or (_09914_, _09913_, _09854_);
  or (_09915_, _09914_, _04790_);
  and (_09916_, _09915_, _04792_);
  and (_09917_, _09916_, _09912_);
  or (_09918_, _09917_, _09857_);
  and (_09919_, _09918_, _03909_);
  or (_09920_, _09854_, _05571_);
  and (_09921_, _09859_, _03908_);
  and (_09922_, _09921_, _09920_);
  or (_09923_, _09922_, _09919_);
  and (_09924_, _09923_, _04785_);
  and (_09925_, _09866_, _04027_);
  and (_09926_, _09925_, _09920_);
  or (_09927_, _09926_, _03914_);
  or (_09928_, _09927_, _09924_);
  nor (_09929_, _06547_, _09905_);
  or (_09930_, _09854_, _06567_);
  or (_09931_, _09930_, _09929_);
  and (_09932_, _09931_, _06572_);
  and (_09933_, _09932_, _09928_);
  nor (_09934_, _06556_, _09905_);
  or (_09935_, _09934_, _09854_);
  and (_09936_, _09935_, _04011_);
  or (_09937_, _09936_, _03773_);
  or (_09938_, _09937_, _09933_);
  or (_09939_, _09863_, _03774_);
  and (_09940_, _09939_, _04060_);
  and (_09941_, _09940_, _09938_);
  and (_09942_, _06077_, _05513_);
  or (_09943_, _09942_, _09854_);
  and (_09944_, _09943_, _03772_);
  or (_09945_, _09944_, _43156_);
  or (_09946_, _09945_, _09941_);
  and (_40696_, _09946_, _09852_);
  or (_09947_, _43152_, \oc8051_golden_model_1.DPH [7]);
  and (_09948_, _09947_, _41894_);
  not (_09949_, \oc8051_golden_model_1.DPH [7]);
  nor (_09950_, _05509_, _09949_);
  and (_09951_, _06557_, _05509_);
  or (_09952_, _09951_, _09950_);
  and (_09953_, _09952_, _04018_);
  and (_09954_, _06348_, _05509_);
  or (_09955_, _09954_, _09950_);
  or (_09956_, _09955_, _04778_);
  and (_09957_, _06160_, _05509_);
  or (_09958_, _09957_, _09950_);
  or (_09959_, _09958_, _04722_);
  and (_09960_, _05509_, \oc8051_golden_model_1.ACC [7]);
  or (_09961_, _09960_, _09950_);
  and (_09962_, _09961_, _04707_);
  nor (_09963_, _04707_, _09949_);
  or (_09964_, _09963_, _03850_);
  or (_09965_, _09964_, _09962_);
  and (_09966_, _09965_, _04733_);
  and (_09967_, _09966_, _09959_);
  and (_09968_, _05568_, _05509_);
  or (_09969_, _09968_, _09950_);
  and (_09970_, _09969_, _03848_);
  or (_09971_, _09970_, _03854_);
  or (_09972_, _09971_, _09967_);
  or (_09973_, _09961_, _03855_);
  and (_09974_, _09973_, _09879_);
  and (_09975_, _09974_, _09972_);
  not (_09976_, \oc8051_golden_model_1.DPH [6]);
  and (_09977_, _09890_, \oc8051_golden_model_1.DPH [0]);
  and (_09978_, _09977_, \oc8051_golden_model_1.DPH [1]);
  and (_09979_, _09978_, \oc8051_golden_model_1.DPH [2]);
  and (_09980_, _09979_, \oc8051_golden_model_1.DPH [3]);
  and (_09981_, _09980_, \oc8051_golden_model_1.DPH [4]);
  nand (_09982_, _09981_, \oc8051_golden_model_1.DPH [5]);
  nor (_09983_, _09982_, _09976_);
  nor (_09984_, _09983_, _09949_);
  and (_09985_, _09983_, _09949_);
  or (_09986_, _09985_, _09984_);
  and (_09987_, _09986_, _09878_);
  or (_09988_, _09987_, _09975_);
  and (_09989_, _09988_, _09861_);
  and (_09990_, _03921_, _03647_);
  or (_09991_, _09990_, _07927_);
  or (_09992_, _09991_, _09989_);
  and (_09993_, _06248_, _05509_);
  or (_09994_, _09950_, _03738_);
  or (_09995_, _09994_, _09993_);
  or (_09996_, _09969_, _07925_);
  and (_09997_, _09996_, _03820_);
  and (_09998_, _09997_, _09995_);
  and (_09999_, _09998_, _09992_);
  not (_10000_, _05509_);
  nor (_10001_, _06536_, _10000_);
  or (_10002_, _10001_, _09950_);
  and (_10003_, _10002_, _03455_);
  or (_10004_, _10003_, _03903_);
  or (_10005_, _10004_, _09999_);
  and (_10006_, _10005_, _09956_);
  or (_10007_, _10006_, _03897_);
  and (_10008_, _06549_, _05509_);
  or (_10009_, _10008_, _09950_);
  or (_10010_, _10009_, _04790_);
  and (_10011_, _10010_, _04792_);
  and (_10012_, _10011_, _10007_);
  or (_10013_, _10012_, _09953_);
  and (_10014_, _10013_, _03909_);
  or (_10015_, _09950_, _05571_);
  and (_10016_, _09955_, _03908_);
  and (_10017_, _10016_, _10015_);
  or (_10018_, _10017_, _10014_);
  and (_10019_, _10018_, _04785_);
  and (_10020_, _09961_, _04027_);
  and (_10021_, _10020_, _10015_);
  or (_10022_, _10021_, _03914_);
  or (_10023_, _10022_, _10019_);
  nor (_10024_, _06547_, _10000_);
  or (_10025_, _09950_, _06567_);
  or (_10026_, _10025_, _10024_);
  and (_10027_, _10026_, _06572_);
  and (_10028_, _10027_, _10023_);
  nor (_10029_, _06556_, _10000_);
  or (_10030_, _10029_, _09950_);
  and (_10031_, _10030_, _04011_);
  or (_10032_, _10031_, _03773_);
  or (_10033_, _10032_, _10028_);
  or (_10034_, _09958_, _03774_);
  and (_10035_, _10034_, _04060_);
  and (_10036_, _10035_, _10033_);
  and (_10037_, _06077_, _05509_);
  or (_10038_, _10037_, _09950_);
  and (_10039_, _10038_, _03772_);
  or (_10040_, _10039_, _43156_);
  or (_10041_, _10040_, _10036_);
  and (_40697_, _10041_, _09948_);
  and (_10042_, _03412_, _03373_);
  and (_10043_, _06253_, _03103_);
  and (_10044_, _10043_, \oc8051_golden_model_1.PC [7]);
  and (_10045_, _10044_, \oc8051_golden_model_1.PC [8]);
  and (_10046_, _10045_, \oc8051_golden_model_1.PC [9]);
  and (_10047_, _10046_, \oc8051_golden_model_1.PC [10]);
  and (_10048_, _10047_, \oc8051_golden_model_1.PC [11]);
  and (_10049_, _10048_, \oc8051_golden_model_1.PC [12]);
  and (_10050_, _10049_, \oc8051_golden_model_1.PC [13]);
  nand (_10051_, _10050_, \oc8051_golden_model_1.PC [14]);
  nand (_10052_, _10051_, _06983_);
  or (_10053_, _10051_, _06983_);
  and (_10054_, _10053_, _10052_);
  and (_10055_, _10054_, _10042_);
  nor (_10056_, _08733_, _03779_);
  not (_10057_, _10056_);
  not (_10058_, _08691_);
  and (_10059_, _07999_, _10058_);
  or (_10060_, _10059_, _10054_);
  and (_10061_, _08599_, _08119_);
  or (_10062_, _10061_, _10054_);
  and (_10063_, _03392_, _03373_);
  not (_10064_, _10063_);
  nor (_10065_, _04011_, _03393_);
  or (_10066_, _10065_, _07003_);
  and (_10067_, _10066_, _10064_);
  or (_10068_, _08573_, _08568_);
  not (_10069_, _10068_);
  not (_10070_, _08563_);
  and (_10071_, _10070_, _08567_);
  and (_10072_, _10071_, _10069_);
  or (_10073_, _10072_, _10054_);
  and (_10074_, _03387_, _03373_);
  not (_10075_, _10074_);
  nor (_10076_, _04027_, _03388_);
  or (_10077_, _10076_, _07003_);
  and (_10078_, _10077_, _10075_);
  nor (_10079_, _08530_, _04016_);
  not (_10080_, _10079_);
  and (_10081_, _08502_, _08520_);
  and (_10082_, _10081_, _08514_);
  or (_10083_, _10082_, _10054_);
  and (_10084_, _06993_, _03455_);
  nor (_10085_, _08320_, _03883_);
  not (_10086_, _10085_);
  and (_10087_, _08153_, _08248_);
  or (_10088_, _10087_, _10054_);
  and (_10089_, _03454_, _03821_);
  not (_10090_, _10089_);
  nor (_10091_, _09878_, _07399_);
  and (_10092_, _10091_, _10090_);
  not (_10093_, _10092_);
  and (_10094_, _10093_, _10054_);
  and (_10095_, _06987_, \oc8051_golden_model_1.PC [12]);
  and (_10096_, _10095_, \oc8051_golden_model_1.PC [13]);
  and (_10097_, _10096_, \oc8051_golden_model_1.PC [14]);
  nor (_10098_, _10096_, \oc8051_golden_model_1.PC [14]);
  nor (_10099_, _10098_, _10097_);
  not (_10100_, _10099_);
  nor (_10101_, _10100_, _06342_);
  and (_10102_, _10100_, _06342_);
  nor (_10103_, _10102_, _10101_);
  nor (_10104_, _10095_, \oc8051_golden_model_1.PC [13]);
  nor (_10105_, _10104_, _10096_);
  not (_10106_, _10105_);
  nor (_10107_, _10106_, _06342_);
  and (_10108_, _10106_, _06342_);
  nor (_10109_, _06987_, \oc8051_golden_model_1.PC [12]);
  nor (_10110_, _10109_, _10095_);
  not (_10111_, _10110_);
  nor (_10112_, _10111_, _06342_);
  nor (_10113_, _06985_, \oc8051_golden_model_1.PC [10]);
  nor (_10114_, _10113_, _06986_);
  not (_10115_, _10114_);
  nor (_10116_, _10115_, _06342_);
  not (_10117_, _10116_);
  nor (_10118_, _06986_, \oc8051_golden_model_1.PC [11]);
  nor (_10119_, _10118_, _06987_);
  not (_10120_, _10119_);
  nor (_10121_, _10120_, _06342_);
  and (_10122_, _10120_, _06342_);
  nor (_10123_, _10122_, _10121_);
  and (_10124_, _10115_, _06342_);
  nor (_10125_, _10124_, _10116_);
  and (_10126_, _10125_, _10123_);
  nor (_10127_, _06984_, \oc8051_golden_model_1.PC [9]);
  nor (_10128_, _10127_, _06985_);
  not (_10129_, _10128_);
  nor (_10130_, _10129_, _06342_);
  and (_10131_, _10129_, _06342_);
  nor (_10132_, _10131_, _10130_);
  nor (_10133_, _06936_, _06342_);
  and (_10134_, _06936_, _06342_);
  and (_10135_, _06931_, _06252_);
  nor (_10136_, _10135_, \oc8051_golden_model_1.PC [6]);
  nor (_10137_, _10136_, _06932_);
  not (_10138_, _10137_);
  nor (_10139_, _10138_, _06379_);
  and (_10140_, _10138_, _06379_);
  nor (_10141_, _10140_, _10139_);
  and (_10142_, _06931_, \oc8051_golden_model_1.PC [4]);
  nor (_10143_, _10142_, \oc8051_golden_model_1.PC [5]);
  nor (_10144_, _10143_, _10135_);
  not (_10145_, _10144_);
  nor (_10146_, _10145_, _06411_);
  and (_10147_, _10145_, _06411_);
  nor (_10148_, _06931_, \oc8051_golden_model_1.PC [4]);
  nor (_10149_, _10148_, _10142_);
  not (_10150_, _10149_);
  nor (_10151_, _10150_, _06442_);
  and (_10152_, _03123_, \oc8051_golden_model_1.PC [2]);
  nor (_10153_, _10152_, \oc8051_golden_model_1.PC [3]);
  nor (_10154_, _10153_, _06931_);
  not (_10155_, _10154_);
  nor (_10156_, _10155_, _04005_);
  and (_10157_, _10155_, _04005_);
  nor (_10158_, _03123_, \oc8051_golden_model_1.PC [2]);
  nor (_10159_, _10158_, _10152_);
  not (_10160_, _10159_);
  nor (_10161_, _10160_, _04180_);
  nor (_10162_, _04595_, _03948_);
  nor (_10163_, _04382_, \oc8051_golden_model_1.PC [0]);
  and (_10164_, _04595_, _03948_);
  nor (_10165_, _10164_, _10162_);
  and (_10166_, _10165_, _10163_);
  nor (_10167_, _10166_, _10162_);
  and (_10168_, _10160_, _04180_);
  nor (_10169_, _10168_, _10161_);
  not (_10170_, _10169_);
  nor (_10171_, _10170_, _10167_);
  nor (_10172_, _10171_, _10161_);
  nor (_10173_, _10172_, _10157_);
  nor (_10174_, _10173_, _10156_);
  and (_10175_, _10150_, _06442_);
  nor (_10176_, _10175_, _10151_);
  not (_10177_, _10176_);
  nor (_10178_, _10177_, _10174_);
  nor (_10179_, _10178_, _10151_);
  nor (_10180_, _10179_, _10147_);
  nor (_10181_, _10180_, _10146_);
  not (_10182_, _10181_);
  and (_10183_, _10182_, _10141_);
  nor (_10184_, _10183_, _10139_);
  nor (_10185_, _10184_, _10134_);
  or (_10186_, _10185_, _10133_);
  nor (_10187_, _06933_, \oc8051_golden_model_1.PC [8]);
  nor (_10188_, _10187_, _06984_);
  not (_10189_, _10188_);
  nor (_10190_, _10189_, _06342_);
  and (_10191_, _10189_, _06342_);
  nor (_10192_, _10191_, _10190_);
  and (_10193_, _10192_, _10186_);
  and (_10194_, _10193_, _10132_);
  and (_10195_, _10194_, _10126_);
  nor (_10196_, _10190_, _10130_);
  not (_10197_, _10196_);
  and (_10198_, _10197_, _10126_);
  or (_10199_, _10198_, _10121_);
  nor (_10200_, _10199_, _10195_);
  and (_10201_, _10200_, _10117_);
  and (_10202_, _10111_, _06342_);
  nor (_10203_, _10202_, _10112_);
  not (_10204_, _10203_);
  nor (_10205_, _10204_, _10201_);
  nor (_10206_, _10205_, _10112_);
  nor (_10207_, _10206_, _10108_);
  nor (_10208_, _10207_, _10107_);
  not (_10209_, _10208_);
  and (_10210_, _10209_, _10103_);
  nor (_10211_, _10210_, _10101_);
  not (_10212_, _06993_);
  and (_10213_, _10212_, _06342_);
  nor (_10214_, _10212_, _06342_);
  nor (_10215_, _10214_, _10213_);
  and (_10216_, _10215_, _10211_);
  nor (_10217_, _10215_, _10211_);
  or (_10218_, _10217_, _10216_);
  nor (_10219_, _06248_, _05421_);
  nor (_10220_, _10219_, _06291_);
  nor (_10221_, _06641_, _03810_);
  and (_10222_, _06641_, _03810_);
  nor (_10223_, _10222_, _10221_);
  and (_10224_, _10223_, _10220_);
  and (_10225_, _06968_, _04093_);
  and (_10226_, _06873_, _05426_);
  nor (_10227_, _10226_, _10225_);
  and (_10228_, _06918_, _05419_);
  and (_10229_, _06969_, _04526_);
  nor (_10230_, _10229_, _10228_);
  and (_10231_, _10230_, _10227_);
  and (_10232_, _10231_, _10224_);
  and (_10233_, _06779_, _03812_);
  not (_10234_, _10233_);
  or (_10235_, _06779_, _03812_);
  and (_10236_, _10235_, _10234_);
  and (_10237_, _06965_, _04139_);
  and (_10238_, _06824_, _05243_);
  nor (_10239_, _10238_, _10237_);
  and (_10240_, _10239_, _10236_);
  or (_10241_, _06733_, _03716_);
  and (_10242_, _06961_, _04563_);
  and (_10243_, _06688_, _04835_);
  nor (_10244_, _10243_, _10242_);
  and (_10245_, _10244_, _10241_);
  or (_10246_, _06962_, _03715_);
  and (_10247_, _10246_, _10245_);
  and (_10248_, _10247_, _10240_);
  and (_10249_, _10248_, _10232_);
  not (_10250_, _10249_);
  and (_10251_, _10250_, _10218_);
  and (_10252_, _10249_, _06993_);
  or (_10253_, _10252_, _10251_);
  and (_10254_, _10253_, _03925_);
  not (_10255_, _03434_);
  nor (_10256_, _03758_, _10255_);
  and (_10257_, _10256_, _03760_);
  or (_10258_, _10257_, _07003_);
  and (_10259_, _07003_, _03854_);
  and (_10260_, _06152_, _05764_);
  and (_10261_, _10260_, _05621_);
  not (_10262_, _05716_);
  and (_10263_, _06070_, _10262_);
  and (_10264_, _10263_, _05669_);
  and (_10265_, _10264_, _10261_);
  or (_10266_, _10265_, _10218_);
  nand (_10267_, _10265_, _10212_);
  and (_10268_, _10267_, _03850_);
  and (_10269_, _10268_, _10266_);
  and (_10270_, _06998_, \oc8051_golden_model_1.PC [12]);
  and (_10271_, _10270_, \oc8051_golden_model_1.PC [13]);
  and (_10272_, _10271_, \oc8051_golden_model_1.PC [14]);
  nor (_10273_, _10271_, \oc8051_golden_model_1.PC [14]);
  nor (_10274_, _10273_, _10272_);
  and (_10275_, _10274_, _03647_);
  nor (_10276_, _10274_, _03647_);
  nor (_10277_, _10276_, _10275_);
  nor (_10278_, _10270_, \oc8051_golden_model_1.PC [13]);
  nor (_10279_, _10278_, _10271_);
  and (_10280_, _10279_, _03647_);
  nor (_10281_, _10279_, _03647_);
  nor (_10282_, _06998_, \oc8051_golden_model_1.PC [12]);
  nor (_10283_, _10282_, _10270_);
  and (_10284_, _10283_, _03647_);
  nor (_10285_, _06997_, \oc8051_golden_model_1.PC [11]);
  nor (_10286_, _10285_, _06998_);
  and (_10287_, _10286_, _03647_);
  nor (_10288_, _10286_, _03647_);
  nor (_10289_, _10288_, _10287_);
  nor (_10290_, _06996_, \oc8051_golden_model_1.PC [10]);
  nor (_10291_, _10290_, _06997_);
  and (_10292_, _10291_, _03647_);
  nor (_10293_, _10291_, _03647_);
  nor (_10294_, _10293_, _10292_);
  and (_10295_, _10294_, _10289_);
  nor (_10296_, _06995_, \oc8051_golden_model_1.PC [9]);
  nor (_10297_, _10296_, _06996_);
  and (_10298_, _10297_, _03647_);
  nor (_10299_, _10297_, _03647_);
  nor (_10300_, _10299_, _10298_);
  and (_10301_, _06257_, _03647_);
  nor (_10302_, _06257_, _03647_);
  and (_10303_, _06252_, _03550_);
  nor (_10304_, _10303_, \oc8051_golden_model_1.PC [6]);
  nor (_10305_, _10304_, _06254_);
  not (_10306_, _10305_);
  nor (_10307_, _10306_, _03810_);
  and (_10308_, _10306_, _03810_);
  nor (_10309_, _10308_, _10307_);
  and (_10310_, _03550_, \oc8051_golden_model_1.PC [4]);
  nor (_10311_, _10310_, \oc8051_golden_model_1.PC [5]);
  nor (_10312_, _10311_, _10303_);
  not (_10313_, _10312_);
  nor (_10314_, _10313_, _04093_);
  and (_10315_, _10313_, _04093_);
  nor (_10316_, _03550_, \oc8051_golden_model_1.PC [4]);
  nor (_10317_, _10316_, _10310_);
  not (_10318_, _10317_);
  nor (_10319_, _10318_, _04526_);
  nor (_10320_, _03678_, _03938_);
  and (_10321_, _03678_, _03938_);
  nor (_10322_, _04139_, _03511_);
  nor (_10323_, _04563_, \oc8051_golden_model_1.PC [1]);
  nor (_10324_, _03715_, _03119_);
  and (_10325_, _04563_, \oc8051_golden_model_1.PC [1]);
  nor (_10326_, _10325_, _10323_);
  and (_10327_, _10326_, _10324_);
  nor (_10328_, _10327_, _10323_);
  and (_10329_, _04139_, _03511_);
  nor (_10330_, _10329_, _10322_);
  not (_10331_, _10330_);
  nor (_10332_, _10331_, _10328_);
  nor (_10333_, _10332_, _10322_);
  nor (_10334_, _10333_, _10321_);
  nor (_10335_, _10334_, _10320_);
  and (_10336_, _10318_, _04526_);
  nor (_10337_, _10336_, _10319_);
  not (_10338_, _10337_);
  nor (_10339_, _10338_, _10335_);
  nor (_10340_, _10339_, _10319_);
  nor (_10341_, _10340_, _10315_);
  nor (_10342_, _10341_, _10314_);
  not (_10343_, _10342_);
  and (_10344_, _10343_, _10309_);
  nor (_10345_, _10344_, _10307_);
  nor (_10346_, _10345_, _10302_);
  or (_10347_, _10346_, _10301_);
  nor (_10348_, _06255_, \oc8051_golden_model_1.PC [8]);
  nor (_10349_, _10348_, _06995_);
  and (_10350_, _10349_, _03647_);
  nor (_10351_, _10349_, _03647_);
  nor (_10352_, _10351_, _10350_);
  and (_10353_, _10352_, _10347_);
  and (_10354_, _10353_, _10300_);
  and (_10355_, _10354_, _10295_);
  nor (_10356_, _10350_, _10298_);
  not (_10357_, _10356_);
  and (_10358_, _10357_, _10295_);
  or (_10359_, _10358_, _10292_);
  or (_10360_, _10359_, _10355_);
  nor (_10361_, _10360_, _10287_);
  nor (_10362_, _10283_, _03647_);
  nor (_10363_, _10362_, _10284_);
  not (_10364_, _10363_);
  nor (_10365_, _10364_, _10361_);
  nor (_10366_, _10365_, _10284_);
  nor (_10367_, _10366_, _10281_);
  nor (_10368_, _10367_, _10280_);
  not (_10369_, _10368_);
  and (_10370_, _10369_, _10277_);
  nor (_10371_, _10370_, _10275_);
  nor (_10372_, _07003_, _03647_);
  and (_10373_, _07003_, _03647_);
  nor (_10374_, _10373_, _10372_);
  and (_10375_, _10374_, _10371_);
  nor (_10376_, _10374_, _10371_);
  or (_10377_, _10376_, _10375_);
  and (_10378_, _06126_, _06124_);
  not (_10379_, _04900_);
  and (_10380_, _10379_, _04700_);
  and (_10381_, _06951_, _10380_);
  and (_10382_, _10381_, _10378_);
  not (_10383_, _10382_);
  and (_10384_, _10383_, _10377_);
  and (_10385_, _10382_, _07003_);
  or (_10386_, _10385_, _10384_);
  and (_10387_, _10386_, _04267_);
  and (_10388_, _10054_, _04263_);
  not (_10389_, _04230_);
  and (_10390_, _07003_, _03420_);
  or (_10391_, _10390_, _10389_);
  and (_10392_, _10054_, _05011_);
  nor (_10393_, _05011_, _06983_);
  or (_10394_, _10393_, _04707_);
  or (_10395_, _10394_, _10392_);
  and (_10396_, _10395_, _10391_);
  or (_10397_, _10396_, _10388_);
  and (_10398_, _10397_, _03770_);
  nand (_10399_, _07003_, _03768_);
  not (_10400_, _08169_);
  nor (_10401_, _08159_, _08162_);
  and (_10402_, _10401_, _10400_);
  nand (_10403_, _10402_, _10399_);
  or (_10404_, _10403_, _10398_);
  or (_10405_, _10402_, _10054_);
  and (_10406_, _10405_, _04266_);
  and (_10407_, _10406_, _10404_);
  or (_10408_, _10407_, _04716_);
  or (_10409_, _10408_, _10387_);
  and (_10410_, _10409_, _04722_);
  and (_10411_, _03762_, _03423_);
  nor (_10412_, _10411_, _08179_);
  not (_10413_, _10412_);
  or (_10414_, _10413_, _10410_);
  or (_10415_, _10414_, _10269_);
  and (_10416_, _03856_, _03431_);
  and (_10417_, _10412_, _04717_);
  or (_10418_, _10417_, _10054_);
  and (_10419_, _10418_, _10416_);
  and (_10420_, _10419_, _10415_);
  and (_10421_, _08157_, _04739_);
  not (_10422_, _07003_);
  or (_10423_, _10416_, _10422_);
  nand (_10424_, _10423_, _10421_);
  or (_10425_, _10424_, _10420_);
  or (_10426_, _10421_, _10054_);
  and (_10427_, _10426_, _03855_);
  and (_10428_, _10427_, _10425_);
  or (_10429_, _10428_, _10259_);
  and (_10430_, _03757_, _03423_);
  nor (_10431_, _10430_, _08224_);
  and (_10432_, _10431_, _10429_);
  not (_10433_, _10257_);
  not (_10434_, _10431_);
  and (_10435_, _10434_, _10054_);
  or (_10436_, _10435_, _10433_);
  or (_10437_, _10436_, _10432_);
  and (_10438_, _10437_, _10258_);
  and (_10439_, _07919_, _04255_);
  nor (_10440_, _10439_, _03427_);
  nor (_10441_, _10440_, _03928_);
  not (_10442_, _10441_);
  or (_10443_, _10442_, _10438_);
  not (_10444_, _03925_);
  nor (_10445_, _05119_, _03678_);
  and (_10446_, _05119_, _03678_);
  nor (_10447_, _10446_, _10445_);
  nor (_10448_, _05307_, _04139_);
  and (_10449_, _05307_, _04139_);
  nor (_10450_, _10449_, _10448_);
  and (_10451_, _10450_, _10447_);
  and (_10452_, _04700_, _03715_);
  not (_10453_, _10452_);
  and (_10454_, _04900_, _04563_);
  nor (_10455_, _04900_, _04563_);
  nor (_10456_, _10455_, _10454_);
  and (_10457_, _10456_, _10453_);
  and (_10458_, _10457_, _10451_);
  nor (_10459_, _04700_, _03715_);
  not (_10460_, _10459_);
  nor (_10461_, _05568_, _05421_);
  nor (_10462_, _10461_, _05569_);
  and (_10463_, _06065_, _03810_);
  nor (_10464_, _06065_, _03810_);
  nor (_10465_, _10464_, _10463_);
  and (_10466_, _10465_, _10462_);
  nor (_10467_, _05857_, _04093_);
  and (_10468_, _05857_, _04093_);
  nor (_10469_, _10468_, _10467_);
  nor (_10470_, _05950_, _04526_);
  and (_10471_, _05950_, _04526_);
  nor (_10472_, _10471_, _10470_);
  and (_10473_, _10472_, _10469_);
  and (_10474_, _10473_, _10466_);
  and (_10475_, _10474_, _10460_);
  and (_10476_, _10475_, _10458_);
  or (_10477_, _10476_, _10218_);
  nand (_10478_, _10476_, _10212_);
  and (_10479_, _10478_, _10477_);
  or (_10480_, _10479_, _10441_);
  and (_10481_, _10480_, _10444_);
  and (_10482_, _10481_, _10443_);
  or (_10483_, _10482_, _03868_);
  or (_10484_, _10483_, _10254_);
  and (_10485_, _03751_, _03423_);
  nor (_10486_, _10485_, _03920_);
  not (_10487_, _08752_);
  and (_10488_, _05716_, _03498_);
  or (_10489_, _10488_, _08753_);
  and (_10490_, _10489_, _10487_);
  nor (_10491_, _08744_, _08742_);
  nor (_10492_, _10491_, _08748_);
  nor (_10493_, _08738_, _08737_);
  nor (_10494_, _10493_, _08741_);
  nor (_10495_, _08736_, _06557_);
  and (_10496_, _10495_, _10494_);
  and (_10497_, _10496_, _10492_);
  and (_10498_, _10497_, _10490_);
  and (_10499_, _10498_, _06993_);
  not (_10500_, _10498_);
  and (_10501_, _10500_, _10218_);
  or (_10502_, _10501_, _03918_);
  or (_10503_, _10502_, _10499_);
  and (_10504_, _10503_, _10486_);
  and (_10505_, _10504_, _10484_);
  and (_10506_, _03715_, _03498_);
  nor (_10507_, _10506_, _08793_);
  nor (_10508_, _10507_, _08792_);
  nor (_10509_, _08784_, _08785_);
  nor (_10510_, _10509_, _08788_);
  nor (_10511_, _08779_, _08783_);
  nor (_10512_, _08776_, _08537_);
  and (_10513_, _10512_, _10511_);
  and (_10514_, _10513_, _10510_);
  and (_10515_, _10514_, _10508_);
  or (_10516_, _10515_, _10218_);
  nand (_10517_, _10515_, _10212_);
  and (_10518_, _10517_, _03920_);
  and (_10519_, _10518_, _10516_);
  nand (_10520_, _10485_, _10054_);
  nor (_10521_, _04939_, _05049_);
  and (_10522_, _10521_, _03844_);
  and (_10523_, _10522_, _03840_);
  nand (_10524_, _10523_, _10520_);
  or (_10525_, _10524_, _10519_);
  or (_10526_, _10525_, _10505_);
  or (_10527_, _10523_, _07003_);
  and (_10528_, _10527_, _10092_);
  and (_10529_, _10528_, _10526_);
  or (_10530_, _10529_, _10094_);
  and (_10531_, _03880_, _03441_);
  and (_10532_, _10531_, _10530_);
  or (_10533_, _10531_, _10422_);
  nand (_10534_, _10533_, _10087_);
  or (_10535_, _10534_, _10532_);
  and (_10536_, _10535_, _10088_);
  or (_10537_, _10536_, _10086_);
  or (_10538_, _10085_, _07003_);
  and (_10539_, _10538_, _03426_);
  and (_10540_, _10539_, _10537_);
  and (_10541_, _10054_, _03425_);
  nor (_10542_, _03746_, _03456_);
  not (_10543_, _10542_);
  or (_10544_, _10543_, _10541_);
  or (_10545_, _10544_, _10540_);
  or (_10546_, _10542_, _07003_);
  and (_10547_, _10546_, _09861_);
  and (_10548_, _10547_, _10545_);
  nand (_10549_, _06993_, _03921_);
  nand (_10550_, _10549_, _07926_);
  or (_10551_, _10550_, _10548_);
  or (_10552_, _07926_, _07003_);
  and (_10553_, _10552_, _03820_);
  and (_10554_, _10553_, _10551_);
  or (_10555_, _10554_, _10084_);
  nor (_10556_, _07010_, _03469_);
  and (_10557_, _10556_, _10555_);
  not (_10558_, _10556_);
  and (_10559_, _10558_, _10054_);
  nor (_10560_, _03816_, _03398_);
  not (_10561_, _10560_);
  or (_10562_, _10561_, _10559_);
  or (_10563_, _10562_, _10557_);
  and (_10564_, _03397_, _03373_);
  not (_10565_, _10564_);
  or (_10566_, _10560_, _07003_);
  and (_10567_, _10566_, _10565_);
  and (_10568_, _10567_, _10563_);
  and (_10569_, _10564_, _10377_);
  or (_10570_, _10569_, _06309_);
  or (_10571_, _10570_, _10568_);
  or (_10572_, _07003_, _06138_);
  and (_10573_, _10572_, _10571_);
  or (_10574_, _10573_, _03903_);
  or (_10575_, _06993_, _04778_);
  and (_10576_, _10575_, _08493_);
  and (_10577_, _10576_, _10574_);
  and (_10578_, _08492_, _07003_);
  or (_10579_, _10578_, _10577_);
  and (_10580_, _03423_, _03400_);
  not (_10581_, _10580_);
  and (_10582_, _10581_, _10579_);
  nor (_10583_, _03815_, _03401_);
  not (_10584_, _10583_);
  not (_10585_, \oc8051_golden_model_1.DPH [0]);
  and (_10586_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_10587_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_10588_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_10589_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_10590_, _10589_, _10588_);
  and (_10591_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_10592_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  and (_10593_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_10594_, _03569_, _03565_);
  not (_10595_, _10594_);
  nor (_10596_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_10597_, _10596_, _10593_);
  and (_10598_, _10597_, _10595_);
  nor (_10599_, _10598_, _10593_);
  nor (_10600_, _10599_, _10592_);
  nor (_10601_, _10600_, _10591_);
  not (_10602_, _10601_);
  and (_10603_, _10602_, _10590_);
  nor (_10604_, _10603_, _10588_);
  nor (_10605_, _10604_, _10587_);
  nor (_10606_, _10605_, _10586_);
  nor (_10607_, _10606_, _10585_);
  and (_10608_, _10607_, \oc8051_golden_model_1.DPH [1]);
  and (_10609_, _10608_, \oc8051_golden_model_1.DPH [2]);
  and (_10610_, _10609_, \oc8051_golden_model_1.DPH [3]);
  and (_10611_, _10610_, \oc8051_golden_model_1.DPH [4]);
  and (_10612_, _10611_, \oc8051_golden_model_1.DPH [5]);
  and (_10613_, _10612_, \oc8051_golden_model_1.DPH [6]);
  nand (_10614_, _10613_, \oc8051_golden_model_1.DPH [7]);
  or (_10615_, _10613_, \oc8051_golden_model_1.DPH [7]);
  and (_10616_, _10615_, _10580_);
  and (_10617_, _10616_, _10614_);
  or (_10618_, _10617_, _10584_);
  or (_10619_, _10618_, _10582_);
  and (_10620_, _03400_, _03373_);
  not (_10621_, _10620_);
  or (_10622_, _10583_, _07003_);
  and (_10623_, _10622_, _10621_);
  and (_10624_, _10623_, _10619_);
  not (_10625_, _10082_);
  or (_10626_, _10377_, _08826_);
  not (_10627_, _08826_);
  or (_10628_, _10627_, _07003_);
  and (_10629_, _10628_, _10620_);
  and (_10630_, _10629_, _10626_);
  or (_10631_, _10630_, _10625_);
  or (_10632_, _10631_, _10624_);
  and (_10633_, _10632_, _10083_);
  or (_10634_, _10633_, _10080_);
  or (_10635_, _10079_, _07003_);
  and (_10636_, _10635_, _04790_);
  and (_10637_, _10636_, _10634_);
  nand (_10638_, _06993_, _03897_);
  nor (_10639_, _04018_, _03405_);
  nand (_10640_, _10639_, _10638_);
  or (_10642_, _10640_, _10637_);
  and (_10643_, _03404_, _03373_);
  not (_10644_, _10643_);
  or (_10645_, _10639_, _07003_);
  and (_10646_, _10645_, _10644_);
  and (_10647_, _10646_, _10642_);
  or (_10648_, _10377_, _10627_);
  or (_10649_, _08826_, _07003_);
  and (_10650_, _10649_, _10643_);
  and (_10651_, _10650_, _10648_);
  or (_10653_, _10651_, _10647_);
  nor (_10654_, _08547_, _08122_);
  and (_10655_, _10654_, _10653_);
  not (_10656_, _10654_);
  and (_10657_, _10656_, _10054_);
  nor (_10658_, _08553_, _04025_);
  not (_10659_, _10658_);
  or (_10660_, _10659_, _10657_);
  or (_10661_, _10660_, _10655_);
  or (_10662_, _10658_, _07003_);
  and (_10664_, _10662_, _03909_);
  and (_10665_, _10664_, _10661_);
  nand (_10666_, _06993_, _03908_);
  nand (_10667_, _10666_, _10076_);
  or (_10668_, _10667_, _10665_);
  and (_10669_, _10668_, _10078_);
  not (_10670_, _10072_);
  or (_10671_, _10377_, \oc8051_golden_model_1.PSW [7]);
  or (_10672_, _07003_, _08297_);
  and (_10673_, _10672_, _10074_);
  and (_10675_, _10673_, _10671_);
  or (_10676_, _10675_, _10670_);
  or (_10677_, _10676_, _10669_);
  and (_10678_, _10677_, _10073_);
  or (_10679_, _10678_, _08582_);
  or (_10680_, _08581_, _07003_);
  and (_10681_, _10680_, _06567_);
  and (_10682_, _10681_, _10679_);
  nand (_10683_, _06993_, _03914_);
  nand (_10684_, _10683_, _10065_);
  or (_10686_, _10684_, _10682_);
  and (_10687_, _10686_, _10067_);
  not (_10688_, _10061_);
  or (_10689_, _10377_, _08297_);
  or (_10690_, _07003_, \oc8051_golden_model_1.PSW [7]);
  and (_10691_, _10690_, _10063_);
  and (_10692_, _10691_, _10689_);
  or (_10693_, _10692_, _10688_);
  or (_10694_, _10693_, _10687_);
  and (_10695_, _10694_, _10062_);
  or (_10697_, _10695_, _08629_);
  or (_10698_, _08628_, _07003_);
  and (_10699_, _10698_, _08658_);
  and (_10700_, _10699_, _10697_);
  and (_10701_, _10054_, _08657_);
  or (_10702_, _10701_, _04034_);
  or (_10703_, _10702_, _10700_);
  not (_10704_, _04034_);
  or (_10705_, _05568_, _10704_);
  and (_10706_, _10705_, _10703_);
  or (_10708_, _10706_, _03383_);
  or (_10709_, _07003_, _03384_);
  and (_10710_, _10709_, _04097_);
  and (_10711_, _10710_, _10708_);
  not (_10712_, _10059_);
  not (_10713_, _05763_);
  and (_10714_, _06085_, \oc8051_golden_model_1.TCON [2]);
  and (_10715_, _06096_, \oc8051_golden_model_1.ACC [2]);
  nor (_10716_, _10715_, _10714_);
  and (_10717_, _06091_, \oc8051_golden_model_1.IP [2]);
  not (_10718_, _10717_);
  and (_10719_, _06094_, \oc8051_golden_model_1.PSW [2]);
  and (_10720_, _06088_, \oc8051_golden_model_1.B [2]);
  nor (_10721_, _10720_, _10719_);
  and (_10722_, _10721_, _10718_);
  and (_10723_, _10722_, _10716_);
  and (_10724_, _06101_, \oc8051_golden_model_1.SCON [2]);
  and (_10725_, _06103_, \oc8051_golden_model_1.IE [2]);
  nor (_10726_, _10725_, _10724_);
  and (_10727_, _06106_, \oc8051_golden_model_1.P2INREG [2]);
  and (_10728_, _06108_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_10729_, _10728_, _10727_);
  and (_10730_, _06112_, \oc8051_golden_model_1.P0INREG [2]);
  and (_10731_, _06114_, \oc8051_golden_model_1.P1INREG [2]);
  nor (_10732_, _10731_, _10730_);
  and (_10733_, _10732_, _10729_);
  and (_10734_, _10733_, _10726_);
  and (_10735_, _10734_, _10723_);
  and (_10736_, _10735_, _10713_);
  and (_10737_, _05477_, _04139_);
  not (_10738_, _10737_);
  nor (_10739_, _10738_, _10736_);
  and (_10740_, _05467_, _04139_);
  not (_10741_, _10740_);
  not (_10742_, _05668_);
  and (_10743_, _06085_, \oc8051_golden_model_1.TCON [1]);
  and (_10744_, _06096_, \oc8051_golden_model_1.ACC [1]);
  nor (_10745_, _10744_, _10743_);
  and (_10746_, _06091_, \oc8051_golden_model_1.IP [1]);
  not (_10747_, _10746_);
  and (_10748_, _06094_, \oc8051_golden_model_1.PSW [1]);
  and (_10749_, _06088_, \oc8051_golden_model_1.B [1]);
  nor (_10750_, _10749_, _10748_);
  and (_10751_, _10750_, _10747_);
  and (_10752_, _10751_, _10745_);
  and (_10753_, _06101_, \oc8051_golden_model_1.SCON [1]);
  and (_10754_, _06103_, \oc8051_golden_model_1.IE [1]);
  nor (_10755_, _10754_, _10753_);
  and (_10756_, _06106_, \oc8051_golden_model_1.P2INREG [1]);
  and (_10757_, _06108_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_10758_, _10757_, _10756_);
  and (_10759_, _06112_, \oc8051_golden_model_1.P0INREG [1]);
  and (_10760_, _06114_, \oc8051_golden_model_1.P1INREG [1]);
  nor (_10761_, _10760_, _10759_);
  and (_10762_, _10761_, _10758_);
  and (_10763_, _10762_, _10755_);
  and (_10764_, _10763_, _10752_);
  and (_10765_, _10764_, _10742_);
  nor (_10766_, _10765_, _10741_);
  nor (_10767_, _10766_, _10739_);
  not (_10768_, _05952_);
  and (_10769_, _06091_, \oc8051_golden_model_1.IP [4]);
  and (_10770_, _06088_, \oc8051_golden_model_1.B [4]);
  nor (_10771_, _10770_, _10769_);
  and (_10772_, _06094_, \oc8051_golden_model_1.PSW [4]);
  and (_10773_, _06096_, \oc8051_golden_model_1.ACC [4]);
  nor (_10774_, _10773_, _10772_);
  and (_10775_, _10774_, _10771_);
  and (_10776_, _06085_, \oc8051_golden_model_1.TCON [4]);
  and (_10777_, _06108_, \oc8051_golden_model_1.P3INREG [4]);
  and (_10778_, _06106_, \oc8051_golden_model_1.P2INREG [4]);
  or (_10779_, _10778_, _10777_);
  nor (_10780_, _10779_, _10776_);
  and (_10781_, _06101_, \oc8051_golden_model_1.SCON [4]);
  and (_10782_, _06103_, \oc8051_golden_model_1.IE [4]);
  nor (_10783_, _10782_, _10781_);
  and (_10784_, _06112_, \oc8051_golden_model_1.P0INREG [4]);
  and (_10785_, _06114_, \oc8051_golden_model_1.P1INREG [4]);
  nor (_10786_, _10785_, _10784_);
  and (_10787_, _10786_, _10783_);
  and (_10788_, _10787_, _10780_);
  and (_10789_, _10788_, _10775_);
  and (_10790_, _10789_, _10768_);
  and (_10791_, _05417_, _05243_);
  not (_10792_, _10791_);
  nor (_10793_, _10792_, _10790_);
  nor (_10794_, _10793_, _06146_);
  and (_10795_, _10794_, _10767_);
  not (_10796_, _05432_);
  not (_10797_, _05715_);
  and (_10798_, _06085_, \oc8051_golden_model_1.TCON [0]);
  and (_10799_, _06096_, \oc8051_golden_model_1.ACC [0]);
  nor (_10800_, _10799_, _10798_);
  and (_10801_, _06091_, \oc8051_golden_model_1.IP [0]);
  not (_10802_, _10801_);
  and (_10803_, _06094_, \oc8051_golden_model_1.PSW [0]);
  and (_10804_, _06088_, \oc8051_golden_model_1.B [0]);
  nor (_10805_, _10804_, _10803_);
  and (_10806_, _10805_, _10802_);
  and (_10807_, _10806_, _10800_);
  and (_10808_, _06101_, \oc8051_golden_model_1.SCON [0]);
  and (_10809_, _06103_, \oc8051_golden_model_1.IE [0]);
  nor (_10810_, _10809_, _10808_);
  and (_10811_, _06106_, \oc8051_golden_model_1.P2INREG [0]);
  and (_10812_, _06108_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_10813_, _10812_, _10811_);
  and (_10814_, _06112_, \oc8051_golden_model_1.P0INREG [0]);
  and (_10815_, _06114_, \oc8051_golden_model_1.P1INREG [0]);
  nor (_10816_, _10815_, _10814_);
  and (_10817_, _10816_, _10813_);
  and (_10818_, _10817_, _10810_);
  and (_10819_, _10818_, _10807_);
  and (_10820_, _10819_, _10797_);
  nor (_10821_, _10820_, _10796_);
  not (_10822_, _06067_);
  and (_10823_, _06085_, \oc8051_golden_model_1.TCON [6]);
  and (_10824_, _06088_, \oc8051_golden_model_1.B [6]);
  nor (_10825_, _10824_, _10823_);
  and (_10826_, _06091_, \oc8051_golden_model_1.IP [6]);
  not (_10827_, _10826_);
  and (_10828_, _06094_, \oc8051_golden_model_1.PSW [6]);
  and (_10829_, _06096_, \oc8051_golden_model_1.ACC [6]);
  nor (_10830_, _10829_, _10828_);
  and (_10831_, _10830_, _10827_);
  and (_10832_, _10831_, _10825_);
  and (_10833_, _06101_, \oc8051_golden_model_1.SCON [6]);
  and (_10834_, _06103_, \oc8051_golden_model_1.IE [6]);
  nor (_10835_, _10834_, _10833_);
  and (_10836_, _06106_, \oc8051_golden_model_1.P2INREG [6]);
  and (_10837_, _06108_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_10838_, _10837_, _10836_);
  and (_10839_, _06112_, \oc8051_golden_model_1.P0INREG [6]);
  and (_10840_, _06114_, \oc8051_golden_model_1.P1INREG [6]);
  nor (_10841_, _10840_, _10839_);
  and (_10842_, _10841_, _10838_);
  and (_10843_, _10842_, _10835_);
  and (_10844_, _10843_, _10832_);
  and (_10845_, _10844_, _10822_);
  and (_10846_, _05477_, _05243_);
  not (_10847_, _10846_);
  nor (_10848_, _10847_, _10845_);
  nor (_10849_, _10848_, _10821_);
  not (_10850_, _05620_);
  and (_10851_, _06085_, \oc8051_golden_model_1.TCON [3]);
  and (_10852_, _06096_, \oc8051_golden_model_1.ACC [3]);
  nor (_10853_, _10852_, _10851_);
  and (_10854_, _06091_, \oc8051_golden_model_1.IP [3]);
  not (_10855_, _10854_);
  and (_10856_, _06094_, \oc8051_golden_model_1.PSW [3]);
  and (_10857_, _06088_, \oc8051_golden_model_1.B [3]);
  nor (_10858_, _10857_, _10856_);
  and (_10859_, _10858_, _10855_);
  and (_10860_, _10859_, _10853_);
  and (_10861_, _06101_, \oc8051_golden_model_1.SCON [3]);
  and (_10862_, _06103_, \oc8051_golden_model_1.IE [3]);
  nor (_10863_, _10862_, _10861_);
  and (_10864_, _06106_, \oc8051_golden_model_1.P2INREG [3]);
  and (_10865_, _06108_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_10866_, _10865_, _10864_);
  and (_10867_, _06112_, \oc8051_golden_model_1.P0INREG [3]);
  and (_10868_, _06114_, \oc8051_golden_model_1.P1INREG [3]);
  nor (_10869_, _10868_, _10867_);
  and (_10870_, _10869_, _10866_);
  and (_10871_, _10870_, _10863_);
  and (_10872_, _10871_, _10860_);
  and (_10873_, _10872_, _10850_);
  and (_10874_, _05457_, _04139_);
  not (_10875_, _10874_);
  nor (_10876_, _10875_, _10873_);
  not (_10877_, _05858_);
  and (_10878_, _06085_, \oc8051_golden_model_1.TCON [5]);
  and (_10879_, _06088_, \oc8051_golden_model_1.B [5]);
  nor (_10880_, _10879_, _10878_);
  and (_10881_, _06094_, \oc8051_golden_model_1.PSW [5]);
  not (_10882_, _10881_);
  and (_10883_, _06091_, \oc8051_golden_model_1.IP [5]);
  and (_10884_, _06096_, \oc8051_golden_model_1.ACC [5]);
  nor (_10885_, _10884_, _10883_);
  and (_10886_, _10885_, _10882_);
  and (_10887_, _10886_, _10880_);
  and (_10888_, _06101_, \oc8051_golden_model_1.SCON [5]);
  and (_10889_, _06103_, \oc8051_golden_model_1.IE [5]);
  nor (_10890_, _10889_, _10888_);
  and (_10891_, _06106_, \oc8051_golden_model_1.P2INREG [5]);
  and (_10892_, _06108_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_10893_, _10892_, _10891_);
  and (_10894_, _06112_, \oc8051_golden_model_1.P0INREG [5]);
  and (_10895_, _06114_, \oc8051_golden_model_1.P1INREG [5]);
  nor (_10896_, _10895_, _10894_);
  and (_10897_, _10896_, _10893_);
  and (_10898_, _10897_, _10890_);
  and (_10899_, _10898_, _10887_);
  and (_10900_, _10899_, _10877_);
  and (_10901_, _05467_, _05243_);
  not (_10902_, _10901_);
  nor (_10903_, _10902_, _10900_);
  nor (_10904_, _10903_, _10876_);
  and (_10905_, _10904_, _10849_);
  and (_10906_, _10905_, _10795_);
  not (_10907_, _10906_);
  or (_10908_, _10218_, _10907_);
  or (_10909_, _06993_, _10906_);
  and (_10910_, _10909_, _03913_);
  and (_10911_, _10910_, _10908_);
  or (_10912_, _10911_, _10712_);
  or (_10913_, _10912_, _10711_);
  and (_10914_, _10913_, _10060_);
  or (_10915_, _10914_, _10057_);
  or (_10916_, _10056_, _07003_);
  and (_10917_, _10916_, _08773_);
  and (_10918_, _10917_, _10915_);
  and (_10919_, _10054_, _08772_);
  or (_10920_, _10919_, _03777_);
  or (_10921_, _10920_, _10918_);
  or (_10922_, _05568_, _03778_);
  and (_10923_, _10922_, _10921_);
  or (_10924_, _10923_, _03410_);
  or (_10925_, _07003_, _03411_);
  and (_10926_, _10925_, _03776_);
  and (_10927_, _10926_, _10924_);
  or (_10928_, _10218_, _10906_);
  nand (_10929_, _10212_, _10906_);
  and (_10930_, _10929_, _10928_);
  and (_10931_, _10930_, _03775_);
  not (_10932_, _03244_);
  nor (_10933_, _07919_, _10932_);
  and (_10934_, _07922_, _03244_);
  nor (_10935_, _10934_, _10933_);
  and (_10936_, _10935_, _04813_);
  not (_10937_, _10936_);
  or (_10938_, _10937_, _10931_);
  or (_10939_, _10938_, _10927_);
  or (_10940_, _10936_, _10054_);
  and (_10941_, _10940_, _03774_);
  and (_10942_, _10941_, _10939_);
  nor (_10943_, _08820_, _08815_);
  nand (_10944_, _07003_, _03773_);
  nand (_10945_, _10944_, _10943_);
  or (_10946_, _10945_, _10942_);
  or (_10947_, _10054_, _10943_);
  and (_10948_, _10947_, _03900_);
  and (_10949_, _10948_, _10946_);
  and (_10950_, _03899_, _03647_);
  or (_10951_, _10950_, _03414_);
  or (_10952_, _10951_, _10949_);
  not (_10953_, _03414_);
  or (_10954_, _07003_, _10953_);
  and (_10955_, _10954_, _03375_);
  and (_10956_, _10955_, _10952_);
  and (_10957_, _10930_, _03374_);
  and (_10958_, _04827_, _04482_);
  not (_10959_, _10958_);
  or (_10960_, _10959_, _10957_);
  or (_10961_, _10960_, _10956_);
  or (_10962_, _10958_, _10054_);
  and (_10963_, _10962_, _04060_);
  and (_10964_, _10963_, _10961_);
  nor (_10965_, _08844_, _08837_);
  nand (_10966_, _07003_, _03772_);
  nand (_10967_, _10966_, _10965_);
  or (_10968_, _10967_, _10964_);
  not (_10969_, _03901_);
  or (_10970_, _10054_, _10965_);
  and (_10971_, _10970_, _10969_);
  and (_10972_, _10971_, _10968_);
  and (_10973_, _03901_, _03647_);
  or (_10974_, _10973_, _03413_);
  or (_10975_, _10974_, _10972_);
  not (_10976_, _10042_);
  not (_10977_, _03413_);
  or (_10978_, _07003_, _10977_);
  and (_10979_, _10978_, _10976_);
  and (_10980_, _10979_, _10975_);
  or (_10981_, _10980_, _10055_);
  or (_10982_, _10981_, _43156_);
  or (_10983_, _43152_, \oc8051_golden_model_1.PC [15]);
  and (_10984_, _10983_, _41894_);
  and (_40698_, _10984_, _10982_);
  not (_10985_, \oc8051_golden_model_1.P2 [7]);
  nor (_10986_, _05498_, _10985_);
  and (_10987_, _05498_, \oc8051_golden_model_1.P2 [7]);
  and (_10988_, _05500_, \oc8051_golden_model_1.P3 [7]);
  nor (_10989_, _10988_, _10987_);
  and (_10990_, _05505_, \oc8051_golden_model_1.P0 [7]);
  and (_10991_, _05455_, \oc8051_golden_model_1.P1 [7]);
  nor (_10992_, _10991_, _10990_);
  and (_10993_, _10992_, _10989_);
  not (_10994_, _05452_);
  and (_10995_, _05482_, _10994_);
  nor (_10996_, _05462_, _05448_);
  and (_10997_, _10996_, _10995_);
  and (_10998_, _10997_, _10993_);
  and (_10999_, _05471_, _05497_);
  and (_11000_, _10999_, _05519_);
  and (_11001_, _11000_, _10998_);
  and (_11002_, _11001_, _05443_);
  and (_11003_, _11002_, _06079_);
  nand (_11004_, _11003_, _06554_);
  or (_11005_, _11003_, _06554_);
  and (_11006_, _11005_, _11004_);
  and (_11007_, _11006_, _05498_);
  or (_11008_, _11007_, _10986_);
  and (_11009_, _11008_, _04018_);
  and (_11010_, _06348_, _05498_);
  or (_11011_, _11010_, _10986_);
  or (_11012_, _11011_, _04778_);
  nor (_11013_, _06106_, _10985_);
  and (_11014_, _06112_, \oc8051_golden_model_1.P0 [7]);
  and (_11015_, _06106_, \oc8051_golden_model_1.P2 [7]);
  nor (_11016_, _11015_, _11014_);
  and (_11017_, _06114_, \oc8051_golden_model_1.P1 [7]);
  and (_11018_, _06108_, \oc8051_golden_model_1.P3 [7]);
  nor (_11019_, _11018_, _11017_);
  and (_11020_, _11019_, _11016_);
  and (_11021_, _11020_, _06105_);
  and (_11022_, _11021_, _06100_);
  and (_11023_, _11022_, _06079_);
  nor (_11024_, _11023_, _05486_);
  and (_11025_, _11024_, _06106_);
  or (_11026_, _11025_, _11013_);
  and (_11027_, _11026_, _03759_);
  not (_11028_, _11003_);
  nor (_11029_, _05976_, _05971_);
  nand (_11030_, _11029_, _05987_);
  nor (_11031_, _11030_, _05970_);
  and (_11032_, _05498_, \oc8051_golden_model_1.P2 [6]);
  and (_11033_, _05500_, \oc8051_golden_model_1.P3 [6]);
  nor (_11034_, _11033_, _11032_);
  and (_11035_, _05505_, \oc8051_golden_model_1.P0 [6]);
  and (_11036_, _05455_, \oc8051_golden_model_1.P1 [6]);
  nor (_11037_, _11036_, _11035_);
  and (_11038_, _11037_, _11034_);
  and (_11039_, _11038_, _05968_);
  and (_11040_, _05983_, _05996_);
  and (_11041_, _11040_, _11039_);
  and (_11042_, _11041_, _06008_);
  and (_11043_, _11042_, _11031_);
  and (_11044_, _11043_, _10822_);
  and (_11045_, _05498_, \oc8051_golden_model_1.P2 [5]);
  and (_11046_, _05500_, \oc8051_golden_model_1.P3 [5]);
  nor (_11047_, _11046_, _11045_);
  and (_11048_, _05505_, \oc8051_golden_model_1.P0 [5]);
  and (_11049_, _05455_, \oc8051_golden_model_1.P1 [5]);
  nor (_11050_, _11049_, _11048_);
  and (_11051_, _11050_, _11047_);
  and (_11052_, _11051_, _05774_);
  and (_11053_, _05784_, _05796_);
  nor (_11054_, _05779_, _05776_);
  nand (_11055_, _11054_, _05787_);
  nor (_11056_, _11055_, _05775_);
  and (_11057_, _11056_, _05808_);
  and (_11058_, _11057_, _11053_);
  and (_11059_, _11058_, _11052_);
  and (_11060_, _11059_, _10877_);
  nor (_11061_, _05871_, _05868_);
  nand (_11062_, _11061_, _05879_);
  nor (_11063_, _11062_, _05867_);
  and (_11064_, _05498_, \oc8051_golden_model_1.P2 [4]);
  and (_11065_, _05500_, \oc8051_golden_model_1.P3 [4]);
  nor (_11066_, _11065_, _11064_);
  and (_11067_, _05505_, \oc8051_golden_model_1.P0 [4]);
  and (_11068_, _05455_, \oc8051_golden_model_1.P1 [4]);
  nor (_11069_, _11068_, _11067_);
  and (_11070_, _11069_, _11066_);
  and (_11071_, _11070_, _05866_);
  and (_11072_, _05876_, _05888_);
  and (_11073_, _11072_, _11071_);
  and (_11074_, _11073_, _05900_);
  and (_11075_, _11074_, _11063_);
  and (_11076_, _11075_, _10768_);
  and (_11077_, _05498_, \oc8051_golden_model_1.P2 [3]);
  and (_11078_, _05500_, \oc8051_golden_model_1.P3 [3]);
  nor (_11079_, _11078_, _11077_);
  and (_11080_, _05505_, \oc8051_golden_model_1.P0 [3]);
  and (_11081_, _05455_, \oc8051_golden_model_1.P1 [3]);
  nor (_11082_, _11081_, _11080_);
  and (_11083_, _11082_, _11079_);
  and (_11084_, _11083_, _05606_);
  and (_11085_, _11084_, _05599_);
  and (_11086_, _11085_, _05593_);
  and (_11087_, _11086_, _10850_);
  and (_11088_, _05498_, \oc8051_golden_model_1.P2 [2]);
  and (_11089_, _05500_, \oc8051_golden_model_1.P3 [2]);
  nor (_11090_, _11089_, _11088_);
  and (_11091_, _05505_, \oc8051_golden_model_1.P0 [2]);
  and (_11092_, _05455_, \oc8051_golden_model_1.P1 [2]);
  nor (_11093_, _11092_, _11091_);
  and (_11094_, _11093_, _11090_);
  and (_11095_, _11094_, _05724_);
  and (_11096_, _05734_, _05746_);
  nor (_11097_, _05729_, _05726_);
  nand (_11098_, _11097_, _05737_);
  nor (_11099_, _11098_, _05725_);
  and (_11100_, _11099_, _05758_);
  and (_11101_, _11100_, _11096_);
  and (_11102_, _11101_, _11095_);
  and (_11103_, _11102_, _10713_);
  and (_11104_, _05505_, \oc8051_golden_model_1.P0 [1]);
  and (_11105_, _05455_, \oc8051_golden_model_1.P1 [1]);
  nor (_11106_, _11105_, _11104_);
  and (_11107_, _05498_, \oc8051_golden_model_1.P2 [1]);
  and (_11108_, _05500_, \oc8051_golden_model_1.P3 [1]);
  nor (_11109_, _11108_, _11107_);
  and (_11110_, _11109_, _05655_);
  and (_11111_, _11110_, _11106_);
  and (_11112_, _11111_, _05653_);
  and (_11113_, _11112_, _05646_);
  and (_11114_, _11113_, _05640_);
  and (_11115_, _11114_, _10742_);
  and (_11116_, _05498_, \oc8051_golden_model_1.P2 [0]);
  and (_11117_, _05500_, \oc8051_golden_model_1.P3 [0]);
  nor (_11118_, _11117_, _11116_);
  and (_11119_, _05505_, \oc8051_golden_model_1.P0 [0]);
  and (_11120_, _05455_, \oc8051_golden_model_1.P1 [0]);
  nor (_11121_, _11120_, _11119_);
  and (_11122_, _11121_, _11118_);
  and (_11123_, _11122_, _05701_);
  and (_11124_, _11123_, _05694_);
  and (_11125_, _11124_, _05688_);
  and (_11126_, _11125_, _10797_);
  and (_11127_, _11126_, _11115_);
  and (_11128_, _11127_, _11103_);
  and (_11129_, _11128_, _11087_);
  and (_11130_, _11129_, _11076_);
  and (_11131_, _11130_, _11060_);
  and (_11132_, _11131_, _11044_);
  or (_11133_, _11132_, _11028_);
  nand (_11134_, _11132_, _11028_);
  and (_11135_, _11134_, _11133_);
  and (_11136_, _11135_, _05498_);
  or (_11137_, _11136_, _10986_);
  or (_11138_, _11137_, _04722_);
  and (_11139_, _05498_, \oc8051_golden_model_1.ACC [7]);
  or (_11140_, _11139_, _10986_);
  and (_11141_, _11140_, _04707_);
  nor (_11142_, _04707_, _10985_);
  or (_11143_, _11142_, _03850_);
  or (_11144_, _11143_, _11141_);
  and (_11145_, _11144_, _03764_);
  and (_11146_, _11145_, _11138_);
  nand (_11147_, _11023_, _06145_);
  and (_11148_, _11147_, _06106_);
  or (_11149_, _11148_, _11013_);
  and (_11150_, _11149_, _03763_);
  or (_11151_, _11150_, _03848_);
  or (_11152_, _11151_, _11146_);
  and (_11153_, _05568_, _05498_);
  or (_11154_, _11153_, _10986_);
  or (_11155_, _11154_, _04733_);
  and (_11156_, _11155_, _11152_);
  or (_11157_, _11156_, _03854_);
  or (_11158_, _11140_, _03855_);
  and (_11159_, _11158_, _03760_);
  and (_11160_, _11159_, _11157_);
  or (_11161_, _11160_, _11027_);
  and (_11162_, _11161_, _03753_);
  or (_11163_, _11023_, _06145_);
  or (_11164_, _11163_, _11013_);
  and (_11165_, _11149_, _03752_);
  and (_11166_, _11165_, _11164_);
  or (_11167_, _11166_, _11162_);
  and (_11168_, _11167_, _03747_);
  or (_11169_, _11024_, _06142_);
  and (_11170_, _11169_, _06106_);
  or (_11171_, _11170_, _11013_);
  and (_11172_, _11171_, _03746_);
  or (_11173_, _11172_, _07927_);
  or (_11174_, _11173_, _11168_);
  and (_11175_, _06248_, _05498_);
  or (_11176_, _10986_, _03738_);
  or (_11177_, _11176_, _11175_);
  or (_11178_, _11154_, _07925_);
  and (_11179_, _11178_, _03820_);
  and (_11180_, _11179_, _11177_);
  and (_11181_, _11180_, _11174_);
  and (_11182_, _06505_, \oc8051_golden_model_1.P1 [7]);
  and (_11183_, _06507_, \oc8051_golden_model_1.P3 [7]);
  or (_11184_, _11183_, _11182_);
  or (_11185_, _11184_, _06513_);
  and (_11186_, _06501_, \oc8051_golden_model_1.P0 [7]);
  and (_11187_, _06515_, \oc8051_golden_model_1.P2 [7]);
  or (_11188_, _11187_, _11186_);
  nor (_11189_, _11188_, _11185_);
  and (_11190_, _11189_, _06531_);
  and (_11191_, _11190_, _06500_);
  nand (_11192_, _11191_, _06487_);
  or (_11193_, _11192_, _06343_);
  and (_11194_, _11193_, _05498_);
  or (_11195_, _11194_, _10986_);
  and (_11196_, _11195_, _03455_);
  or (_11197_, _11196_, _03903_);
  or (_11198_, _11197_, _11181_);
  and (_11199_, _11198_, _11012_);
  or (_11200_, _11199_, _03897_);
  nand (_11201_, _11003_, _06342_);
  or (_11202_, _11003_, _06342_);
  and (_11203_, _11202_, _11201_);
  and (_11204_, _11203_, _05498_);
  or (_11205_, _10986_, _04790_);
  or (_11206_, _11205_, _11204_);
  and (_11207_, _11206_, _04792_);
  and (_11208_, _11207_, _11200_);
  or (_11209_, _11208_, _11009_);
  and (_11210_, _11209_, _03909_);
  or (_11211_, _11028_, _10986_);
  and (_11212_, _11011_, _03908_);
  and (_11213_, _11212_, _11211_);
  or (_11214_, _11213_, _11210_);
  and (_11215_, _11214_, _04785_);
  and (_11216_, _11140_, _04027_);
  and (_11217_, _11216_, _11211_);
  or (_11218_, _11217_, _03914_);
  or (_11219_, _11218_, _11215_);
  and (_11220_, _11201_, _05498_);
  or (_11221_, _10986_, _06567_);
  or (_11222_, _11221_, _11220_);
  and (_11223_, _11222_, _06572_);
  and (_11224_, _11223_, _11219_);
  and (_11225_, _11004_, _05498_);
  or (_11226_, _11225_, _10986_);
  and (_11227_, _11226_, _04011_);
  or (_11228_, _11227_, _03773_);
  or (_11229_, _11228_, _11224_);
  or (_11230_, _11137_, _03774_);
  and (_11231_, _11230_, _03375_);
  and (_11232_, _11231_, _11229_);
  and (_11233_, _11026_, _03374_);
  or (_11234_, _11233_, _03772_);
  or (_11235_, _11234_, _11232_);
  not (_11236_, _11044_);
  not (_11237_, _11060_);
  not (_11238_, _11076_);
  not (_11239_, _11087_);
  not (_11240_, _11103_);
  nor (_11241_, _11126_, _11115_);
  and (_11242_, _11241_, _11240_);
  and (_11243_, _11242_, _11239_);
  and (_11244_, _11243_, _11238_);
  and (_11245_, _11244_, _11237_);
  nand (_11246_, _11245_, _11236_);
  nand (_11247_, _11246_, _11003_);
  or (_11248_, _11246_, _11003_);
  and (_11249_, _11248_, _11247_);
  and (_11250_, _11249_, _05498_);
  or (_11251_, _10986_, _04060_);
  or (_11252_, _11251_, _11250_);
  and (_11253_, _11252_, _43152_);
  and (_11254_, _11253_, _11235_);
  nor (_11255_, _43152_, _10985_);
  or (_11256_, _11255_, rst);
  or (_40699_, _11256_, _11254_);
  not (_11257_, _05500_);
  and (_11258_, _11257_, \oc8051_golden_model_1.P3 [7]);
  and (_11259_, _11006_, _05500_);
  or (_11260_, _11259_, _11258_);
  and (_11261_, _11260_, _04018_);
  and (_11262_, _06348_, _05500_);
  or (_11263_, _11262_, _11258_);
  or (_11264_, _11263_, _04778_);
  not (_11265_, _06108_);
  and (_11266_, _11265_, \oc8051_golden_model_1.P3 [7]);
  and (_11267_, _11024_, _06108_);
  or (_11268_, _11267_, _11266_);
  and (_11269_, _11268_, _03759_);
  and (_11270_, _11135_, _05500_);
  or (_11271_, _11270_, _11258_);
  or (_11272_, _11271_, _04722_);
  and (_11273_, _05500_, \oc8051_golden_model_1.ACC [7]);
  or (_11274_, _11273_, _11258_);
  and (_11275_, _11274_, _04707_);
  and (_11276_, _04708_, \oc8051_golden_model_1.P3 [7]);
  or (_11277_, _11276_, _03850_);
  or (_11278_, _11277_, _11275_);
  and (_11279_, _11278_, _03764_);
  and (_11280_, _11279_, _11272_);
  and (_11281_, _11147_, _06108_);
  or (_11282_, _11281_, _11266_);
  and (_11283_, _11282_, _03763_);
  or (_11284_, _11283_, _03848_);
  or (_11285_, _11284_, _11280_);
  and (_11286_, _05568_, _05500_);
  or (_11287_, _11286_, _11258_);
  or (_11288_, _11287_, _04733_);
  and (_11289_, _11288_, _11285_);
  or (_11290_, _11289_, _03854_);
  or (_11291_, _11274_, _03855_);
  and (_11292_, _11291_, _03760_);
  and (_11293_, _11292_, _11290_);
  or (_11294_, _11293_, _11269_);
  and (_11295_, _11294_, _03753_);
  or (_11296_, _11266_, _11163_);
  and (_11297_, _11296_, _03752_);
  and (_11298_, _11297_, _11282_);
  or (_11299_, _11298_, _11295_);
  and (_11300_, _11299_, _03747_);
  and (_11301_, _11169_, _06108_);
  or (_11302_, _11301_, _11266_);
  and (_11303_, _11302_, _03746_);
  or (_11304_, _11303_, _07927_);
  or (_11305_, _11304_, _11300_);
  and (_11306_, _06248_, _05500_);
  or (_11307_, _11258_, _03738_);
  or (_11308_, _11307_, _11306_);
  or (_11309_, _11287_, _07925_);
  and (_11310_, _11309_, _03820_);
  and (_11311_, _11310_, _11308_);
  and (_11312_, _11311_, _11305_);
  and (_11313_, _11193_, _05500_);
  or (_11314_, _11313_, _11258_);
  and (_11315_, _11314_, _03455_);
  or (_11316_, _11315_, _03903_);
  or (_11317_, _11316_, _11312_);
  and (_11318_, _11317_, _11264_);
  or (_11319_, _11318_, _03897_);
  and (_11320_, _11203_, _05500_);
  or (_11321_, _11320_, _11258_);
  or (_11322_, _11321_, _04790_);
  and (_11323_, _11322_, _04792_);
  and (_11324_, _11323_, _11319_);
  or (_11325_, _11324_, _11261_);
  and (_11326_, _11325_, _03909_);
  or (_11327_, _11258_, _11028_);
  and (_11328_, _11263_, _03908_);
  and (_11329_, _11328_, _11327_);
  or (_11330_, _11329_, _11326_);
  and (_11331_, _11330_, _04785_);
  and (_11332_, _11274_, _04027_);
  and (_11333_, _11332_, _11327_);
  or (_11334_, _11333_, _03914_);
  or (_11335_, _11334_, _11331_);
  and (_11336_, _11201_, _05500_);
  or (_11337_, _11258_, _06567_);
  or (_11338_, _11337_, _11336_);
  and (_11339_, _11338_, _06572_);
  and (_11340_, _11339_, _11335_);
  and (_11341_, _11004_, _05500_);
  or (_11342_, _11341_, _11258_);
  and (_11343_, _11342_, _04011_);
  or (_11344_, _11343_, _03773_);
  or (_11345_, _11344_, _11340_);
  or (_11346_, _11271_, _03774_);
  and (_11347_, _11346_, _03375_);
  and (_11348_, _11347_, _11345_);
  and (_11349_, _11268_, _03374_);
  or (_11350_, _11349_, _03772_);
  or (_11351_, _11350_, _11348_);
  and (_11352_, _11249_, _05500_);
  or (_11353_, _11258_, _04060_);
  or (_11354_, _11353_, _11352_);
  and (_11355_, _11354_, _43152_);
  and (_11356_, _11355_, _11351_);
  nor (_11357_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_11358_, _11357_, _05397_);
  or (_40701_, _11358_, _11356_);
  not (_11359_, _05505_);
  and (_11360_, _11359_, \oc8051_golden_model_1.P0 [7]);
  and (_11361_, _11006_, _05505_);
  or (_11362_, _11361_, _11360_);
  and (_11363_, _11362_, _04018_);
  and (_11364_, _06348_, _05505_);
  or (_11365_, _11364_, _11360_);
  or (_11366_, _11365_, _04778_);
  not (_11367_, _06112_);
  and (_11368_, _11367_, \oc8051_golden_model_1.P0 [7]);
  and (_11369_, _11024_, _06112_);
  or (_11370_, _11369_, _11368_);
  and (_11371_, _11370_, _03759_);
  and (_11372_, _11135_, _05505_);
  or (_11373_, _11372_, _11360_);
  or (_11374_, _11373_, _04722_);
  and (_11375_, _05505_, \oc8051_golden_model_1.ACC [7]);
  or (_11376_, _11375_, _11360_);
  and (_11377_, _11376_, _04707_);
  and (_11378_, _04708_, \oc8051_golden_model_1.P0 [7]);
  or (_11379_, _11378_, _03850_);
  or (_11380_, _11379_, _11377_);
  and (_11381_, _11380_, _03764_);
  and (_11382_, _11381_, _11374_);
  and (_11383_, _11147_, _06112_);
  or (_11384_, _11383_, _11368_);
  and (_11385_, _11384_, _03763_);
  or (_11386_, _11385_, _03848_);
  or (_11387_, _11386_, _11382_);
  and (_11388_, _05568_, _05505_);
  or (_11389_, _11388_, _11360_);
  or (_11390_, _11389_, _04733_);
  and (_11391_, _11390_, _11387_);
  or (_11392_, _11391_, _03854_);
  or (_11393_, _11376_, _03855_);
  and (_11394_, _11393_, _03760_);
  and (_11395_, _11394_, _11392_);
  or (_11396_, _11395_, _11371_);
  and (_11397_, _11396_, _03753_);
  or (_11398_, _11368_, _11163_);
  and (_11399_, _11398_, _03752_);
  and (_11400_, _11399_, _11384_);
  or (_11401_, _11400_, _11397_);
  and (_11402_, _11401_, _03747_);
  and (_11403_, _11169_, _06112_);
  or (_11404_, _11403_, _11368_);
  and (_11405_, _11404_, _03746_);
  or (_11406_, _11405_, _07927_);
  or (_11407_, _11406_, _11402_);
  and (_11408_, _06248_, _05505_);
  or (_11409_, _11360_, _03738_);
  or (_11410_, _11409_, _11408_);
  or (_11411_, _11389_, _07925_);
  and (_11412_, _11411_, _03820_);
  and (_11413_, _11412_, _11410_);
  and (_11414_, _11413_, _11407_);
  and (_11415_, _11193_, _05505_);
  or (_11416_, _11415_, _11360_);
  and (_11417_, _11416_, _03455_);
  or (_11418_, _11417_, _03903_);
  or (_11419_, _11418_, _11414_);
  and (_11420_, _11419_, _11366_);
  or (_11421_, _11420_, _03897_);
  and (_11422_, _11203_, _05505_);
  or (_11423_, _11360_, _04790_);
  or (_11424_, _11423_, _11422_);
  and (_11425_, _11424_, _04792_);
  and (_11426_, _11425_, _11421_);
  or (_11427_, _11426_, _11363_);
  and (_11428_, _11427_, _03909_);
  or (_11429_, _11360_, _11028_);
  and (_11430_, _11365_, _03908_);
  and (_11431_, _11430_, _11429_);
  or (_11432_, _11431_, _11428_);
  and (_11433_, _11432_, _04785_);
  and (_11434_, _11376_, _04027_);
  and (_11435_, _11434_, _11429_);
  or (_11436_, _11435_, _03914_);
  or (_11437_, _11436_, _11433_);
  and (_11438_, _11201_, _05505_);
  or (_11439_, _11360_, _06567_);
  or (_11440_, _11439_, _11438_);
  and (_11441_, _11440_, _06572_);
  and (_11442_, _11441_, _11437_);
  and (_11443_, _11004_, _05505_);
  or (_11444_, _11443_, _11360_);
  and (_11445_, _11444_, _04011_);
  or (_11446_, _11445_, _03773_);
  or (_11447_, _11446_, _11442_);
  or (_11448_, _11373_, _03774_);
  and (_11449_, _11448_, _03375_);
  and (_11450_, _11449_, _11447_);
  and (_11451_, _11370_, _03374_);
  or (_11452_, _11451_, _03772_);
  or (_11453_, _11452_, _11450_);
  and (_11454_, _11249_, _05505_);
  or (_11455_, _11360_, _04060_);
  or (_11456_, _11455_, _11454_);
  and (_11457_, _11456_, _43152_);
  and (_11458_, _11457_, _11453_);
  nor (_11459_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_11460_, _11459_, _05397_);
  or (_40702_, _11460_, _11458_);
  not (_11461_, _05455_);
  and (_11462_, _11461_, \oc8051_golden_model_1.P1 [7]);
  and (_11463_, _11006_, _05455_);
  or (_11464_, _11463_, _11462_);
  and (_11465_, _11464_, _04018_);
  and (_11466_, _06348_, _05455_);
  or (_11467_, _11466_, _11462_);
  or (_11468_, _11467_, _04778_);
  not (_11469_, _06114_);
  and (_11470_, _11469_, \oc8051_golden_model_1.P1 [7]);
  and (_11471_, _11024_, _06114_);
  or (_11472_, _11471_, _11470_);
  and (_11473_, _11472_, _03759_);
  and (_11474_, _11135_, _05455_);
  or (_11475_, _11474_, _11462_);
  or (_11476_, _11475_, _04722_);
  and (_11477_, _05455_, \oc8051_golden_model_1.ACC [7]);
  or (_11478_, _11477_, _11462_);
  and (_11479_, _11478_, _04707_);
  and (_11480_, _04708_, \oc8051_golden_model_1.P1 [7]);
  or (_11481_, _11480_, _03850_);
  or (_11482_, _11481_, _11479_);
  and (_11483_, _11482_, _03764_);
  and (_11484_, _11483_, _11476_);
  and (_11485_, _11147_, _06114_);
  or (_11486_, _11485_, _11470_);
  and (_11487_, _11486_, _03763_);
  or (_11488_, _11487_, _03848_);
  or (_11489_, _11488_, _11484_);
  and (_11490_, _05568_, _05455_);
  or (_11491_, _11490_, _11462_);
  or (_11492_, _11491_, _04733_);
  and (_11493_, _11492_, _11489_);
  or (_11494_, _11493_, _03854_);
  or (_11495_, _11478_, _03855_);
  and (_11496_, _11495_, _03760_);
  and (_11497_, _11496_, _11494_);
  or (_11498_, _11497_, _11473_);
  and (_11499_, _11498_, _03753_);
  or (_11500_, _11470_, _11163_);
  and (_11501_, _11486_, _03752_);
  and (_11502_, _11501_, _11500_);
  or (_11503_, _11502_, _11499_);
  and (_11504_, _11503_, _03747_);
  and (_11505_, _11169_, _06114_);
  or (_11506_, _11505_, _11470_);
  and (_11507_, _11506_, _03746_);
  or (_11508_, _11507_, _07927_);
  or (_11509_, _11508_, _11504_);
  and (_11510_, _06248_, _05455_);
  or (_11511_, _11462_, _03738_);
  or (_11512_, _11511_, _11510_);
  or (_11513_, _11491_, _07925_);
  and (_11514_, _11513_, _03820_);
  and (_11515_, _11514_, _11512_);
  and (_11516_, _11515_, _11509_);
  and (_11517_, _11193_, _05455_);
  or (_11518_, _11517_, _11462_);
  and (_11519_, _11518_, _03455_);
  or (_11520_, _11519_, _03903_);
  or (_11521_, _11520_, _11516_);
  and (_11522_, _11521_, _11468_);
  or (_11523_, _11522_, _03897_);
  and (_11524_, _11203_, _05455_);
  or (_11525_, _11462_, _04790_);
  or (_11526_, _11525_, _11524_);
  and (_11527_, _11526_, _04792_);
  and (_11528_, _11527_, _11523_);
  or (_11529_, _11528_, _11465_);
  and (_11530_, _11529_, _03909_);
  or (_11531_, _11462_, _11028_);
  and (_11532_, _11467_, _03908_);
  and (_11533_, _11532_, _11531_);
  or (_11534_, _11533_, _11530_);
  and (_11535_, _11534_, _04785_);
  and (_11536_, _11478_, _04027_);
  and (_11537_, _11536_, _11531_);
  or (_11538_, _11537_, _03914_);
  or (_11539_, _11538_, _11535_);
  and (_11540_, _11201_, _05455_);
  or (_11541_, _11462_, _06567_);
  or (_11542_, _11541_, _11540_);
  and (_11543_, _11542_, _06572_);
  and (_11544_, _11543_, _11539_);
  and (_11545_, _11004_, _05455_);
  or (_11546_, _11545_, _11462_);
  and (_11547_, _11546_, _04011_);
  or (_11548_, _11547_, _03773_);
  or (_11549_, _11548_, _11544_);
  or (_11550_, _11475_, _03774_);
  and (_11551_, _11550_, _03375_);
  and (_11552_, _11551_, _11549_);
  and (_11553_, _11472_, _03374_);
  or (_11554_, _11553_, _03772_);
  or (_11555_, _11554_, _11552_);
  and (_11556_, _11249_, _05455_);
  or (_11557_, _11462_, _04060_);
  or (_11558_, _11557_, _11556_);
  and (_11559_, _11558_, _43152_);
  and (_11560_, _11559_, _11555_);
  nor (_11561_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_11562_, _11561_, _05397_);
  or (_40703_, _11562_, _11560_);
  not (_11563_, \oc8051_golden_model_1.SP [7]);
  nor (_11564_, _43152_, _11563_);
  and (_11565_, _05127_, \oc8051_golden_model_1.SP [4]);
  and (_11566_, _11565_, \oc8051_golden_model_1.SP [5]);
  and (_11567_, _11566_, \oc8051_golden_model_1.SP [6]);
  or (_11568_, _11567_, \oc8051_golden_model_1.SP [7]);
  nand (_11569_, _11567_, \oc8051_golden_model_1.SP [7]);
  and (_11570_, _11569_, _11568_);
  or (_11571_, _11570_, _04819_);
  nor (_11572_, _05516_, _11563_);
  and (_11573_, _06557_, _05516_);
  or (_11574_, _11573_, _11572_);
  and (_11575_, _11574_, _04018_);
  and (_11576_, _05568_, _05516_);
  or (_11577_, _11572_, _03737_);
  or (_11578_, _11577_, _11576_);
  and (_11579_, _11578_, _07927_);
  and (_11580_, _06160_, _05516_);
  or (_11581_, _11580_, _11572_);
  or (_11582_, _11581_, _04722_);
  and (_11583_, _05516_, \oc8051_golden_model_1.ACC [7]);
  or (_11584_, _11583_, _11572_);
  or (_11585_, _11584_, _04708_);
  or (_11586_, _04707_, \oc8051_golden_model_1.SP [7]);
  and (_11587_, _11586_, _03770_);
  and (_11588_, _11587_, _11585_);
  and (_11589_, _11570_, _03768_);
  or (_11590_, _11589_, _03850_);
  or (_11591_, _11590_, _11588_);
  and (_11592_, _11591_, _03431_);
  and (_11593_, _11592_, _11582_);
  and (_11594_, _11570_, _05045_);
  or (_11595_, _11594_, _03848_);
  or (_11596_, _11595_, _11593_);
  not (_11597_, \oc8051_golden_model_1.SP [6]);
  not (_11598_, \oc8051_golden_model_1.SP [5]);
  not (_11599_, \oc8051_golden_model_1.SP [4]);
  and (_11600_, _06166_, _11599_);
  and (_11601_, _11600_, _11598_);
  and (_11602_, _11601_, _11597_);
  and (_11603_, _11602_, _03683_);
  nor (_11604_, _11603_, _11563_);
  and (_11605_, _11603_, _11563_);
  nor (_11606_, _11605_, _11604_);
  nand (_11607_, _11606_, _03848_);
  and (_11608_, _11607_, _11596_);
  or (_11609_, _11608_, _03854_);
  or (_11610_, _11584_, _03855_);
  and (_11611_, _11610_, _04845_);
  and (_11612_, _11611_, _11609_);
  and (_11613_, _11566_, \oc8051_golden_model_1.SP [0]);
  and (_11614_, _11613_, \oc8051_golden_model_1.SP [6]);
  or (_11615_, _11614_, \oc8051_golden_model_1.SP [7]);
  nand (_11616_, _11614_, \oc8051_golden_model_1.SP [7]);
  and (_11617_, _11616_, _11615_);
  nand (_11618_, _11617_, _03758_);
  nand (_11619_, _11618_, _05050_);
  or (_11620_, _11619_, _11612_);
  or (_11621_, _11570_, _05050_);
  and (_11622_, _11621_, _07925_);
  and (_11623_, _11622_, _11620_);
  or (_11624_, _11623_, _11579_);
  and (_11625_, _06248_, _05516_);
  or (_11626_, _11572_, _03738_);
  or (_11627_, _11626_, _11625_);
  and (_11628_, _11627_, _03820_);
  and (_11629_, _11628_, _11624_);
  not (_11630_, _05516_);
  nor (_11631_, _06536_, _11630_);
  or (_11632_, _11631_, _11572_);
  and (_11633_, _11632_, _03455_);
  or (_11634_, _11633_, _03903_);
  or (_11635_, _11634_, _11629_);
  and (_11636_, _06348_, _05516_);
  or (_11637_, _11636_, _11572_);
  or (_11638_, _11637_, _04778_);
  and (_11639_, _11638_, _11635_);
  or (_11640_, _11639_, _03401_);
  not (_11641_, _03401_);
  or (_11642_, _11570_, _11641_);
  and (_11643_, _11642_, _11640_);
  or (_11644_, _11643_, _03897_);
  and (_11645_, _06549_, _05516_);
  or (_11646_, _11572_, _04790_);
  or (_11647_, _11646_, _11645_);
  and (_11648_, _11647_, _04792_);
  and (_11649_, _11648_, _11644_);
  or (_11650_, _11649_, _11575_);
  and (_11651_, _11650_, _03909_);
  or (_11652_, _11572_, _05571_);
  and (_11653_, _11637_, _03908_);
  and (_11654_, _11653_, _11652_);
  or (_11655_, _11654_, _11651_);
  and (_11656_, _11655_, _10076_);
  and (_11657_, _11584_, _04027_);
  and (_11658_, _11657_, _11652_);
  and (_11659_, _11570_, _03388_);
  or (_11660_, _11659_, _03914_);
  or (_11661_, _11660_, _11658_);
  or (_11662_, _11661_, _11656_);
  nor (_11663_, _06547_, _11630_);
  or (_11664_, _11663_, _11572_);
  or (_11665_, _11664_, _06567_);
  and (_11666_, _11665_, _11662_);
  or (_11667_, _11666_, _04011_);
  nor (_11668_, _06556_, _11630_);
  or (_11669_, _11572_, _06572_);
  or (_11670_, _11669_, _11668_);
  and (_11671_, _11670_, _10704_);
  and (_11672_, _11671_, _11667_);
  or (_11673_, _11602_, \oc8051_golden_model_1.SP [7]);
  nand (_11674_, _11602_, \oc8051_golden_model_1.SP [7]);
  and (_11675_, _11674_, _11673_);
  and (_11676_, _11675_, _04034_);
  or (_11677_, _11676_, _03383_);
  or (_11678_, _11677_, _11672_);
  or (_11679_, _11570_, _03384_);
  and (_11680_, _11679_, _11678_);
  or (_11681_, _11680_, _03777_);
  or (_11682_, _11675_, _03778_);
  and (_11683_, _11682_, _03774_);
  and (_11684_, _11683_, _11681_);
  and (_11685_, _11581_, _03773_);
  or (_11686_, _11685_, _05223_);
  or (_11687_, _11686_, _11684_);
  and (_11688_, _11687_, _11571_);
  or (_11689_, _11688_, _03772_);
  and (_11690_, _06077_, _05516_);
  or (_11691_, _11572_, _04060_);
  or (_11692_, _11691_, _11690_);
  and (_11693_, _11692_, _43152_);
  and (_11694_, _11693_, _11689_);
  or (_11695_, _11694_, _11564_);
  and (_40704_, _11695_, _41894_);
  nor (_11696_, _43152_, _08297_);
  nor (_11697_, _06094_, _08297_);
  and (_11698_, _06121_, _06094_);
  or (_11699_, _11698_, _11697_);
  or (_11700_, _11699_, _03375_);
  and (_11701_, _08044_, \oc8051_golden_model_1.ACC [7]);
  or (_11702_, _11701_, _08109_);
  or (_11703_, _08119_, _08041_);
  or (_11704_, _11703_, _11702_);
  nor (_11705_, _05424_, _08297_);
  and (_11706_, _06557_, _05424_);
  or (_11707_, _11706_, _11705_);
  and (_11708_, _11707_, _04018_);
  not (_11709_, _05424_);
  nor (_11710_, _06536_, _11709_);
  or (_11711_, _11710_, _11705_);
  and (_11712_, _11711_, _03455_);
  and (_11713_, _08338_, _08335_);
  and (_11714_, _11713_, _06071_);
  and (_11715_, _08334_, _08330_);
  nor (_11716_, _11715_, _08328_);
  nand (_11717_, _08384_, _08330_);
  or (_11718_, _11717_, _08382_);
  and (_11719_, _11718_, _11716_);
  or (_11720_, _11719_, _11714_);
  and (_11721_, _11720_, _03883_);
  and (_11722_, _08260_, _08255_);
  nor (_11723_, _11722_, _08253_);
  nand (_11724_, _08310_, _08255_);
  or (_11725_, _11724_, _08308_);
  and (_11726_, _11725_, _11723_);
  and (_11727_, _08249_, _06248_);
  or (_11728_, _11727_, _08248_);
  or (_11729_, _11728_, _11726_);
  not (_11730_, _03878_);
  not (_11731_, _03879_);
  nor (_11732_, _10906_, _11731_);
  or (_11733_, _10245_, _10243_);
  and (_11734_, _11733_, _10240_);
  and (_11735_, _10238_, _10235_);
  or (_11736_, _11735_, _10233_);
  or (_11737_, _11736_, _11734_);
  and (_11738_, _11737_, _10232_);
  nor (_11739_, _10228_, _10226_);
  nor (_11740_, _11739_, _10225_);
  and (_11741_, _11740_, _10224_);
  nor (_11742_, _10221_, _10219_);
  nor (_11743_, _11742_, _06291_);
  or (_11744_, _11743_, _11741_);
  or (_11745_, _11744_, _11738_);
  and (_11746_, _11745_, _10250_);
  or (_11747_, _11746_, _10444_);
  and (_11748_, _06160_, _05424_);
  or (_11749_, _11748_, _11705_);
  or (_11750_, _11749_, _04722_);
  not (_11751_, _08179_);
  and (_11752_, _05424_, \oc8051_golden_model_1.ACC [7]);
  or (_11753_, _11752_, _11705_);
  and (_11754_, _11753_, _04707_);
  nor (_11755_, _04707_, _08297_);
  or (_11756_, _11755_, _03850_);
  or (_11757_, _11756_, _11754_);
  and (_11758_, _11757_, _11751_);
  and (_11759_, _11758_, _11750_);
  nor (_11760_, _08189_, \oc8051_golden_model_1.PSW [7]);
  not (_11761_, _11760_);
  nor (_11762_, _11761_, _08199_);
  nor (_11763_, _11762_, _11751_);
  not (_11764_, _10411_);
  nand (_11765_, _11764_, _03856_);
  or (_11766_, _11765_, _11763_);
  or (_11767_, _11766_, _11759_);
  and (_11768_, _06148_, _06094_);
  or (_11769_, _11768_, _11697_);
  or (_11770_, _11769_, _03764_);
  and (_11771_, _05568_, _05424_);
  or (_11772_, _11771_, _11705_);
  or (_11773_, _11772_, _04733_);
  and (_11774_, _11773_, _11770_);
  and (_11775_, _11774_, _11767_);
  or (_11776_, _11775_, _03854_);
  nor (_11777_, _11753_, _03855_);
  nor (_11778_, _11777_, _10430_);
  and (_11779_, _11778_, _11776_);
  or (_11780_, _11779_, _03759_);
  or (_11781_, _11699_, _03760_);
  and (_11782_, _11781_, _10441_);
  and (_11783_, _11782_, _11780_);
  and (_11784_, _10447_, _10448_);
  or (_11785_, _11784_, _10445_);
  or (_11786_, _10457_, _10455_);
  and (_11787_, _11786_, _10451_);
  or (_11788_, _11787_, _11785_);
  and (_11789_, _11788_, _10474_);
  or (_11790_, _10470_, _10467_);
  nand (_11791_, _11790_, _10466_);
  nor (_11792_, _11791_, _10468_);
  and (_11793_, _10464_, _06079_);
  or (_11794_, _11793_, _10461_);
  or (_11795_, _11794_, _11792_);
  or (_11796_, _11795_, _11789_);
  nor (_11797_, _10476_, _10441_);
  and (_11798_, _11797_, _11796_);
  or (_11799_, _11798_, _03925_);
  or (_11800_, _11799_, _11783_);
  and (_11801_, _11800_, _03918_);
  and (_11802_, _11801_, _11747_);
  nor (_11803_, _05669_, \oc8051_golden_model_1.ACC [1]);
  and (_11804_, _05716_, \oc8051_golden_model_1.ACC [0]);
  nor (_11805_, _11804_, _08752_);
  or (_11806_, _11805_, _11803_);
  and (_11807_, _11806_, _10497_);
  nor (_11808_, _05570_, \oc8051_golden_model_1.ACC [7]);
  or (_11809_, _06068_, \oc8051_golden_model_1.ACC [6]);
  nor (_11810_, _11809_, _06557_);
  or (_11811_, _11810_, _11808_);
  nand (_11812_, _05859_, \oc8051_golden_model_1.ACC [5]);
  nor (_11813_, _05859_, \oc8051_golden_model_1.ACC [5]);
  nor (_11814_, _05953_, \oc8051_golden_model_1.ACC [4]);
  or (_11815_, _11814_, _11813_);
  and (_11816_, _11815_, _11812_);
  and (_11817_, _11816_, _10495_);
  or (_11818_, _11817_, _11811_);
  nand (_11819_, _05621_, \oc8051_golden_model_1.ACC [3]);
  nor (_11820_, _05621_, \oc8051_golden_model_1.ACC [3]);
  nor (_11821_, _05764_, \oc8051_golden_model_1.ACC [2]);
  or (_11822_, _11821_, _11820_);
  and (_11823_, _11822_, _11819_);
  and (_11824_, _11823_, _10496_);
  or (_11825_, _11824_, _11818_);
  or (_11826_, _11825_, _11807_);
  nor (_11827_, _10498_, _03918_);
  and (_11828_, _11827_, _11826_);
  or (_11829_, _11828_, _11802_);
  and (_11830_, _11829_, _10486_);
  and (_11831_, _10485_, _08297_);
  or (_11832_, _03810_, \oc8051_golden_model_1.ACC [6]);
  nor (_11833_, _11832_, _08537_);
  and (_11834_, _03647_, _06554_);
  or (_11835_, _11834_, _11833_);
  nand (_11836_, _04093_, \oc8051_golden_model_1.ACC [5]);
  nor (_11837_, _04093_, \oc8051_golden_model_1.ACC [5]);
  nor (_11838_, _04526_, \oc8051_golden_model_1.ACC [4]);
  or (_11839_, _11838_, _11837_);
  and (_11840_, _11839_, _11836_);
  and (_11841_, _11840_, _10512_);
  or (_11842_, _11841_, _11835_);
  nor (_11843_, _04563_, \oc8051_golden_model_1.ACC [1]);
  and (_11844_, _04563_, \oc8051_golden_model_1.ACC [1]);
  and (_11845_, _03715_, \oc8051_golden_model_1.ACC [0]);
  nor (_11846_, _11845_, _11844_);
  or (_11847_, _11846_, _11843_);
  and (_11848_, _11847_, _10510_);
  nand (_11849_, _03678_, \oc8051_golden_model_1.ACC [3]);
  nor (_11850_, _03678_, \oc8051_golden_model_1.ACC [3]);
  nor (_11851_, _04139_, \oc8051_golden_model_1.ACC [2]);
  or (_11852_, _11851_, _11850_);
  and (_11853_, _11852_, _11849_);
  or (_11854_, _11853_, _11848_);
  and (_11855_, _11854_, _10513_);
  or (_11856_, _11855_, _11842_);
  not (_11857_, _03920_);
  nor (_11858_, _10515_, _11857_);
  and (_11859_, _11858_, _11856_);
  or (_11860_, _11859_, _11831_);
  or (_11861_, _11860_, _11830_);
  and (_11862_, _11861_, _03844_);
  and (_11863_, _10906_, \oc8051_golden_model_1.PSW [7]);
  and (_11864_, _11863_, _03843_);
  or (_11865_, _11697_, _06147_);
  and (_11866_, _11865_, _03752_);
  and (_11867_, _11866_, _11769_);
  or (_11868_, _11867_, _11864_);
  or (_11869_, _11868_, _11862_);
  nor (_11870_, _07399_, _03879_);
  and (_11871_, _11870_, _11869_);
  or (_11872_, _11871_, _11732_);
  and (_11873_, _11872_, _11730_);
  or (_11874_, _10906_, \oc8051_golden_model_1.PSW [7]);
  and (_11875_, _11874_, _03878_);
  nand (_11876_, _03825_, _03424_);
  or (_11877_, _08150_, _04333_);
  nor (_11878_, _11877_, _08151_);
  and (_11879_, _11878_, _11876_);
  not (_11880_, _11879_);
  or (_11881_, _11880_, _11875_);
  or (_11882_, _11881_, _11873_);
  not (_11883_, _04335_);
  and (_11884_, _08051_, _08047_);
  nor (_11885_, _11884_, _08045_);
  and (_11886_, _08053_, _08047_);
  not (_11887_, _11886_);
  or (_11888_, _11887_, _08142_);
  and (_11889_, _11888_, _11885_);
  or (_11890_, _11889_, _08041_);
  or (_11891_, _11890_, _11879_);
  and (_11892_, _11891_, _11883_);
  and (_11893_, _11892_, _11882_);
  and (_11894_, _11890_, _04335_);
  or (_11895_, _11894_, _04330_);
  or (_11896_, _11895_, _11893_);
  and (_11897_, _11896_, _11729_);
  and (_11898_, _11897_, _03888_);
  or (_11899_, _11898_, _11721_);
  and (_11900_, _11899_, _08321_);
  and (_11901_, _08400_, _05422_);
  and (_11902_, _08409_, _08405_);
  nor (_11903_, _11902_, _08403_);
  and (_11904_, _08411_, _08405_);
  and (_11905_, _11904_, _08453_);
  not (_11906_, _11905_);
  and (_11907_, _11906_, _11903_);
  or (_11908_, _11907_, _11901_);
  and (_11909_, _11908_, _08320_);
  or (_11910_, _11909_, _07927_);
  or (_11911_, _11910_, _11900_);
  and (_11912_, _06248_, _05424_);
  or (_11913_, _11705_, _03738_);
  or (_11914_, _11913_, _11912_);
  or (_11915_, _11772_, _07925_);
  and (_11916_, _11915_, _03820_);
  and (_11917_, _11916_, _11914_);
  and (_11918_, _11917_, _11911_);
  or (_11919_, _11918_, _11712_);
  nor (_11920_, _07010_, _03816_);
  and (_11921_, _11920_, _11919_);
  nor (_11922_, _10906_, _08297_);
  and (_11923_, _11922_, _03816_);
  or (_11924_, _11923_, _03903_);
  or (_11925_, _11924_, _11921_);
  and (_11926_, _06348_, _05424_);
  or (_11927_, _11926_, _11705_);
  or (_11928_, _11927_, _04778_);
  and (_11929_, _11928_, _11925_);
  and (_11930_, _11929_, _04391_);
  nand (_11931_, _10906_, _08297_);
  and (_11932_, _11931_, _03815_);
  or (_11933_, _11932_, _11930_);
  or (_11934_, _11933_, _03897_);
  and (_11935_, _06549_, _05424_);
  or (_11936_, _11935_, _11705_);
  or (_11937_, _11936_, _04790_);
  and (_11938_, _11937_, _04792_);
  and (_11939_, _11938_, _11934_);
  or (_11940_, _11939_, _11708_);
  and (_11941_, _11940_, _03909_);
  or (_11942_, _11705_, _05571_);
  and (_11943_, _11927_, _03908_);
  and (_11944_, _11943_, _11942_);
  or (_11945_, _11944_, _11941_);
  and (_11946_, _11945_, _04785_);
  and (_11947_, _11753_, _04027_);
  and (_11948_, _11947_, _11942_);
  or (_11949_, _11948_, _03914_);
  or (_11950_, _11949_, _11946_);
  nor (_11951_, _06547_, _11709_);
  or (_11952_, _11705_, _06567_);
  or (_11953_, _11952_, _11951_);
  and (_11954_, _11953_, _06572_);
  and (_11955_, _11954_, _11950_);
  nor (_11956_, _06556_, _11709_);
  or (_11957_, _11956_, _11705_);
  and (_11958_, _11957_, _04011_);
  or (_11959_, _11958_, _08590_);
  or (_11960_, _11959_, _11955_);
  and (_11961_, _11960_, _11704_);
  or (_11962_, _11961_, _08597_);
  or (_11963_, _11727_, _08599_);
  nor (_11964_, _08252_, _06554_);
  or (_11965_, _11964_, _08621_);
  or (_11966_, _11965_, _11963_);
  and (_11967_, _11966_, _04023_);
  and (_11968_, _11967_, _11962_);
  nor (_11969_, _08327_, _06554_);
  or (_11970_, _11969_, _08651_);
  or (_11971_, _11970_, _11714_);
  and (_11972_, _11971_, _04022_);
  or (_11973_, _11972_, _08627_);
  or (_11974_, _11973_, _11968_);
  and (_11975_, _08402_, \oc8051_golden_model_1.ACC [7]);
  or (_11976_, _11975_, _08681_);
  or (_11977_, _11976_, _11901_);
  or (_11978_, _11977_, _08659_);
  and (_11979_, _11978_, _08658_);
  and (_11980_, _11979_, _11974_);
  nand (_11981_, _08657_, \oc8051_golden_model_1.ACC [7]);
  and (_11982_, _08115_, _03409_);
  not (_11983_, _11982_);
  and (_11984_, _11983_, _07997_);
  nand (_11985_, _11984_, _11981_);
  or (_11986_, _11985_, _11980_);
  not (_11987_, _04456_);
  not (_11988_, _08001_);
  or (_11989_, _08034_, _08000_);
  nand (_11990_, _11989_, _11988_);
  or (_11991_, _11990_, _11984_);
  and (_11992_, _11991_, _11987_);
  and (_11993_, _11992_, _11986_);
  and (_11994_, _11990_, _04456_);
  or (_11995_, _11994_, _08691_);
  or (_11996_, _11995_, _11993_);
  and (_11997_, _08725_, _08526_);
  nor (_11998_, _08695_, _08525_);
  nor (_11999_, _11998_, _08524_);
  or (_12000_, _11999_, _10058_);
  or (_12001_, _12000_, _11997_);
  and (_12002_, _12001_, _04140_);
  and (_12003_, _12002_, _11996_);
  not (_12004_, _06556_);
  not (_12005_, _06555_);
  nand (_12006_, _08765_, _12005_);
  and (_12007_, _12006_, _03779_);
  and (_12008_, _12007_, _12004_);
  or (_12009_, _12008_, _08733_);
  or (_12010_, _12009_, _12003_);
  or (_12011_, _08805_, _08535_);
  nand (_12012_, _12011_, _08733_);
  or (_12013_, _12012_, _08536_);
  and (_12014_, _12013_, _12010_);
  or (_12015_, _12014_, _03773_);
  not (_12016_, _08820_);
  or (_12017_, _11749_, _03774_);
  and (_12018_, _12017_, _12016_);
  and (_12019_, _12018_, _12015_);
  and (_12020_, _08820_, \oc8051_golden_model_1.ACC [0]);
  or (_12021_, _12020_, _03374_);
  or (_12022_, _12021_, _12019_);
  and (_12023_, _12022_, _11700_);
  or (_12024_, _12023_, _03772_);
  and (_12025_, _06077_, _05424_);
  or (_12026_, _11705_, _04060_);
  or (_12027_, _12026_, _12025_);
  and (_12028_, _12027_, _43152_);
  and (_12029_, _12028_, _12024_);
  or (_12030_, _12029_, _11696_);
  and (_40705_, _12030_, _41894_);
  and (_12031_, _43156_, \oc8051_golden_model_1.P0INREG [7]);
  or (_12032_, _12031_, _01158_);
  and (_40707_, _12032_, _41894_);
  and (_12033_, _43156_, \oc8051_golden_model_1.P1INREG [7]);
  or (_12034_, _12033_, _01313_);
  and (_40708_, _12034_, _41894_);
  and (_12035_, _43156_, \oc8051_golden_model_1.P2INREG [7]);
  or (_12036_, _12035_, _01225_);
  and (_40709_, _12036_, _41894_);
  and (_12037_, _43156_, \oc8051_golden_model_1.P3INREG [7]);
  or (_12038_, _12037_, _01371_);
  and (_40710_, _12038_, _41894_);
  and (_12039_, _05071_, _04834_);
  nor (_12040_, _12039_, _05073_);
  nor (_12041_, _05242_, _05072_);
  nor (_12042_, _12041_, _05386_);
  and (_12043_, _12042_, _05071_);
  and (_12044_, _12043_, _12040_);
  or (_12045_, _12044_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_12046_, _05399_, _04990_);
  not (_12047_, _12046_);
  not (_12048_, _04838_);
  and (_12049_, _12046_, _05393_);
  and (_12050_, _12046_, _05396_);
  or (_12051_, _12050_, _12049_);
  or (_12052_, _12051_, _12048_);
  or (_12053_, _12052_, _12047_);
  and (_12054_, _12053_, _12045_);
  not (_12055_, _12044_);
  nand (_12056_, _03414_, _03119_);
  nand (_12057_, _10488_, _06573_);
  nor (_12058_, _05716_, _04382_);
  and (_12059_, _12058_, _04788_);
  or (_12060_, _03735_, _04700_);
  and (_12061_, _06962_, _05421_);
  or (_12062_, _12061_, _05714_);
  and (_12063_, _12062_, _04939_);
  nand (_12064_, _10820_, _10796_);
  nand (_12065_, _12064_, _03755_);
  nor (_12066_, _12065_, _10821_);
  and (_12067_, _03768_, \oc8051_golden_model_1.PC [0]);
  nor (_12068_, _03768_, _03498_);
  or (_12069_, _12068_, _12067_);
  or (_12070_, _12069_, _04267_);
  nand (_12071_, _04700_, _04267_);
  and (_12072_, _12071_, _12070_);
  and (_12073_, _12072_, _06250_);
  and (_12074_, _05716_, _04723_);
  or (_12075_, _12074_, _12073_);
  or (_12076_, _12075_, _04721_);
  or (_12077_, _12064_, _05152_);
  and (_12078_, _12077_, _12076_);
  and (_12079_, _12078_, _03431_);
  nor (_12080_, _03431_, _03119_);
  or (_12081_, _04734_, _12080_);
  or (_12082_, _12081_, _12079_);
  or (_12083_, _05132_, _04700_);
  and (_12084_, _12083_, _05005_);
  and (_12085_, _12084_, _12082_);
  nor (_12086_, _10820_, _05432_);
  and (_12087_, _12086_, _04743_);
  or (_12088_, _12087_, _03758_);
  or (_12089_, _12088_, _12085_);
  nand (_12090_, _05716_, _03758_);
  and (_12091_, _12090_, _03756_);
  and (_12092_, _12091_, _12089_);
  or (_12093_, _12092_, _12066_);
  and (_12094_, _12093_, _03428_);
  or (_12095_, _03428_, _03119_);
  nand (_12096_, _03840_, _12095_);
  or (_12097_, _12096_, _12094_);
  nand (_12098_, _05716_, _03841_);
  and (_12099_, _12098_, _04940_);
  and (_12100_, _12099_, _12097_);
  or (_12101_, _12100_, _12063_);
  and (_12102_, _12101_, _05183_);
  and (_12103_, _05432_, \oc8051_golden_model_1.PSW [7]);
  nor (_12104_, _12103_, _12086_);
  nor (_12105_, _12104_, _05183_);
  or (_12106_, _12105_, _12102_);
  and (_12107_, _12106_, _06141_);
  nand (_12108_, _03456_, \oc8051_golden_model_1.PC [0]);
  nand (_12109_, _03735_, _12108_);
  or (_12110_, _12109_, _12107_);
  and (_12111_, _12110_, _12060_);
  or (_12112_, _12111_, _03739_);
  or (_12113_, _06962_, _06305_);
  and (_12114_, _12113_, _06304_);
  and (_12115_, _12114_, _12112_);
  and (_12116_, _06342_, _04700_);
  and (_12117_, _06519_, \oc8051_golden_model_1.SP [0]);
  not (_12118_, _12117_);
  and (_12119_, _06522_, \oc8051_golden_model_1.IE [0]);
  not (_12120_, _12119_);
  and (_12121_, _06525_, \oc8051_golden_model_1.SCON [0]);
  and (_12122_, _06527_, \oc8051_golden_model_1.SBUF [0]);
  nor (_12123_, _12122_, _12121_);
  and (_12124_, _12123_, _12120_);
  and (_12125_, _06512_, \oc8051_golden_model_1.TMOD [0]);
  not (_12126_, _12125_);
  and (_12127_, _06505_, \oc8051_golden_model_1.P1INREG [0]);
  and (_12128_, _06507_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_12129_, _12128_, _12127_);
  and (_12130_, _12129_, _12126_);
  and (_12131_, _12130_, _12124_);
  and (_12132_, _12131_, _12118_);
  and (_12133_, _06477_, \oc8051_golden_model_1.DPH [0]);
  and (_12134_, _06483_, \oc8051_golden_model_1.TH1 [0]);
  nor (_12135_, _12134_, _12133_);
  and (_12136_, _06472_, \oc8051_golden_model_1.TL0 [0]);
  not (_12137_, _12136_);
  and (_12138_, _06501_, \oc8051_golden_model_1.P0INREG [0]);
  and (_12139_, _06515_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_12140_, _12139_, _12138_);
  and (_12141_, _12140_, _12137_);
  and (_12142_, _12141_, _12135_);
  and (_12143_, _12142_, _12132_);
  and (_12144_, _06488_, \oc8051_golden_model_1.TH0 [0]);
  and (_12145_, _06490_, \oc8051_golden_model_1.TL1 [0]);
  nor (_12146_, _12145_, _12144_);
  and (_12147_, _06493_, \oc8051_golden_model_1.TCON [0]);
  and (_12148_, _06497_, \oc8051_golden_model_1.PCON [0]);
  nor (_12149_, _12148_, _12147_);
  and (_12150_, _12149_, _12146_);
  and (_12151_, _06469_, \oc8051_golden_model_1.DPL [0]);
  not (_12152_, _12151_);
  and (_12153_, _06445_, \oc8051_golden_model_1.IP [0]);
  and (_12154_, _06460_, \oc8051_golden_model_1.B [0]);
  nor (_12155_, _12154_, _12153_);
  and (_12156_, _06458_, \oc8051_golden_model_1.PSW [0]);
  and (_12157_, _06453_, \oc8051_golden_model_1.ACC [0]);
  nor (_12158_, _12157_, _12156_);
  and (_12159_, _12158_, _12155_);
  and (_12160_, _12159_, _12152_);
  and (_12161_, _12160_, _12150_);
  and (_12162_, _12161_, _12143_);
  not (_12163_, _12162_);
  nor (_12164_, _12163_, _12116_);
  nor (_12165_, _12164_, _06311_);
  or (_12166_, _12165_, _06309_);
  or (_12167_, _12166_, _12115_);
  and (_12168_, _06309_, _03715_);
  nor (_12169_, _12168_, _04779_);
  and (_12170_, _12169_, _12167_);
  and (_12171_, _04779_, _06479_);
  or (_12172_, _12171_, _03401_);
  or (_12173_, _12172_, _12170_);
  and (_12174_, _03401_, _03119_);
  nor (_12175_, _12174_, _04791_);
  and (_12176_, _12175_, _12173_);
  and (_12177_, _05716_, _04382_);
  nor (_12178_, _12177_, _12058_);
  nor (_12179_, _12178_, _04793_);
  nor (_12180_, _12179_, _04794_);
  or (_12181_, _12180_, _12176_);
  nand (_12182_, _10489_, _04793_);
  and (_12183_, _12182_, _04789_);
  and (_12184_, _12183_, _12181_);
  or (_12185_, _12184_, _12059_);
  and (_12186_, _12185_, _04787_);
  and (_12187_, _08753_, _04786_);
  or (_12188_, _12187_, _03388_);
  or (_12189_, _12188_, _12186_);
  and (_12190_, _03388_, _03119_);
  nor (_12191_, _12190_, _06568_);
  and (_12192_, _12191_, _12189_);
  nor (_12193_, _12177_, _06574_);
  or (_12194_, _12193_, _06573_);
  or (_12195_, _12194_, _12192_);
  and (_12196_, _12195_, _12057_);
  or (_12197_, _12196_, _03383_);
  nand (_12198_, _03383_, _03119_);
  and (_12199_, _12198_, _10935_);
  and (_12200_, _12199_, _12197_);
  nor (_12201_, _10935_, _04700_);
  or (_12202_, _12201_, _12200_);
  and (_12203_, _12202_, _04813_);
  and (_12204_, _06733_, _04812_);
  or (_12205_, _12204_, _04811_);
  or (_12206_, _12205_, _12203_);
  or (_12207_, _05716_, _06595_);
  and (_12208_, _12207_, _03900_);
  and (_12209_, _12208_, _12206_);
  and (_12210_, _03899_, _03119_);
  or (_12211_, _12210_, _03414_);
  or (_12212_, _12211_, _12209_);
  and (_12213_, _12212_, _12056_);
  or (_12214_, _12213_, _03681_);
  or (_12215_, _12086_, _03682_);
  and (_12216_, _12215_, _04482_);
  and (_12217_, _12216_, _12214_);
  nor (_12218_, _04700_, _04482_);
  or (_12219_, _12218_, _04826_);
  or (_12220_, _12219_, _12217_);
  or (_12221_, _06733_, _04827_);
  and (_12222_, _12221_, _12220_);
  or (_12223_, _12222_, _04831_);
  or (_12224_, _05716_, _06960_);
  and (_12225_, _12224_, _05071_);
  and (_12226_, _12225_, _12223_);
  or (_12227_, _12226_, _12055_);
  and (_12228_, _12227_, _12054_);
  and (_12229_, _05400_, _05393_);
  nor (_12230_, _12229_, _05401_);
  and (_12231_, _05400_, _04838_);
  and (_12232_, _12231_, _12230_);
  nand (_12233_, _10189_, _03899_);
  or (_12234_, _10349_, _03899_);
  and (_12235_, _12234_, _12233_);
  and (_12236_, _12235_, _05400_);
  and (_12237_, _12236_, _12232_);
  or (_40726_, _12237_, _12228_);
  or (_12238_, _12044_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_12239_, _12238_, _12053_);
  nor (_12240_, _06963_, _06734_);
  or (_12241_, _12240_, _04827_);
  nand (_12242_, _03899_, _03948_);
  and (_12243_, _12242_, _10953_);
  nor (_12244_, _05669_, _04595_);
  and (_12245_, _12244_, _04788_);
  or (_12246_, _04900_, _03735_);
  nand (_12247_, _05669_, _03841_);
  not (_12248_, _10766_);
  nand (_12249_, _10765_, _10741_);
  and (_12250_, _12249_, _03755_);
  and (_12251_, _12250_, _12248_);
  nor (_12252_, _10765_, _10740_);
  or (_12253_, _12252_, _05005_);
  nor (_12254_, _06945_, _06125_);
  nand (_12255_, _12254_, _04267_);
  and (_12256_, _03768_, _03087_);
  or (_12257_, _03768_, _03474_);
  nand (_12258_, _12257_, _04266_);
  or (_12259_, _12258_, _12256_);
  and (_12260_, _12259_, _12255_);
  and (_12261_, _12260_, _06250_);
  nor (_12262_, _06153_, _05717_);
  nor (_12263_, _12262_, _06250_);
  or (_12264_, _12263_, _12261_);
  or (_12265_, _12264_, _04721_);
  or (_12266_, _12249_, _05152_);
  and (_12267_, _12266_, _12265_);
  or (_12268_, _12267_, _05045_);
  nor (_12269_, _03431_, _03087_);
  nor (_12270_, _12269_, _04734_);
  and (_12271_, _12270_, _12268_);
  and (_12272_, _04900_, _04734_);
  or (_12273_, _12272_, _04743_);
  or (_12274_, _12273_, _12271_);
  and (_12275_, _12274_, _12253_);
  or (_12276_, _12275_, _03758_);
  nand (_12277_, _05669_, _03758_);
  and (_12278_, _12277_, _03756_);
  and (_12279_, _12278_, _12276_);
  or (_12280_, _12279_, _12251_);
  and (_12281_, _12280_, _03428_);
  or (_12282_, _03428_, \oc8051_golden_model_1.PC [1]);
  nand (_12283_, _03840_, _12282_);
  or (_12284_, _12283_, _12281_);
  and (_12285_, _12284_, _12247_);
  or (_12286_, _12285_, _05131_);
  and (_12287_, _06961_, _05421_);
  nand (_12288_, _05666_, _04939_);
  or (_12289_, _12288_, _12287_);
  and (_12290_, _12289_, _12286_);
  or (_12291_, _12290_, _04759_);
  and (_12292_, _10740_, \oc8051_golden_model_1.PSW [7]);
  nor (_12293_, _12292_, _12252_);
  nand (_12294_, _12293_, _04759_);
  and (_12295_, _12294_, _06141_);
  and (_12296_, _12295_, _12291_);
  nand (_12297_, _03456_, _03087_);
  nand (_12298_, _03735_, _12297_);
  or (_12299_, _12298_, _12296_);
  and (_12300_, _12299_, _12246_);
  or (_12301_, _12300_, _03739_);
  or (_12302_, _06961_, _06305_);
  and (_12303_, _12302_, _06304_);
  and (_12304_, _12303_, _12301_);
  and (_12305_, _06342_, _04900_);
  and (_12306_, _06453_, \oc8051_golden_model_1.ACC [1]);
  and (_12307_, _06458_, \oc8051_golden_model_1.PSW [1]);
  and (_12308_, _06460_, \oc8051_golden_model_1.B [1]);
  or (_12309_, _12308_, _12307_);
  nor (_12310_, _12309_, _12306_);
  and (_12311_, _06488_, \oc8051_golden_model_1.TH0 [1]);
  not (_12312_, _12311_);
  and (_12313_, _06493_, \oc8051_golden_model_1.TCON [1]);
  and (_12314_, _06445_, \oc8051_golden_model_1.IP [1]);
  nor (_12315_, _12314_, _12313_);
  and (_12316_, _12315_, _12312_);
  and (_12317_, _06497_, \oc8051_golden_model_1.PCON [1]);
  and (_12318_, _06490_, \oc8051_golden_model_1.TL1 [1]);
  nor (_12319_, _12318_, _12317_);
  and (_12320_, _12319_, _12316_);
  and (_12321_, _12320_, _12310_);
  and (_12322_, _06472_, \oc8051_golden_model_1.TL0 [1]);
  and (_12323_, _06483_, \oc8051_golden_model_1.TH1 [1]);
  nor (_12324_, _12323_, _12322_);
  and (_12325_, _06469_, \oc8051_golden_model_1.DPL [1]);
  and (_12326_, _06477_, \oc8051_golden_model_1.DPH [1]);
  nor (_12327_, _12326_, _12325_);
  and (_12328_, _12327_, _12324_);
  and (_12329_, _06512_, \oc8051_golden_model_1.TMOD [1]);
  not (_12330_, _12329_);
  and (_12331_, _06505_, \oc8051_golden_model_1.P1INREG [1]);
  and (_12332_, _06507_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_12333_, _12332_, _12331_);
  and (_12334_, _12333_, _12330_);
  and (_12335_, _06501_, \oc8051_golden_model_1.P0INREG [1]);
  and (_12336_, _06515_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_12337_, _12336_, _12335_);
  and (_12338_, _12337_, _12334_);
  and (_12339_, _06519_, \oc8051_golden_model_1.SP [1]);
  not (_12340_, _12339_);
  and (_12341_, _06522_, \oc8051_golden_model_1.IE [1]);
  not (_12342_, _12341_);
  and (_12343_, _06525_, \oc8051_golden_model_1.SCON [1]);
  and (_12344_, _06527_, \oc8051_golden_model_1.SBUF [1]);
  nor (_12345_, _12344_, _12343_);
  and (_12346_, _12345_, _12342_);
  and (_12347_, _12346_, _12340_);
  and (_12348_, _12347_, _12338_);
  and (_12349_, _12348_, _12328_);
  and (_12350_, _12349_, _12321_);
  not (_12351_, _12350_);
  nor (_12352_, _12351_, _12305_);
  nor (_12353_, _12352_, _06311_);
  or (_12354_, _12353_, _06309_);
  or (_12355_, _12354_, _12304_);
  and (_12356_, _06309_, _04563_);
  nor (_12357_, _12356_, _04779_);
  and (_12358_, _12357_, _12355_);
  and (_12359_, _04779_, _06467_);
  or (_12360_, _12359_, _03401_);
  or (_12361_, _12360_, _12358_);
  and (_12362_, _03401_, \oc8051_golden_model_1.PC [1]);
  nor (_12363_, _12362_, _04791_);
  and (_12364_, _12363_, _12361_);
  and (_12365_, _05669_, _04595_);
  nor (_12366_, _12365_, _12244_);
  nor (_12367_, _12366_, _04793_);
  nor (_12368_, _12367_, _04794_);
  or (_12369_, _12368_, _12364_);
  or (_12370_, _08752_, _06553_);
  and (_12371_, _12370_, _04789_);
  and (_12372_, _12371_, _12369_);
  or (_12373_, _12372_, _12245_);
  and (_12374_, _12373_, _04787_);
  and (_12375_, _08750_, _04786_);
  or (_12376_, _12375_, _03388_);
  or (_12377_, _12376_, _12374_);
  and (_12378_, _03388_, \oc8051_golden_model_1.PC [1]);
  nor (_12379_, _12378_, _06568_);
  and (_12380_, _12379_, _12377_);
  nor (_12381_, _12365_, _06574_);
  or (_12382_, _12381_, _06573_);
  or (_12383_, _12382_, _12380_);
  nand (_12384_, _08751_, _06573_);
  and (_12385_, _12384_, _03384_);
  and (_12386_, _12385_, _12383_);
  and (_12387_, _03383_, _03087_);
  or (_12388_, _04200_, _12387_);
  or (_12389_, _12388_, _12386_);
  nand (_12390_, _12254_, _04200_);
  nor (_12391_, _04632_, _04196_);
  and (_12392_, _12391_, _12390_);
  and (_12393_, _12392_, _12389_);
  nor (_12394_, _12391_, _12254_);
  or (_12395_, _12394_, _05053_);
  or (_12396_, _12395_, _12393_);
  and (_12397_, _04760_, _03244_);
  not (_12398_, _12397_);
  nand (_12399_, _12254_, _05053_);
  and (_12400_, _12399_, _12398_);
  and (_12401_, _12400_, _12396_);
  or (_12402_, _06963_, _06734_);
  or (_12403_, _12402_, _03275_);
  and (_12404_, _12403_, _04812_);
  or (_12405_, _12404_, _12401_);
  not (_12406_, _04471_);
  or (_12407_, _12402_, _12406_);
  and (_12408_, _12407_, _06595_);
  and (_12409_, _12408_, _12405_);
  nor (_12410_, _12262_, _06595_);
  or (_12411_, _12410_, _03899_);
  or (_12412_, _12411_, _12409_);
  and (_12413_, _12412_, _12243_);
  and (_12414_, _03414_, _03087_);
  or (_12415_, _03681_, _12414_);
  or (_12416_, _12415_, _12413_);
  and (_12417_, _03724_, _03412_);
  not (_12418_, _12417_);
  or (_12419_, _12252_, _03682_);
  and (_12420_, _12419_, _12418_);
  and (_12421_, _12420_, _12416_);
  and (_12422_, _12254_, _12417_);
  or (_12423_, _12422_, _04629_);
  or (_12424_, _12423_, _12421_);
  and (_12425_, _04485_, _03307_);
  not (_12426_, _12254_);
  and (_12427_, _12426_, _04485_);
  nor (_12428_, _12427_, _12425_);
  and (_12429_, _12428_, _12424_);
  and (_12430_, _12254_, _12425_);
  or (_12431_, _12430_, _04826_);
  or (_12432_, _12431_, _12429_);
  and (_12433_, _12432_, _12241_);
  or (_12434_, _12433_, _04831_);
  or (_12435_, _12262_, _06960_);
  and (_12436_, _12435_, _05071_);
  and (_12437_, _12436_, _12434_);
  or (_12438_, _12437_, _12055_);
  and (_12439_, _12438_, _12239_);
  nand (_12440_, _10129_, _03899_);
  or (_12441_, _10297_, _03899_);
  and (_12442_, _12441_, _12440_);
  and (_12443_, _12442_, _05400_);
  and (_12444_, _12443_, _12232_);
  or (_40727_, _12444_, _12439_);
  or (_12445_, _12044_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_12446_, _12445_, _12053_);
  nor (_12447_, _05411_, _04989_);
  nor (_12448_, _12447_, _05408_);
  nor (_12449_, _05411_, _05385_);
  nor (_12450_, _12449_, _05412_);
  and (_12451_, _12450_, _05407_);
  nand (_12452_, _12451_, _12448_);
  nor (_12453_, _06963_, _06965_);
  nor (_12454_, _12453_, _08279_);
  or (_12455_, _12454_, _04827_);
  and (_12456_, _06734_, _06824_);
  nor (_12457_, _06734_, _06824_);
  or (_12458_, _12457_, _12456_);
  and (_12459_, _12458_, _12397_);
  nor (_12460_, _05764_, _04180_);
  and (_12461_, _12460_, _04788_);
  or (_12462_, _05307_, _03735_);
  not (_12463_, _10739_);
  nand (_12464_, _10738_, _10736_);
  and (_12465_, _12464_, _03755_);
  and (_12466_, _12465_, _12463_);
  nor (_12467_, _10737_, _10736_);
  or (_12468_, _12467_, _05005_);
  and (_12469_, _06153_, _05764_);
  nor (_12470_, _06153_, _05764_);
  nor (_12471_, _12470_, _12469_);
  nand (_12472_, _12471_, _04723_);
  not (_12473_, _05307_);
  and (_12474_, _06125_, _12473_);
  nor (_12475_, _06125_, _12473_);
  nor (_12476_, _12475_, _12474_);
  nor (_12477_, _12476_, _04266_);
  and (_12478_, _03768_, _03510_);
  nor (_12479_, _03768_, _07190_);
  or (_12480_, _12479_, _12478_);
  and (_12481_, _12480_, _04266_);
  or (_12482_, _12481_, _04723_);
  or (_12483_, _12482_, _12477_);
  and (_12484_, _12483_, _05152_);
  and (_12485_, _12484_, _12472_);
  and (_12486_, _12464_, _04721_);
  or (_12487_, _12486_, _05045_);
  or (_12488_, _12487_, _12485_);
  nor (_12489_, _03510_, _03431_);
  nor (_12490_, _12489_, _04734_);
  and (_12491_, _12490_, _12488_);
  and (_12492_, _05307_, _04734_);
  or (_12493_, _12492_, _04743_);
  or (_12494_, _12493_, _12491_);
  and (_12495_, _12494_, _12468_);
  or (_12496_, _12495_, _03758_);
  nand (_12497_, _05764_, _03758_);
  and (_12498_, _12497_, _03756_);
  and (_12499_, _12498_, _12496_);
  or (_12500_, _12499_, _12466_);
  and (_12501_, _12500_, _03428_);
  or (_12502_, _03511_, _03428_);
  nand (_12503_, _03840_, _12502_);
  or (_12504_, _12503_, _12501_);
  nand (_12505_, _05764_, _03841_);
  and (_12506_, _12505_, _12504_);
  or (_12507_, _12506_, _05131_);
  and (_12508_, _06965_, _05421_);
  nand (_12509_, _05761_, _04939_);
  or (_12510_, _12509_, _12508_);
  and (_12511_, _12510_, _12507_);
  or (_12512_, _12511_, _04759_);
  and (_12513_, _10737_, \oc8051_golden_model_1.PSW [7]);
  nor (_12514_, _12513_, _12467_);
  nand (_12515_, _12514_, _04759_);
  and (_12516_, _12515_, _06141_);
  and (_12517_, _12516_, _12512_);
  nand (_12518_, _03510_, _03456_);
  nand (_12519_, _03735_, _12518_);
  or (_12520_, _12519_, _12517_);
  and (_12521_, _12520_, _12462_);
  or (_12522_, _12521_, _03739_);
  or (_12523_, _06965_, _06305_);
  and (_12524_, _12523_, _06304_);
  and (_12525_, _12524_, _12522_);
  and (_12526_, _06342_, _05307_);
  and (_12527_, _06477_, \oc8051_golden_model_1.DPH [2]);
  and (_12528_, _06483_, \oc8051_golden_model_1.TH1 [2]);
  nor (_12529_, _12528_, _12527_);
  and (_12530_, _06515_, \oc8051_golden_model_1.P2INREG [2]);
  not (_12531_, _12530_);
  and (_12532_, _06512_, \oc8051_golden_model_1.TMOD [2]);
  and (_12533_, _06472_, \oc8051_golden_model_1.TL0 [2]);
  nor (_12534_, _12533_, _12532_);
  and (_12535_, _12534_, _12531_);
  and (_12536_, _06522_, \oc8051_golden_model_1.IE [2]);
  not (_12537_, _12536_);
  and (_12538_, _06525_, \oc8051_golden_model_1.SCON [2]);
  and (_12539_, _06527_, \oc8051_golden_model_1.SBUF [2]);
  nor (_12540_, _12539_, _12538_);
  and (_12541_, _12540_, _12537_);
  and (_12542_, _06501_, \oc8051_golden_model_1.P0INREG [2]);
  not (_12543_, _12542_);
  and (_12544_, _06505_, \oc8051_golden_model_1.P1INREG [2]);
  and (_12545_, _06507_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_12546_, _12545_, _12544_);
  and (_12547_, _12546_, _12543_);
  and (_12548_, _12547_, _12541_);
  and (_12549_, _12548_, _12535_);
  and (_12550_, _12549_, _12529_);
  and (_12551_, _06488_, \oc8051_golden_model_1.TH0 [2]);
  and (_12552_, _06490_, \oc8051_golden_model_1.TL1 [2]);
  nor (_12553_, _12552_, _12551_);
  and (_12554_, _06493_, \oc8051_golden_model_1.TCON [2]);
  and (_12555_, _06497_, \oc8051_golden_model_1.PCON [2]);
  nor (_12556_, _12555_, _12554_);
  and (_12557_, _12556_, _12553_);
  and (_12558_, _06453_, \oc8051_golden_model_1.ACC [2]);
  and (_12559_, _06460_, \oc8051_golden_model_1.B [2]);
  nor (_12560_, _12559_, _12558_);
  and (_12561_, _06445_, \oc8051_golden_model_1.IP [2]);
  and (_12562_, _06458_, \oc8051_golden_model_1.PSW [2]);
  nor (_12563_, _12562_, _12561_);
  and (_12564_, _12563_, _12560_);
  and (_12565_, _06519_, \oc8051_golden_model_1.SP [2]);
  and (_12566_, _06469_, \oc8051_golden_model_1.DPL [2]);
  nor (_12567_, _12566_, _12565_);
  and (_12568_, _12567_, _12564_);
  and (_12569_, _12568_, _12557_);
  and (_12570_, _12569_, _12550_);
  not (_12571_, _12570_);
  nor (_12572_, _12571_, _12526_);
  nor (_12573_, _12572_, _06311_);
  or (_12574_, _12573_, _06309_);
  or (_12575_, _12574_, _12525_);
  and (_12576_, _06309_, _04139_);
  nor (_12577_, _12576_, _04779_);
  and (_12578_, _12577_, _12575_);
  and (_12579_, _04779_, _06495_);
  or (_12580_, _12579_, _03401_);
  or (_12581_, _12580_, _12578_);
  and (_12582_, _03511_, _03401_);
  nor (_12583_, _12582_, _04791_);
  and (_12584_, _12583_, _12581_);
  and (_12585_, _05764_, _04180_);
  nor (_12586_, _12585_, _12460_);
  nor (_12587_, _12586_, _04793_);
  nor (_12588_, _12587_, _04794_);
  or (_12589_, _12588_, _12584_);
  or (_12590_, _08748_, _06553_);
  and (_12591_, _12590_, _04789_);
  and (_12592_, _12591_, _12589_);
  or (_12593_, _12592_, _12461_);
  and (_12594_, _12593_, _04787_);
  and (_12595_, _08746_, _04786_);
  or (_12596_, _12595_, _03388_);
  or (_12597_, _12596_, _12594_);
  and (_12598_, _03511_, _03388_);
  nor (_12599_, _12598_, _06568_);
  and (_12600_, _12599_, _12597_);
  nor (_12601_, _12585_, _06574_);
  or (_12602_, _12601_, _06573_);
  or (_12603_, _12602_, _12600_);
  nand (_12604_, _08747_, _06573_);
  and (_12605_, _12604_, _03384_);
  and (_12606_, _12605_, _12603_);
  or (_12607_, _03732_, _03719_);
  and (_12608_, _12607_, _03244_);
  nand (_12609_, _03510_, _03383_);
  nand (_12610_, _06585_, _12609_);
  or (_12611_, _12610_, _12608_);
  or (_12612_, _12611_, _12606_);
  not (_12613_, _10935_);
  nand (_12614_, _12476_, _12613_);
  and (_12615_, _12614_, _12398_);
  and (_12616_, _12615_, _12612_);
  or (_12617_, _12616_, _12459_);
  and (_12618_, _12617_, _12406_);
  and (_12619_, _12458_, _04471_);
  or (_12620_, _12619_, _12618_);
  and (_12621_, _12620_, _06595_);
  nor (_12622_, _12471_, _06595_);
  or (_12623_, _12622_, _03899_);
  or (_12624_, _12623_, _12621_);
  nand (_12625_, _10160_, _03899_);
  and (_12626_, _12625_, _10953_);
  and (_12627_, _12626_, _12624_);
  and (_12628_, _03510_, _03414_);
  or (_12629_, _03681_, _12628_);
  or (_12630_, _12629_, _12627_);
  or (_12631_, _12467_, _03682_);
  and (_12632_, _12631_, _04482_);
  and (_12633_, _12632_, _12630_);
  nor (_12634_, _06945_, _05307_);
  nor (_12635_, _12634_, _08072_);
  and (_12636_, _12635_, _04483_);
  or (_12637_, _12636_, _04826_);
  or (_12638_, _12637_, _12633_);
  and (_12639_, _12638_, _12455_);
  or (_12640_, _12639_, _04831_);
  nor (_12641_, _05765_, _05717_);
  nor (_12642_, _12641_, _05766_);
  or (_12643_, _12642_, _06960_);
  and (_12644_, _12643_, _05407_);
  and (_12645_, _12644_, _12640_);
  or (_12646_, _12645_, _12452_);
  and (_12647_, _12646_, _12446_);
  nand (_12648_, _10115_, _03899_);
  or (_12649_, _10291_, _03899_);
  and (_12650_, _12649_, _12648_);
  and (_12651_, _12650_, _05400_);
  and (_12652_, _12651_, _12232_);
  or (_40729_, _12652_, _12647_);
  or (_12653_, _12044_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_12655_, _12653_, _12053_);
  nor (_12656_, _08072_, _05119_);
  nor (_12657_, _12656_, _06947_);
  and (_12658_, _12657_, _04827_);
  or (_12659_, _12658_, _05038_);
  nor (_12660_, _12456_, _06779_);
  or (_12661_, _12660_, _06826_);
  and (_12662_, _12661_, _04812_);
  and (_12663_, _03552_, _03383_);
  nor (_12664_, _05621_, _04005_);
  and (_12665_, _12664_, _04788_);
  and (_12666_, _10874_, \oc8051_golden_model_1.PSW [7]);
  nor (_12667_, _10874_, _10873_);
  nor (_12668_, _12667_, _12666_);
  nor (_12669_, _12668_, _05183_);
  and (_12670_, _06964_, _05421_);
  or (_12671_, _12670_, _05619_);
  and (_12672_, _12671_, _04939_);
  not (_12673_, _10876_);
  nand (_12674_, _10875_, _10873_);
  and (_12676_, _12674_, _12673_);
  and (_12677_, _12676_, _03755_);
  or (_12678_, _12667_, _05005_);
  or (_12679_, _12674_, _05152_);
  nor (_12680_, _12469_, _05621_);
  nor (_12681_, _12680_, _06155_);
  nor (_12682_, _12681_, _06250_);
  not (_12683_, _05119_);
  nor (_12684_, _12474_, _12683_);
  or (_12685_, _12684_, _06127_);
  and (_12686_, _12685_, _04267_);
  nor (_12687_, _03768_, _07184_);
  and (_12688_, _03768_, _03552_);
  or (_12689_, _12688_, _12687_);
  and (_12690_, _12689_, _04266_);
  or (_12691_, _12690_, _12686_);
  and (_12692_, _12691_, _06250_);
  or (_12693_, _12692_, _12682_);
  or (_12694_, _12693_, _04721_);
  and (_12695_, _12694_, _12679_);
  or (_12696_, _12695_, _05045_);
  nor (_12697_, _03552_, _03431_);
  nor (_12698_, _12697_, _04734_);
  and (_12699_, _12698_, _12696_);
  and (_12700_, _05119_, _04734_);
  or (_12701_, _12700_, _04743_);
  or (_12702_, _12701_, _12699_);
  and (_12703_, _12702_, _12678_);
  or (_12704_, _12703_, _03758_);
  nand (_12705_, _05621_, _03758_);
  and (_12706_, _12705_, _03756_);
  and (_12707_, _12706_, _12704_);
  or (_12708_, _12707_, _12677_);
  and (_12709_, _12708_, _03428_);
  or (_12710_, _03938_, _03428_);
  nand (_12711_, _03840_, _12710_);
  or (_12712_, _12711_, _12709_);
  nand (_12713_, _05621_, _03841_);
  and (_12714_, _12713_, _04940_);
  and (_12715_, _12714_, _12712_);
  or (_12716_, _12715_, _12672_);
  and (_12717_, _12716_, _05183_);
  or (_12718_, _12717_, _12669_);
  and (_12719_, _12718_, _06141_);
  nand (_12720_, _03552_, _03456_);
  nand (_12721_, _03735_, _12720_);
  or (_12722_, _12721_, _12719_);
  or (_12723_, _05119_, _03735_);
  and (_12724_, _12723_, _12722_);
  or (_12725_, _12724_, _03739_);
  or (_12726_, _06964_, _06305_);
  and (_12727_, _12726_, _06304_);
  and (_12728_, _12727_, _12725_);
  and (_12729_, _06342_, _05119_);
  and (_12730_, _06453_, \oc8051_golden_model_1.ACC [3]);
  and (_12731_, _06460_, \oc8051_golden_model_1.B [3]);
  nor (_12732_, _12731_, _12730_);
  and (_12733_, _06445_, \oc8051_golden_model_1.IP [3]);
  and (_12734_, _06458_, \oc8051_golden_model_1.PSW [3]);
  nor (_12735_, _12734_, _12733_);
  and (_12736_, _12735_, _12732_);
  and (_12737_, _06469_, \oc8051_golden_model_1.DPL [3]);
  and (_12738_, _06472_, \oc8051_golden_model_1.TL0 [3]);
  nor (_12739_, _12738_, _12737_);
  and (_12740_, _06477_, \oc8051_golden_model_1.DPH [3]);
  and (_12741_, _06483_, \oc8051_golden_model_1.TH1 [3]);
  nor (_12742_, _12741_, _12740_);
  and (_12743_, _12742_, _12739_);
  and (_12744_, _12743_, _12736_);
  and (_12745_, _06493_, \oc8051_golden_model_1.TCON [3]);
  and (_12746_, _06488_, \oc8051_golden_model_1.TH0 [3]);
  nor (_12747_, _12746_, _12745_);
  and (_12748_, _06497_, \oc8051_golden_model_1.PCON [3]);
  and (_12749_, _06490_, \oc8051_golden_model_1.TL1 [3]);
  nor (_12750_, _12749_, _12748_);
  and (_12751_, _12750_, _12747_);
  and (_12752_, _06501_, \oc8051_golden_model_1.P0INREG [3]);
  not (_12753_, _12752_);
  and (_12754_, _06505_, \oc8051_golden_model_1.P1INREG [3]);
  and (_12755_, _06507_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_12756_, _12755_, _12754_);
  and (_12757_, _12756_, _12753_);
  and (_12758_, _06512_, \oc8051_golden_model_1.TMOD [3]);
  and (_12759_, _06515_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_12760_, _12759_, _12758_);
  and (_12761_, _12760_, _12757_);
  and (_12762_, _06519_, \oc8051_golden_model_1.SP [3]);
  not (_12763_, _12762_);
  and (_12764_, _06522_, \oc8051_golden_model_1.IE [3]);
  not (_12765_, _12764_);
  and (_12766_, _06525_, \oc8051_golden_model_1.SCON [3]);
  and (_12767_, _06527_, \oc8051_golden_model_1.SBUF [3]);
  nor (_12768_, _12767_, _12766_);
  and (_12769_, _12768_, _12765_);
  and (_12770_, _12769_, _12763_);
  and (_12771_, _12770_, _12761_);
  and (_12772_, _12771_, _12751_);
  and (_12773_, _12772_, _12744_);
  not (_12774_, _12773_);
  nor (_12775_, _12774_, _12729_);
  nor (_12776_, _12775_, _06311_);
  or (_12777_, _12776_, _06309_);
  or (_12778_, _12777_, _12728_);
  and (_12779_, _06309_, _03678_);
  nor (_12780_, _12779_, _04779_);
  and (_12781_, _12780_, _12778_);
  and (_12782_, _04779_, _06345_);
  or (_12783_, _12782_, _03401_);
  or (_12784_, _12783_, _12781_);
  and (_12785_, _03938_, _03401_);
  nor (_12786_, _12785_, _04791_);
  and (_12787_, _12786_, _12784_);
  and (_12788_, _05621_, _04005_);
  nor (_12789_, _12788_, _12664_);
  nor (_12790_, _12789_, _04793_);
  nor (_12791_, _12790_, _04794_);
  or (_12792_, _12791_, _12787_);
  or (_12793_, _10491_, _06553_);
  and (_12794_, _12793_, _04789_);
  and (_12795_, _12794_, _12792_);
  or (_12796_, _12795_, _12665_);
  and (_12797_, _12796_, _04787_);
  and (_12798_, _08744_, _04786_);
  or (_12799_, _12798_, _03388_);
  or (_12800_, _12799_, _12797_);
  and (_12801_, _03938_, _03388_);
  nor (_12802_, _12801_, _06568_);
  and (_12803_, _12802_, _12800_);
  nor (_12804_, _12788_, _06574_);
  or (_12805_, _12804_, _06573_);
  or (_12806_, _12805_, _12803_);
  nand (_12807_, _08742_, _06573_);
  and (_12808_, _12807_, _03384_);
  and (_12809_, _12808_, _12806_);
  nor (_12810_, _12809_, _12663_);
  nor (_12811_, _12810_, _10933_);
  and (_12812_, _12685_, _10933_);
  or (_12813_, _12812_, _10934_);
  or (_12814_, _12813_, _12811_);
  not (_12815_, _10934_);
  or (_12816_, _12685_, _12815_);
  and (_12817_, _12816_, _04813_);
  and (_12818_, _12817_, _12814_);
  or (_12819_, _12818_, _12662_);
  and (_12820_, _12819_, _06595_);
  nor (_12821_, _12681_, _06595_);
  or (_12822_, _12821_, _03899_);
  or (_12823_, _12822_, _12820_);
  nand (_12824_, _10155_, _03899_);
  and (_12825_, _12824_, _10953_);
  and (_12826_, _12825_, _12823_);
  and (_12827_, _03552_, _03414_);
  or (_12828_, _03681_, _12827_);
  or (_12829_, _12828_, _12826_);
  or (_12830_, _12667_, _03682_);
  and (_12831_, _03834_, _03412_);
  and (_12832_, _08115_, _03412_);
  nor (_12833_, _12832_, _12831_);
  nand (_12834_, _12833_, _12418_);
  not (_12835_, _12834_);
  and (_12836_, _12835_, _12830_);
  and (_12837_, _12836_, _12829_);
  and (_12838_, _12834_, _12657_);
  or (_12839_, _12838_, _12837_);
  or (_12840_, _12839_, _05037_);
  and (_12841_, _12840_, _12659_);
  or (_12842_, _08279_, _06964_);
  nor (_12843_, _06967_, _04827_);
  and (_12844_, _12843_, _12842_);
  or (_12845_, _12844_, _04831_);
  or (_12846_, _12845_, _12841_);
  nor (_12847_, _05766_, _05622_);
  nor (_12848_, _12847_, _05767_);
  or (_12849_, _12848_, _06960_);
  and (_12850_, _12849_, _05071_);
  and (_12851_, _12850_, _12846_);
  or (_12852_, _12851_, _12055_);
  and (_12853_, _12852_, _12655_);
  nand (_12854_, _10120_, _03899_);
  or (_12855_, _10286_, _03899_);
  and (_12856_, _12855_, _12854_);
  and (_12857_, _12856_, _05400_);
  and (_12858_, _12857_, _12232_);
  or (_40730_, _12858_, _12853_);
  or (_12859_, _12044_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_12860_, _12859_, _12053_);
  nor (_12861_, _06967_, _06969_);
  nor (_12862_, _12861_, _08261_);
  or (_12863_, _12862_, _04827_);
  not (_12864_, _05950_);
  nor (_12865_, _06127_, _12864_);
  and (_12866_, _06127_, _12864_);
  or (_12867_, _12866_, _12865_);
  or (_12868_, _12867_, _06587_);
  or (_12869_, _08739_, _04787_);
  nor (_12870_, _10791_, _10790_);
  and (_12871_, _10791_, \oc8051_golden_model_1.PSW [7]);
  nor (_12872_, _12871_, _12870_);
  nor (_12873_, _12872_, _05183_);
  not (_12874_, _10793_);
  nand (_12875_, _10792_, _10790_);
  and (_12876_, _12875_, _12874_);
  and (_12877_, _12876_, _03755_);
  or (_12878_, _12870_, _05005_);
  nor (_12879_, _03768_, _07090_);
  and (_12880_, _10317_, _03768_);
  or (_12881_, _12880_, _12879_);
  and (_12882_, _12881_, _04266_);
  and (_12883_, _12867_, _04267_);
  or (_12884_, _12883_, _12882_);
  and (_12885_, _12884_, _04717_);
  and (_12886_, _06969_, _04716_);
  or (_12887_, _12886_, _12885_);
  and (_12888_, _12887_, _06250_);
  nor (_12889_, _06155_, _05953_);
  and (_12890_, _06155_, _05953_);
  nor (_12891_, _12890_, _12889_);
  nor (_12892_, _12891_, _06250_);
  or (_12893_, _12892_, _12888_);
  and (_12894_, _12893_, _05152_);
  and (_12895_, _12875_, _04721_);
  or (_12896_, _12895_, _05045_);
  or (_12897_, _12896_, _12894_);
  nor (_12898_, _10317_, _03431_);
  nor (_12899_, _12898_, _04734_);
  and (_12900_, _12899_, _12897_);
  and (_12901_, _05950_, _04734_);
  or (_12902_, _12901_, _04743_);
  or (_12903_, _12902_, _12900_);
  and (_12904_, _12903_, _12878_);
  or (_12905_, _12904_, _03758_);
  nand (_12906_, _05953_, _03758_);
  and (_12907_, _12906_, _03756_);
  and (_12908_, _12907_, _12905_);
  or (_12909_, _12908_, _12877_);
  and (_12910_, _12909_, _03428_);
  or (_12911_, _10318_, _03428_);
  nand (_12912_, _12911_, _03840_);
  or (_12913_, _12912_, _12910_);
  nand (_12914_, _05953_, _03841_);
  and (_12915_, _12914_, _12913_);
  or (_12916_, _12915_, _05131_);
  and (_12917_, _06969_, _05421_);
  nand (_12918_, _05903_, _04939_);
  or (_12919_, _12918_, _12917_);
  and (_12920_, _12919_, _05183_);
  and (_12921_, _12920_, _12916_);
  or (_12922_, _12921_, _12873_);
  and (_12923_, _12922_, _06141_);
  nand (_12924_, _10317_, _03456_);
  nand (_12925_, _12924_, _03735_);
  or (_12926_, _12925_, _12923_);
  or (_12927_, _05950_, _03735_);
  and (_12928_, _12927_, _12926_);
  or (_12929_, _12928_, _03739_);
  nand (_12930_, _03721_, _03736_);
  or (_12931_, _06969_, _12930_);
  and (_12932_, _12931_, _06311_);
  and (_12933_, _12932_, _12929_);
  and (_12934_, _06342_, _05950_);
  and (_12935_, _06477_, \oc8051_golden_model_1.DPH [4]);
  and (_12936_, _06483_, \oc8051_golden_model_1.TH1 [4]);
  nor (_12937_, _12936_, _12935_);
  and (_12938_, _06453_, \oc8051_golden_model_1.ACC [4]);
  and (_12939_, _06460_, \oc8051_golden_model_1.B [4]);
  nor (_12940_, _12939_, _12938_);
  and (_12941_, _06445_, \oc8051_golden_model_1.IP [4]);
  and (_12942_, _06458_, \oc8051_golden_model_1.PSW [4]);
  nor (_12943_, _12942_, _12941_);
  and (_12944_, _12943_, _12940_);
  and (_12945_, _06515_, \oc8051_golden_model_1.P2INREG [4]);
  not (_12946_, _12945_);
  and (_12947_, _06512_, \oc8051_golden_model_1.TMOD [4]);
  and (_12948_, _06472_, \oc8051_golden_model_1.TL0 [4]);
  nor (_12949_, _12948_, _12947_);
  and (_12950_, _12949_, _12946_);
  and (_12951_, _12950_, _12944_);
  and (_12952_, _12951_, _12937_);
  and (_12953_, _06493_, \oc8051_golden_model_1.TCON [4]);
  and (_12954_, _06488_, \oc8051_golden_model_1.TH0 [4]);
  nor (_12955_, _12954_, _12953_);
  and (_12956_, _06497_, \oc8051_golden_model_1.PCON [4]);
  and (_12957_, _06490_, \oc8051_golden_model_1.TL1 [4]);
  nor (_12958_, _12957_, _12956_);
  and (_12959_, _12958_, _12955_);
  and (_12960_, _06469_, \oc8051_golden_model_1.DPL [4]);
  not (_12961_, _12960_);
  and (_12962_, _06501_, \oc8051_golden_model_1.P0INREG [4]);
  not (_12963_, _12962_);
  and (_12964_, _06505_, \oc8051_golden_model_1.P1INREG [4]);
  and (_12965_, _06507_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_12966_, _12965_, _12964_);
  and (_12967_, _12966_, _12963_);
  and (_12968_, _12967_, _12961_);
  and (_12969_, _06519_, \oc8051_golden_model_1.SP [4]);
  not (_12970_, _12969_);
  and (_12971_, _06522_, \oc8051_golden_model_1.IE [4]);
  not (_12972_, _12971_);
  and (_12973_, _06525_, \oc8051_golden_model_1.SCON [4]);
  and (_12974_, _06527_, \oc8051_golden_model_1.SBUF [4]);
  nor (_12975_, _12974_, _12973_);
  and (_12976_, _12975_, _12972_);
  and (_12977_, _12976_, _12970_);
  and (_12978_, _12977_, _12968_);
  and (_12979_, _12978_, _12959_);
  and (_12980_, _12979_, _12952_);
  not (_12981_, _12980_);
  nor (_12982_, _12981_, _12934_);
  nor (_12983_, _12982_, _06311_);
  or (_12984_, _12983_, _06309_);
  or (_12985_, _12984_, _12933_);
  and (_12986_, _06309_, _04526_);
  nor (_12987_, _12986_, _04779_);
  and (_12988_, _12987_, _12985_);
  and (_12989_, _06456_, _04779_);
  or (_12990_, _12989_, _03401_);
  or (_12991_, _12990_, _12988_);
  and (_12992_, _10318_, _03401_);
  nor (_12993_, _12992_, _04791_);
  and (_12994_, _12993_, _12991_);
  nor (_12995_, _06442_, _05953_);
  and (_12996_, _06442_, _05953_);
  nor (_12997_, _12996_, _12995_);
  and (_12998_, _12997_, _04791_);
  or (_12999_, _12998_, _04793_);
  or (_13000_, _12999_, _12994_);
  or (_13001_, _08741_, _06553_);
  and (_13002_, _13001_, _04789_);
  and (_13003_, _13002_, _13000_);
  and (_13004_, _12995_, _04788_);
  or (_13005_, _13004_, _04786_);
  or (_13006_, _13005_, _13003_);
  and (_13007_, _13006_, _12869_);
  or (_13008_, _13007_, _03388_);
  and (_13009_, _10318_, _03388_);
  nor (_13010_, _13009_, _06568_);
  and (_13011_, _13010_, _13008_);
  nor (_13012_, _12996_, _06574_);
  or (_13013_, _13012_, _06573_);
  or (_13014_, _13013_, _13011_);
  nand (_13015_, _08740_, _06573_);
  and (_13016_, _13015_, _03384_);
  and (_13017_, _13016_, _13014_);
  nand (_13018_, _10317_, _03383_);
  nand (_13019_, _13018_, _06587_);
  or (_13020_, _13019_, _13017_);
  and (_13021_, _13020_, _12868_);
  or (_13022_, _13021_, _05053_);
  or (_13023_, _12867_, _06590_);
  and (_13024_, _13023_, _12398_);
  and (_13025_, _13024_, _13022_);
  and (_13026_, _06826_, _06918_);
  nor (_13027_, _06826_, _06918_);
  or (_13028_, _13027_, _13026_);
  or (_13029_, _13028_, _03275_);
  and (_13030_, _13029_, _04812_);
  or (_13031_, _13030_, _13025_);
  or (_13032_, _13028_, _12406_);
  and (_13033_, _13032_, _06595_);
  and (_13034_, _13033_, _13031_);
  nor (_13035_, _12891_, _06595_);
  or (_13036_, _13035_, _03899_);
  or (_13037_, _13036_, _13034_);
  nand (_13038_, _10150_, _03899_);
  and (_13039_, _13038_, _10953_);
  and (_13040_, _13039_, _13037_);
  and (_13041_, _10317_, _03414_);
  or (_13042_, _13041_, _03681_);
  or (_13043_, _13042_, _13040_);
  or (_13044_, _12870_, _03682_);
  and (_13045_, _13044_, _04482_);
  and (_13046_, _13045_, _13043_);
  nor (_13047_, _06947_, _05950_);
  nor (_13048_, _13047_, _08055_);
  and (_13049_, _13048_, _04483_);
  or (_13050_, _13049_, _04826_);
  or (_13051_, _13050_, _13046_);
  and (_13052_, _13051_, _12863_);
  or (_13053_, _13052_, _04831_);
  and (_13054_, _08336_, _05767_);
  nor (_13055_, _08336_, _05767_);
  nor (_13056_, _13055_, _13054_);
  or (_13057_, _13056_, _06960_);
  and (_13058_, _13057_, _05071_);
  and (_13059_, _13058_, _13053_);
  or (_13060_, _13059_, _12055_);
  and (_13061_, _13060_, _12860_);
  nand (_13062_, _10111_, _03899_);
  or (_13063_, _10283_, _03899_);
  and (_13064_, _13063_, _13062_);
  and (_13065_, _13064_, _05400_);
  and (_13066_, _13065_, _12232_);
  or (_40731_, _13066_, _13061_);
  or (_13067_, _12044_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_13068_, _13067_, _12053_);
  nor (_13069_, _06411_, _05859_);
  and (_13070_, _13069_, _04788_);
  nor (_13071_, _10901_, _10900_);
  and (_13072_, _10901_, \oc8051_golden_model_1.PSW [7]);
  nor (_13073_, _13072_, _13071_);
  nor (_13074_, _13073_, _05183_);
  or (_13075_, _13071_, _05005_);
  nor (_13076_, _03768_, _07084_);
  and (_13077_, _10312_, _03768_);
  or (_13078_, _13077_, _13076_);
  and (_13079_, _13078_, _04266_);
  not (_13080_, _05857_);
  nor (_13081_, _12866_, _13080_);
  or (_13082_, _13081_, _06128_);
  and (_13083_, _13082_, _04267_);
  or (_13084_, _13083_, _13079_);
  and (_13085_, _13084_, _04717_);
  and (_13086_, _06968_, _04716_);
  or (_13087_, _13086_, _13085_);
  and (_13088_, _13087_, _06250_);
  nor (_13089_, _12890_, _05859_);
  nor (_13090_, _13089_, _06156_);
  nor (_13091_, _13090_, _06250_);
  or (_13092_, _13091_, _13088_);
  and (_13093_, _13092_, _05152_);
  nand (_13094_, _10902_, _10900_);
  and (_13095_, _13094_, _04721_);
  or (_13096_, _13095_, _05045_);
  or (_13097_, _13096_, _13093_);
  nor (_13098_, _10312_, _03431_);
  nor (_13099_, _13098_, _04734_);
  and (_13100_, _13099_, _13097_);
  and (_13101_, _05857_, _04734_);
  or (_13102_, _13101_, _04743_);
  or (_13103_, _13102_, _13100_);
  and (_13104_, _13103_, _13075_);
  or (_13105_, _13104_, _03758_);
  nand (_13106_, _05859_, _03758_);
  and (_13107_, _13106_, _03756_);
  and (_13108_, _13107_, _13105_);
  not (_13109_, _10903_);
  and (_13110_, _13094_, _13109_);
  and (_13111_, _13110_, _03755_);
  or (_13112_, _13111_, _13108_);
  and (_13113_, _13112_, _03428_);
  or (_13114_, _10313_, _03428_);
  nand (_13115_, _13114_, _03840_);
  or (_13116_, _13115_, _13113_);
  nand (_13117_, _05859_, _03841_);
  and (_13118_, _13117_, _13116_);
  or (_13119_, _13118_, _05131_);
  and (_13120_, _06968_, _05421_);
  nand (_13121_, _05811_, _05131_);
  or (_13122_, _13121_, _13120_);
  and (_13123_, _13122_, _05183_);
  and (_13124_, _13123_, _13119_);
  or (_13125_, _13124_, _13074_);
  and (_13126_, _13125_, _06141_);
  nand (_13127_, _10312_, _03456_);
  nand (_13128_, _13127_, _03735_);
  or (_13129_, _13128_, _13126_);
  or (_13130_, _05857_, _03735_);
  and (_13131_, _13130_, _13129_);
  or (_13132_, _13131_, _03739_);
  or (_13133_, _06968_, _06305_);
  and (_13134_, _13133_, _06304_);
  and (_13135_, _13134_, _13132_);
  and (_13136_, _06342_, _05857_);
  and (_13137_, _06477_, \oc8051_golden_model_1.DPH [5]);
  and (_13138_, _06483_, \oc8051_golden_model_1.TH1 [5]);
  nor (_13139_, _13138_, _13137_);
  and (_13140_, _06515_, \oc8051_golden_model_1.P2INREG [5]);
  not (_13141_, _13140_);
  and (_13142_, _06512_, \oc8051_golden_model_1.TMOD [5]);
  and (_13143_, _06472_, \oc8051_golden_model_1.TL0 [5]);
  nor (_13144_, _13143_, _13142_);
  and (_13145_, _13144_, _13141_);
  and (_13146_, _06522_, \oc8051_golden_model_1.IE [5]);
  not (_13147_, _13146_);
  and (_13148_, _06525_, \oc8051_golden_model_1.SCON [5]);
  and (_13149_, _06527_, \oc8051_golden_model_1.SBUF [5]);
  nor (_13150_, _13149_, _13148_);
  and (_13151_, _13150_, _13147_);
  and (_13152_, _06501_, \oc8051_golden_model_1.P0INREG [5]);
  not (_13153_, _13152_);
  and (_13154_, _06505_, \oc8051_golden_model_1.P1INREG [5]);
  and (_13155_, _06507_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_13156_, _13155_, _13154_);
  and (_13157_, _13156_, _13153_);
  and (_13158_, _13157_, _13151_);
  and (_13159_, _13158_, _13145_);
  and (_13160_, _13159_, _13139_);
  and (_13161_, _06488_, \oc8051_golden_model_1.TH0 [5]);
  and (_13162_, _06490_, \oc8051_golden_model_1.TL1 [5]);
  nor (_13163_, _13162_, _13161_);
  and (_13164_, _06493_, \oc8051_golden_model_1.TCON [5]);
  and (_13165_, _06497_, \oc8051_golden_model_1.PCON [5]);
  nor (_13166_, _13165_, _13164_);
  and (_13167_, _13166_, _13163_);
  and (_13168_, _06453_, \oc8051_golden_model_1.ACC [5]);
  and (_13169_, _06460_, \oc8051_golden_model_1.B [5]);
  nor (_13170_, _13169_, _13168_);
  and (_13171_, _06445_, \oc8051_golden_model_1.IP [5]);
  and (_13172_, _06458_, \oc8051_golden_model_1.PSW [5]);
  nor (_13173_, _13172_, _13171_);
  and (_13174_, _13173_, _13170_);
  and (_13175_, _06519_, \oc8051_golden_model_1.SP [5]);
  and (_13176_, _06469_, \oc8051_golden_model_1.DPL [5]);
  nor (_13177_, _13176_, _13175_);
  and (_13178_, _13177_, _13174_);
  and (_13179_, _13178_, _13167_);
  and (_13180_, _13179_, _13160_);
  not (_13181_, _13180_);
  nor (_13182_, _13181_, _13136_);
  nor (_13183_, _13182_, _06311_);
  or (_13184_, _13183_, _06309_);
  or (_13185_, _13184_, _13135_);
  and (_13186_, _06309_, _04093_);
  nor (_13187_, _13186_, _04779_);
  and (_13188_, _13187_, _13185_);
  and (_13189_, _06447_, _04779_);
  or (_13190_, _13189_, _03401_);
  or (_13191_, _13190_, _13188_);
  and (_13192_, _10313_, _03401_);
  nor (_13193_, _13192_, _04791_);
  and (_13194_, _13193_, _13191_);
  and (_13195_, _06411_, _05859_);
  nor (_13196_, _13195_, _13069_);
  nor (_13197_, _13196_, _04793_);
  nor (_13198_, _13197_, _04794_);
  or (_13199_, _13198_, _13194_);
  or (_13200_, _10493_, _06553_);
  and (_13201_, _13200_, _04789_);
  and (_13202_, _13201_, _13199_);
  or (_13203_, _13202_, _13070_);
  and (_13204_, _13203_, _04787_);
  and (_13205_, _08737_, _04786_);
  or (_13206_, _13205_, _03388_);
  or (_13207_, _13206_, _13204_);
  and (_13208_, _10313_, _03388_);
  nor (_13209_, _13208_, _06568_);
  and (_13210_, _13209_, _13207_);
  nor (_13211_, _13195_, _06574_);
  or (_13212_, _13211_, _06573_);
  or (_13213_, _13212_, _13210_);
  nand (_13214_, _08738_, _06573_);
  and (_13215_, _13214_, _03384_);
  and (_13216_, _13215_, _13213_);
  and (_13217_, _08115_, _03244_);
  and (_13218_, _10312_, _03383_);
  or (_13219_, _13218_, _13217_);
  or (_13220_, _13219_, _10933_);
  or (_13221_, _13220_, _13216_);
  or (_13222_, _13082_, _10935_);
  and (_13223_, _13222_, _13221_);
  and (_13224_, _13082_, _04472_);
  or (_13225_, _13224_, _04812_);
  or (_13226_, _13225_, _13223_);
  nor (_13227_, _13026_, _06873_);
  or (_13228_, _06920_, _04813_);
  or (_13229_, _13228_, _13227_);
  and (_13230_, _13229_, _06595_);
  and (_13231_, _13230_, _13226_);
  nor (_13232_, _13090_, _06595_);
  or (_13233_, _13232_, _03899_);
  or (_13234_, _13233_, _13231_);
  nand (_13235_, _10145_, _03899_);
  and (_13236_, _13235_, _10953_);
  and (_13237_, _13236_, _13234_);
  and (_13238_, _10312_, _03414_);
  or (_13239_, _13238_, _03681_);
  or (_13240_, _13239_, _13237_);
  or (_13241_, _13071_, _03682_);
  and (_13242_, _13241_, _04482_);
  and (_13243_, _13242_, _13240_);
  or (_13244_, _08055_, _05857_);
  nor (_13245_, _06949_, _04482_);
  and (_13246_, _13245_, _13244_);
  or (_13247_, _13246_, _13243_);
  and (_13248_, _13247_, _04827_);
  or (_13249_, _08261_, _06968_);
  nor (_13250_, _06971_, _04827_);
  and (_13251_, _13250_, _13249_);
  or (_13252_, _13251_, _04831_);
  or (_13253_, _13252_, _13248_);
  nor (_13254_, _13054_, _08335_);
  nor (_13255_, _13254_, _05956_);
  or (_13256_, _13255_, _06960_);
  and (_13257_, _13256_, _05071_);
  and (_13258_, _13257_, _13253_);
  or (_13259_, _13258_, _12055_);
  and (_13260_, _13259_, _13068_);
  nand (_13261_, _10106_, _03899_);
  or (_13262_, _10279_, _03899_);
  and (_13263_, _13262_, _13261_);
  and (_13264_, _13263_, _05400_);
  and (_13265_, _13264_, _12232_);
  or (_40733_, _13265_, _13260_);
  or (_13266_, _12044_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_13267_, _13266_, _12053_);
  nand (_13268_, _06949_, _06065_);
  or (_13269_, _06949_, _06065_);
  and (_13270_, _13269_, _04483_);
  and (_13271_, _13270_, _13268_);
  nor (_13272_, _06128_, _06123_);
  or (_13273_, _13272_, _06129_);
  or (_13274_, _13273_, _06587_);
  nor (_13275_, _06379_, _06068_);
  and (_13276_, _13275_, _04788_);
  nor (_13277_, _10846_, _10845_);
  and (_13278_, _10846_, \oc8051_golden_model_1.PSW [7]);
  nor (_13279_, _13278_, _13277_);
  nor (_13280_, _13279_, _05183_);
  or (_13281_, _13277_, _05005_);
  or (_13282_, _13273_, _04266_);
  nor (_13283_, _03768_, _07036_);
  and (_13284_, _10305_, _03768_);
  or (_13285_, _13284_, _13283_);
  or (_13286_, _13285_, _04267_);
  and (_13287_, _13286_, _13282_);
  or (_13288_, _13287_, _04716_);
  or (_13289_, _06641_, _04717_);
  and (_13290_, _13289_, _13288_);
  and (_13291_, _13290_, _06250_);
  nor (_13292_, _06156_, _06068_);
  nor (_13293_, _13292_, _06157_);
  nor (_13294_, _13293_, _06250_);
  or (_13295_, _13294_, _13291_);
  and (_13296_, _13295_, _05152_);
  nand (_13297_, _10847_, _10845_);
  and (_13298_, _13297_, _04721_);
  or (_13299_, _13298_, _05045_);
  or (_13300_, _13299_, _13296_);
  nor (_13301_, _10305_, _03431_);
  nor (_13302_, _13301_, _04734_);
  and (_13303_, _13302_, _13300_);
  and (_13304_, _06065_, _04734_);
  or (_13305_, _13304_, _04743_);
  or (_13306_, _13305_, _13303_);
  and (_13307_, _13306_, _13281_);
  or (_13308_, _13307_, _03758_);
  nand (_13309_, _06068_, _03758_);
  and (_13310_, _13309_, _03756_);
  and (_13311_, _13310_, _13308_);
  not (_13312_, _10848_);
  and (_13313_, _13297_, _13312_);
  and (_13314_, _13313_, _03755_);
  or (_13315_, _13314_, _13311_);
  and (_13316_, _13315_, _03428_);
  or (_13317_, _10306_, _03428_);
  nand (_13318_, _13317_, _03840_);
  or (_13319_, _13318_, _13316_);
  nand (_13320_, _06068_, _03841_);
  and (_13321_, _13320_, _13319_);
  or (_13322_, _13321_, _05131_);
  and (_13323_, _06641_, _05421_);
  nand (_13324_, _06011_, _04939_);
  or (_13325_, _13324_, _13323_);
  and (_13326_, _13325_, _05183_);
  and (_13327_, _13326_, _13322_);
  or (_13328_, _13327_, _13280_);
  and (_13329_, _13328_, _06141_);
  nand (_13330_, _10305_, _03456_);
  nand (_13331_, _13330_, _03735_);
  or (_13332_, _13331_, _13329_);
  or (_13333_, _06065_, _03735_);
  and (_13334_, _13333_, _13332_);
  or (_13335_, _13334_, _03739_);
  or (_13336_, _06641_, _12930_);
  and (_13337_, _13336_, _06311_);
  and (_13338_, _13337_, _13335_);
  and (_13339_, _06342_, _06065_);
  and (_13340_, _06469_, \oc8051_golden_model_1.DPL [6]);
  not (_13341_, _13340_);
  and (_13342_, _06472_, \oc8051_golden_model_1.TL0 [6]);
  not (_13343_, _13342_);
  and (_13344_, _06505_, \oc8051_golden_model_1.P1INREG [6]);
  and (_13345_, _06507_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_13346_, _13345_, _13344_);
  and (_13347_, _13346_, _13343_);
  and (_13348_, _06501_, \oc8051_golden_model_1.P0INREG [6]);
  and (_13349_, _06515_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_13350_, _13349_, _13348_);
  and (_13351_, _13350_, _13347_);
  and (_13352_, _13351_, _13341_);
  and (_13353_, _06453_, \oc8051_golden_model_1.ACC [6]);
  and (_13354_, _06460_, \oc8051_golden_model_1.B [6]);
  nor (_13355_, _13354_, _13353_);
  and (_13356_, _06445_, \oc8051_golden_model_1.IP [6]);
  and (_13357_, _06458_, \oc8051_golden_model_1.PSW [6]);
  nor (_13358_, _13357_, _13356_);
  and (_13359_, _13358_, _13355_);
  and (_13360_, _06490_, \oc8051_golden_model_1.TL1 [6]);
  and (_13361_, _06488_, \oc8051_golden_model_1.TH0 [6]);
  nor (_13362_, _13361_, _13360_);
  and (_13363_, _13362_, _13359_);
  and (_13364_, _13363_, _13352_);
  and (_13365_, _06512_, \oc8051_golden_model_1.TMOD [6]);
  and (_13366_, _06483_, \oc8051_golden_model_1.TH1 [6]);
  nor (_13367_, _13366_, _13365_);
  and (_13368_, _06519_, \oc8051_golden_model_1.SP [6]);
  and (_13369_, _06477_, \oc8051_golden_model_1.DPH [6]);
  nor (_13370_, _13369_, _13368_);
  and (_13371_, _13370_, _13367_);
  and (_13372_, _06497_, \oc8051_golden_model_1.PCON [6]);
  not (_13373_, _13372_);
  and (_13374_, _06522_, \oc8051_golden_model_1.IE [6]);
  not (_13375_, _13374_);
  and (_13376_, _06493_, \oc8051_golden_model_1.TCON [6]);
  not (_13377_, _13376_);
  and (_13378_, _06525_, \oc8051_golden_model_1.SCON [6]);
  and (_13379_, _06527_, \oc8051_golden_model_1.SBUF [6]);
  nor (_13380_, _13379_, _13378_);
  and (_13381_, _13380_, _13377_);
  and (_13382_, _13381_, _13375_);
  and (_13383_, _13382_, _13373_);
  and (_13384_, _13383_, _13371_);
  and (_13385_, _13384_, _13364_);
  not (_13386_, _13385_);
  nor (_13387_, _13386_, _13339_);
  nor (_13388_, _13387_, _06311_);
  or (_13389_, _13388_, _06309_);
  or (_13390_, _13389_, _13338_);
  and (_13391_, _06309_, _03810_);
  nor (_13392_, _13391_, _04779_);
  and (_13393_, _13392_, _13390_);
  not (_13394_, _06379_);
  and (_13395_, _13394_, _04779_);
  or (_13396_, _13395_, _03401_);
  or (_13397_, _13396_, _13393_);
  and (_13398_, _10306_, _03401_);
  nor (_13399_, _13398_, _04791_);
  and (_13400_, _13399_, _13397_);
  and (_13401_, _06379_, _06068_);
  nor (_13402_, _13401_, _13275_);
  and (_13403_, _13402_, _04791_);
  or (_13404_, _13403_, _04793_);
  or (_13405_, _13404_, _13400_);
  or (_13406_, _08736_, _06553_);
  and (_13407_, _13406_, _04789_);
  and (_13408_, _13407_, _13405_);
  or (_13409_, _13408_, _13276_);
  and (_13410_, _13409_, _04787_);
  and (_13411_, _08734_, _04786_);
  or (_13412_, _13411_, _03388_);
  or (_13413_, _13412_, _13410_);
  and (_13414_, _10306_, _03388_);
  nor (_13415_, _13414_, _06568_);
  and (_13416_, _13415_, _13413_);
  nor (_13417_, _13401_, _06574_);
  or (_13418_, _13417_, _06573_);
  or (_13419_, _13418_, _13416_);
  nand (_13420_, _08735_, _06573_);
  and (_13421_, _13420_, _03384_);
  and (_13422_, _13421_, _13419_);
  nand (_13423_, _10305_, _03383_);
  nand (_13424_, _13423_, _06587_);
  or (_13425_, _13424_, _13422_);
  and (_13426_, _13425_, _13274_);
  or (_13427_, _13426_, _05053_);
  or (_13428_, _13273_, _06590_);
  and (_13429_, _13428_, _12398_);
  and (_13430_, _13429_, _13427_);
  nor (_13431_, _06920_, _06642_);
  or (_13432_, _13431_, _06921_);
  or (_13433_, _13432_, _04471_);
  and (_13434_, _13433_, _04812_);
  or (_13435_, _13434_, _13430_);
  or (_13436_, _13432_, _12406_);
  and (_13437_, _13436_, _06595_);
  and (_13438_, _13437_, _13435_);
  nor (_13439_, _13293_, _06595_);
  or (_13440_, _13439_, _03899_);
  or (_13441_, _13440_, _13438_);
  nand (_13442_, _10138_, _03899_);
  and (_13443_, _13442_, _10953_);
  and (_13444_, _13443_, _13441_);
  and (_13445_, _10305_, _03414_);
  or (_13446_, _13445_, _03681_);
  or (_13447_, _13446_, _13444_);
  or (_13448_, _13277_, _03682_);
  and (_13449_, _13448_, _04482_);
  and (_13450_, _13449_, _13447_);
  or (_13451_, _13450_, _13271_);
  and (_13452_, _13451_, _04827_);
  or (_13453_, _06971_, _06641_);
  nor (_13454_, _06972_, _04827_);
  and (_13455_, _13454_, _13453_);
  or (_13456_, _13455_, _04831_);
  or (_13457_, _13456_, _13452_);
  nor (_13458_, _06068_, _05956_);
  and (_13459_, _06068_, _05956_);
  nor (_13460_, _13459_, _13458_);
  nand (_13461_, _13460_, _04831_);
  and (_13462_, _13461_, _05071_);
  and (_13463_, _13462_, _13457_);
  or (_13464_, _13463_, _12055_);
  and (_13465_, _13464_, _13267_);
  or (_13466_, _10099_, _03900_);
  or (_13467_, _10274_, _03899_);
  and (_13468_, _13467_, _13466_);
  and (_13469_, _13468_, _05400_);
  and (_13470_, _13469_, _12232_);
  or (_40734_, _13470_, _13465_);
  or (_13471_, _12044_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_13472_, _13471_, _12053_);
  or (_13473_, _12055_, _06979_);
  and (_13474_, _13473_, _13472_);
  and (_13475_, _12232_, _07006_);
  or (_40735_, _13475_, _13474_);
  and (_13476_, _05408_, _04989_);
  and (_13477_, _13476_, _12450_);
  or (_13478_, _13477_, \oc8051_golden_model_1.IRAM[1] [0]);
  not (_13479_, _05123_);
  or (_13480_, _12051_, _13479_);
  or (_13481_, _13480_, _12047_);
  and (_13482_, _13481_, _13478_);
  and (_13483_, _12224_, _05407_);
  and (_13484_, _13483_, _12223_);
  not (_13485_, _13477_);
  or (_13486_, _13485_, _13484_);
  and (_13487_, _13486_, _13482_);
  and (_13488_, _05400_, _05123_);
  and (_13489_, _13488_, _12230_);
  and (_13490_, _13489_, _12236_);
  or (_40740_, _13490_, _13487_);
  or (_13491_, _13477_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_13492_, _13491_, _13481_);
  and (_13493_, _12435_, _05407_);
  and (_13494_, _13493_, _12434_);
  or (_13495_, _13485_, _13494_);
  and (_13496_, _13495_, _13492_);
  and (_13497_, _13489_, _12443_);
  or (_40741_, _13497_, _13496_);
  or (_13498_, _13477_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_13499_, _13498_, _13481_);
  or (_13500_, _13485_, _12645_);
  and (_13501_, _13500_, _13499_);
  and (_13502_, _13489_, _12651_);
  or (_40742_, _13502_, _13501_);
  or (_13503_, _13477_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_13504_, _13503_, _13481_);
  and (_13505_, _12849_, _05407_);
  and (_13506_, _13505_, _12846_);
  or (_13507_, _13485_, _13506_);
  and (_13508_, _13507_, _13504_);
  and (_13509_, _13489_, _12857_);
  or (_40743_, _13509_, _13508_);
  or (_13510_, _13477_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_13511_, _13510_, _13481_);
  and (_13512_, _13057_, _05407_);
  and (_13513_, _13512_, _13053_);
  or (_13514_, _13485_, _13513_);
  and (_13515_, _13514_, _13511_);
  and (_13516_, _13489_, _13065_);
  or (_40745_, _13516_, _13515_);
  and (_13517_, _13256_, _05407_);
  and (_13518_, _13517_, _13253_);
  or (_13519_, _13485_, _13518_);
  nor (_13520_, _13477_, \oc8051_golden_model_1.IRAM[1] [5]);
  nor (_13521_, _13520_, _13489_);
  and (_13522_, _13521_, _13519_);
  and (_13523_, _13489_, _13264_);
  or (_40746_, _13523_, _13522_);
  or (_13524_, _13477_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_13525_, _13524_, _13481_);
  and (_13526_, _13461_, _05407_);
  and (_13527_, _13526_, _13457_);
  or (_13528_, _13485_, _13527_);
  and (_13529_, _13528_, _13525_);
  and (_13530_, _13489_, _13469_);
  or (_40747_, _13530_, _13529_);
  or (_13531_, _13477_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_13532_, _13531_, _13481_);
  or (_13533_, _13485_, _06980_);
  and (_13534_, _13533_, _13532_);
  and (_13535_, _13489_, _07006_);
  or (_40748_, _13535_, _13534_);
  not (_13536_, _04834_);
  and (_13537_, _05073_, _13536_);
  and (_13538_, _13537_, _12042_);
  or (_13539_, _13538_, \oc8051_golden_model_1.IRAM[2] [0]);
  not (_13540_, _06162_);
  or (_13541_, _12051_, _13540_);
  or (_13542_, _13541_, _12047_);
  and (_13543_, _13542_, _13539_);
  not (_13544_, _13538_);
  or (_13545_, _13544_, _12226_);
  and (_13546_, _13545_, _13543_);
  and (_13547_, _06162_, _05400_);
  and (_13548_, _13547_, _12230_);
  and (_13549_, _13548_, _12236_);
  or (_40752_, _13549_, _13546_);
  or (_13550_, _13538_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_13551_, _13550_, _13542_);
  or (_13552_, _13544_, _12437_);
  and (_13553_, _13552_, _13551_);
  and (_13554_, _13548_, _12443_);
  or (_40754_, _13554_, _13553_);
  or (_13555_, _13538_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_13556_, _13555_, _13542_);
  and (_13557_, _12447_, _13536_);
  nand (_13558_, _13557_, _12450_);
  or (_13559_, _13558_, _12645_);
  and (_13560_, _13559_, _13556_);
  and (_13561_, _13548_, _12651_);
  or (_40755_, _13561_, _13560_);
  or (_13562_, _13538_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_13563_, _13562_, _13542_);
  or (_13564_, _13544_, _12851_);
  and (_13565_, _13564_, _13563_);
  and (_13566_, _13548_, _12857_);
  or (_40756_, _13566_, _13565_);
  or (_13567_, _13538_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_13568_, _13567_, _13542_);
  or (_13569_, _13544_, _13059_);
  and (_13570_, _13569_, _13568_);
  and (_13571_, _13548_, _13065_);
  or (_40757_, _13571_, _13570_);
  or (_13572_, _13538_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_13573_, _13572_, _13542_);
  or (_13574_, _13544_, _13258_);
  and (_13575_, _13574_, _13573_);
  and (_13576_, _13548_, _13264_);
  or (_40758_, _13576_, _13575_);
  or (_13578_, _13538_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_13579_, _13578_, _13542_);
  or (_13580_, _13544_, _13463_);
  and (_13581_, _13580_, _13579_);
  and (_13582_, _13548_, _13469_);
  or (_40760_, _13582_, _13581_);
  or (_13583_, _13538_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_13584_, _13583_, _13542_);
  or (_13585_, _13558_, _06980_);
  and (_13586_, _13585_, _13584_);
  and (_13588_, _13548_, _07006_);
  or (_40761_, _13588_, _13586_);
  and (_13589_, _12042_, _05074_);
  or (_13590_, _13589_, \oc8051_golden_model_1.IRAM[3] [0]);
  not (_13591_, _04837_);
  or (_13592_, _12051_, _13591_);
  or (_13593_, _13592_, _12047_);
  and (_13594_, _13593_, _13590_);
  not (_13595_, _13589_);
  or (_13596_, _13595_, _12226_);
  and (_13598_, _13596_, _13594_);
  and (_13599_, _05400_, _04837_);
  and (_13600_, _13599_, _12230_);
  and (_13601_, _13600_, _12236_);
  or (_40765_, _13601_, _13598_);
  or (_13602_, _13589_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_13603_, _13602_, _13593_);
  or (_13604_, _13595_, _12437_);
  and (_13605_, _13604_, _13603_);
  and (_13606_, _13600_, _12443_);
  or (_40766_, _13606_, _13605_);
  or (_13608_, _13589_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_13609_, _13608_, _13593_);
  nand (_13610_, _12450_, _05409_);
  or (_13611_, _13610_, _12645_);
  and (_13612_, _13611_, _13609_);
  and (_13613_, _13600_, _12651_);
  or (_40767_, _13613_, _13612_);
  or (_13614_, _13589_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_13615_, _13614_, _13593_);
  or (_13617_, _13595_, _12851_);
  and (_13618_, _13617_, _13615_);
  and (_13619_, _13600_, _12857_);
  or (_40768_, _13619_, _13618_);
  or (_13620_, _13610_, _13513_);
  or (_13621_, _13589_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_13622_, _13621_, _13593_);
  and (_13623_, _13622_, _13620_);
  and (_13624_, _13600_, _13065_);
  or (_40770_, _13624_, _13623_);
  or (_13626_, _13589_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_13627_, _13626_, _13593_);
  or (_13628_, _13595_, _13258_);
  and (_13629_, _13628_, _13627_);
  and (_13630_, _13600_, _13264_);
  or (_40771_, _13630_, _13629_);
  or (_13631_, _13589_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_13632_, _13631_, _13593_);
  or (_13633_, _13595_, _13463_);
  and (_13634_, _13633_, _13632_);
  and (_13636_, _13600_, _13469_);
  or (_40772_, _13636_, _13634_);
  or (_13637_, _13589_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_13638_, _13637_, _13593_);
  or (_13639_, _13610_, _06980_);
  and (_13640_, _13639_, _13638_);
  and (_13641_, _13600_, _07006_);
  or (_40773_, _13641_, _13640_);
  and (_13642_, _05386_, _05242_);
  and (_13643_, _13642_, _12040_);
  nor (_13645_, _13643_, _04666_);
  and (_13646_, _13643_, _12226_);
  or (_13647_, _13646_, _13645_);
  not (_13648_, _05396_);
  and (_13649_, _12229_, _13648_);
  and (_13650_, _13649_, _04838_);
  or (_13651_, _13650_, _13647_);
  not (_13652_, _13650_);
  or (_13653_, _13652_, _12236_);
  and (_40777_, _13653_, _13651_);
  not (_13655_, _13643_);
  or (_13656_, _13655_, _12437_);
  and (_13657_, _12049_, _13648_);
  nand (_13658_, _13657_, _04838_);
  or (_13659_, _13643_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_13660_, _13659_, _13658_);
  and (_13661_, _13660_, _13656_);
  and (_13662_, _13650_, _12443_);
  or (_40779_, _13662_, _13661_);
  or (_13663_, _13655_, _12645_);
  or (_13665_, _13643_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_13666_, _13665_, _13658_);
  and (_13667_, _13666_, _13663_);
  and (_13668_, _13650_, _12651_);
  or (_40780_, _13668_, _13667_);
  or (_13669_, _13655_, _12851_);
  or (_13670_, _13643_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_13671_, _13670_, _13658_);
  and (_13672_, _13671_, _13669_);
  and (_13673_, _13650_, _12857_);
  or (_40781_, _13673_, _13672_);
  or (_13675_, _13655_, _13059_);
  or (_13676_, _13643_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_13677_, _13676_, _13658_);
  and (_13678_, _13677_, _13675_);
  and (_13679_, _13650_, _13065_);
  or (_40782_, _13679_, _13678_);
  or (_13680_, _13655_, _13518_);
  or (_13681_, _13643_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_13682_, _13681_, _13652_);
  and (_13684_, _13682_, _13680_);
  and (_13685_, _13650_, _13264_);
  or (_40783_, _13685_, _13684_);
  or (_13686_, _13643_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_13687_, _13686_, _13658_);
  or (_13688_, _13655_, _13463_);
  and (_13689_, _13688_, _13687_);
  and (_13690_, _13650_, _13469_);
  or (_40785_, _13690_, _13689_);
  or (_13691_, _13655_, _06980_);
  or (_13693_, _13643_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_13694_, _13693_, _13658_);
  and (_13695_, _13694_, _13691_);
  and (_13696_, _13650_, _07006_);
  or (_40786_, _13696_, _13695_);
  and (_13697_, _12449_, _05242_);
  nand (_13698_, _13697_, _13476_);
  or (_13699_, _13698_, _13484_);
  and (_13700_, _13657_, _05123_);
  not (_13701_, _13700_);
  nand (_13703_, _13698_, _04668_);
  and (_13704_, _13703_, _13701_);
  and (_13705_, _13704_, _13699_);
  and (_13706_, _13700_, _12236_);
  or (_40790_, _13706_, _13705_);
  and (_13707_, _13700_, _12443_);
  and (_13708_, _12039_, _04989_);
  and (_13709_, _13642_, _13708_);
  or (_13710_, _13709_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_13711_, _13710_, _13701_);
  not (_13712_, _13709_);
  or (_13713_, _13712_, _12437_);
  and (_13714_, _13713_, _13711_);
  or (_40791_, _13714_, _13707_);
  or (_13715_, _13698_, _12645_);
  or (_13716_, _13709_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_13717_, _13716_, _13701_);
  and (_13718_, _13717_, _13715_);
  and (_13719_, _13700_, _12651_);
  or (_40792_, _13719_, _13718_);
  or (_13720_, _13698_, _13506_);
  or (_13721_, _13709_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_13722_, _13721_, _13701_);
  and (_13723_, _13722_, _13720_);
  and (_13724_, _13700_, _12857_);
  or (_40793_, _13724_, _13723_);
  and (_13725_, _13700_, _13065_);
  or (_13726_, _13698_, _13513_);
  or (_13727_, _13709_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_13728_, _13727_, _13701_);
  and (_13729_, _13728_, _13726_);
  or (_40794_, _13729_, _13725_);
  or (_13730_, _13698_, _13518_);
  nand (_13731_, _13698_, _06861_);
  and (_13732_, _13731_, _13701_);
  and (_13733_, _13732_, _13730_);
  and (_13734_, _13700_, _13264_);
  or (_40796_, _13734_, _13733_);
  or (_13735_, _13709_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_13736_, _13735_, _13701_);
  or (_13737_, _13712_, _13463_);
  and (_13738_, _13737_, _13736_);
  and (_13739_, _13700_, _13469_);
  or (_40797_, _13739_, _13738_);
  or (_13740_, _13698_, _06980_);
  or (_13741_, _13709_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_13742_, _13741_, _13701_);
  and (_13743_, _13742_, _13740_);
  and (_13744_, _13700_, _07006_);
  or (_40798_, _13744_, _13743_);
  and (_13745_, _13697_, _13557_);
  not (_13746_, _13745_);
  or (_13747_, _13746_, _13484_);
  and (_13748_, _13657_, _06162_);
  not (_13749_, _13748_);
  or (_13750_, _13745_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_13751_, _13750_, _13749_);
  and (_13752_, _13751_, _13747_);
  and (_13753_, _13748_, _12236_);
  or (_40802_, _13753_, _13752_);
  and (_13754_, _13642_, _13537_);
  not (_13755_, _13754_);
  or (_13756_, _13755_, _12437_);
  or (_13757_, _13754_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_13758_, _13757_, _13749_);
  and (_13759_, _13758_, _13756_);
  and (_13760_, _13748_, _12443_);
  or (_40803_, _13760_, _13759_);
  or (_13761_, _13754_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_13762_, _13761_, _13749_);
  or (_13763_, _13746_, _12645_);
  and (_13764_, _13763_, _13762_);
  and (_13765_, _13748_, _12651_);
  or (_40804_, _13765_, _13764_);
  or (_13766_, _13754_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_13767_, _13766_, _13749_);
  or (_13768_, _13755_, _12851_);
  and (_13769_, _13768_, _13767_);
  and (_13770_, _13748_, _12857_);
  or (_40805_, _13770_, _13769_);
  or (_13771_, _13754_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_13772_, _13771_, _13749_);
  or (_13773_, _13755_, _13059_);
  and (_13774_, _13773_, _13772_);
  and (_13775_, _13748_, _13065_);
  or (_40806_, _13775_, _13774_);
  or (_13776_, _13754_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_13777_, _13776_, _13749_);
  or (_13778_, _13755_, _13258_);
  and (_13779_, _13778_, _13777_);
  and (_13780_, _13748_, _13264_);
  or (_40808_, _13780_, _13779_);
  or (_13781_, _13754_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_13782_, _13781_, _13749_);
  or (_13783_, _13755_, _13463_);
  and (_13784_, _13783_, _13782_);
  and (_13785_, _13748_, _13469_);
  or (_40809_, _13785_, _13784_);
  or (_13786_, _13754_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_13787_, _13786_, _13749_);
  or (_13788_, _13746_, _06980_);
  and (_13789_, _13788_, _13787_);
  and (_13790_, _13748_, _07006_);
  or (_40810_, _13790_, _13789_);
  and (_13791_, _13697_, _05409_);
  not (_13792_, _13791_);
  or (_13793_, _13792_, _13484_);
  and (_13794_, _13649_, _04837_);
  nor (_13795_, _13791_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_13796_, _13795_, _13794_);
  and (_13797_, _13796_, _13793_);
  and (_13798_, _13794_, _12236_);
  or (_40814_, _13798_, _13797_);
  nand (_13799_, _13657_, _04837_);
  or (_13800_, _13791_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_13801_, _13800_, _13799_);
  or (_13802_, _13792_, _13494_);
  and (_13803_, _13802_, _13801_);
  and (_13804_, _13794_, _12443_);
  or (_40815_, _13804_, _13803_);
  or (_13805_, _13791_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_13806_, _13805_, _13799_);
  or (_13807_, _13792_, _12645_);
  and (_13808_, _13807_, _13806_);
  and (_13809_, _13794_, _12651_);
  or (_40816_, _13809_, _13808_);
  or (_13810_, _13791_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_13811_, _13810_, _13799_);
  or (_13812_, _13792_, _13506_);
  and (_13813_, _13812_, _13811_);
  and (_13814_, _13794_, _12857_);
  or (_40817_, _13814_, _13813_);
  or (_13815_, _13791_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_13816_, _13815_, _13799_);
  or (_13817_, _13792_, _13513_);
  and (_13818_, _13817_, _13816_);
  and (_13819_, _13794_, _13065_);
  or (_40819_, _13819_, _13818_);
  or (_13820_, _13791_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_13821_, _13820_, _13799_);
  or (_13822_, _13792_, _13518_);
  and (_13823_, _13822_, _13821_);
  and (_13824_, _13794_, _13264_);
  or (_40820_, _13824_, _13823_);
  or (_13825_, _13791_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_13826_, _13825_, _13799_);
  or (_13827_, _13792_, _13527_);
  and (_13828_, _13827_, _13826_);
  and (_13829_, _13794_, _13469_);
  or (_40821_, _13829_, _13828_);
  or (_13830_, _13791_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_13831_, _13830_, _13799_);
  or (_13832_, _13792_, _06980_);
  and (_13833_, _13832_, _13831_);
  and (_13834_, _13794_, _07006_);
  or (_40822_, _13834_, _13833_);
  and (_13835_, _12041_, _05385_);
  and (_13836_, _13835_, _12040_);
  nor (_13837_, _13836_, _04681_);
  nand (_13838_, _12050_, _05391_);
  nand (_13839_, _13836_, _12226_);
  nand (_13840_, _13839_, _13838_);
  or (_13841_, _13840_, _13837_);
  not (_13842_, _05393_);
  and (_13843_, _05401_, _13842_);
  and (_13844_, _13843_, _04838_);
  not (_13845_, _13844_);
  or (_13846_, _13845_, _12236_);
  and (_40826_, _13846_, _13841_);
  and (_13847_, _05412_, _05385_);
  and (_13848_, _13847_, _12448_);
  or (_13849_, _13848_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_13850_, _13849_, _13845_);
  not (_13851_, _13848_);
  or (_13852_, _13851_, _13494_);
  and (_13853_, _13852_, _13850_);
  and (_13854_, _13844_, _12443_);
  or (_40828_, _13854_, _13853_);
  or (_13855_, _13848_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_13856_, _13855_, _13845_);
  or (_13857_, _13851_, _12645_);
  and (_13858_, _13857_, _13856_);
  and (_13859_, _13844_, _12651_);
  or (_40829_, _13859_, _13858_);
  or (_13860_, _13848_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_13861_, _13860_, _13845_);
  or (_13862_, _13851_, _13506_);
  and (_13863_, _13862_, _13861_);
  and (_13864_, _13844_, _12857_);
  or (_40830_, _13864_, _13863_);
  or (_13865_, _13848_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_13866_, _13865_, _13845_);
  or (_13867_, _13851_, _13513_);
  and (_13868_, _13867_, _13866_);
  and (_13869_, _13844_, _13065_);
  or (_40831_, _13869_, _13868_);
  or (_13870_, _13851_, _13518_);
  or (_13871_, _13848_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_13872_, _13871_, _13845_);
  and (_13873_, _13872_, _13870_);
  and (_13874_, _13844_, _13264_);
  or (_40832_, _13874_, _13873_);
  or (_13875_, _13848_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_13876_, _13875_, _13845_);
  or (_13877_, _13851_, _13527_);
  and (_13878_, _13877_, _13876_);
  and (_13879_, _13844_, _13469_);
  or (_40834_, _13879_, _13878_);
  or (_13880_, _13848_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_13881_, _13880_, _13845_);
  or (_13882_, _13851_, _06980_);
  and (_13883_, _13882_, _13881_);
  and (_13884_, _13844_, _07006_);
  or (_40835_, _13884_, _13883_);
  and (_13885_, _13847_, _13476_);
  not (_13886_, _13885_);
  or (_13887_, _13886_, _13484_);
  and (_13888_, _13843_, _05123_);
  nor (_13889_, _13885_, \oc8051_golden_model_1.IRAM[9] [0]);
  nor (_13890_, _13889_, _13888_);
  and (_13891_, _13890_, _13887_);
  and (_13892_, _13888_, _12236_);
  or (_40839_, _13892_, _13891_);
  nand (_13893_, _12050_, _05124_);
  or (_13894_, _13885_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_13895_, _13894_, _13893_);
  or (_13896_, _13886_, _13494_);
  and (_13897_, _13896_, _13895_);
  and (_13898_, _13888_, _12443_);
  or (_40840_, _13898_, _13897_);
  or (_13899_, _13885_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_13900_, _13899_, _13893_);
  or (_13901_, _13886_, _12645_);
  and (_13902_, _13901_, _13900_);
  and (_13903_, _13888_, _12651_);
  or (_40841_, _13903_, _13902_);
  or (_13904_, _13885_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_13905_, _13904_, _13893_);
  or (_13906_, _13886_, _13506_);
  and (_13907_, _13906_, _13905_);
  and (_13908_, _13888_, _12857_);
  or (_40842_, _13908_, _13907_);
  or (_13909_, _13885_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_13910_, _13909_, _13893_);
  or (_13911_, _13886_, _13513_);
  and (_13912_, _13911_, _13910_);
  and (_13913_, _13888_, _13065_);
  or (_40843_, _13913_, _13912_);
  or (_13914_, _13886_, _13518_);
  nor (_13915_, _13885_, \oc8051_golden_model_1.IRAM[9] [5]);
  nor (_13916_, _13915_, _13888_);
  and (_13917_, _13916_, _13914_);
  and (_13918_, _13888_, _13264_);
  or (_40845_, _13918_, _13917_);
  or (_13919_, _13885_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_13920_, _13919_, _13893_);
  or (_13921_, _13886_, _13527_);
  and (_13922_, _13921_, _13920_);
  and (_13923_, _13888_, _13469_);
  or (_40846_, _13923_, _13922_);
  or (_13924_, _13885_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_13925_, _13924_, _13893_);
  or (_13926_, _13886_, _06980_);
  and (_13927_, _13926_, _13925_);
  and (_13928_, _13888_, _07006_);
  or (_40847_, _13928_, _13927_);
  and (_13929_, _13847_, _13557_);
  not (_13930_, _13929_);
  or (_13931_, _13930_, _13484_);
  and (_13932_, _13843_, _06162_);
  not (_13933_, _13932_);
  or (_13934_, _13929_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_13935_, _13934_, _13933_);
  and (_13936_, _13935_, _13931_);
  and (_13937_, _13932_, _12236_);
  or (_40851_, _13937_, _13936_);
  or (_13938_, _13929_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_13939_, _13938_, _13933_);
  or (_13940_, _13930_, _13494_);
  and (_13941_, _13940_, _13939_);
  and (_13942_, _13932_, _12443_);
  or (_40852_, _13942_, _13941_);
  or (_13943_, _13929_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_13944_, _13943_, _13933_);
  or (_13945_, _13930_, _12645_);
  and (_13946_, _13945_, _13944_);
  and (_13947_, _13932_, _12651_);
  or (_40853_, _13947_, _13946_);
  or (_13948_, _13929_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_13949_, _13948_, _13933_);
  or (_13950_, _13930_, _13506_);
  and (_13951_, _13950_, _13949_);
  and (_13952_, _13932_, _12857_);
  or (_40854_, _13952_, _13951_);
  or (_13953_, _13930_, _13513_);
  or (_13954_, _13929_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_13955_, _13954_, _13933_);
  and (_13956_, _13955_, _13953_);
  and (_13957_, _13932_, _13065_);
  or (_40855_, _13957_, _13956_);
  or (_13958_, _13929_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_13959_, _13958_, _13933_);
  or (_13960_, _13930_, _13518_);
  and (_13961_, _13960_, _13959_);
  and (_13962_, _13932_, _13264_);
  or (_40857_, _13962_, _13961_);
  or (_13963_, _13929_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_13964_, _13963_, _13933_);
  or (_13965_, _13930_, _13527_);
  and (_13966_, _13965_, _13964_);
  and (_13967_, _13932_, _13469_);
  or (_40858_, _13967_, _13966_);
  or (_13968_, _13929_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_13969_, _13968_, _13933_);
  or (_13970_, _13930_, _06980_);
  and (_13971_, _13970_, _13969_);
  and (_13972_, _13932_, _07006_);
  or (_40859_, _13972_, _13971_);
  and (_13973_, _13847_, _05409_);
  not (_13974_, _13973_);
  or (_13975_, _13974_, _13484_);
  and (_13976_, _13843_, _04837_);
  not (_13977_, _13976_);
  or (_13978_, _13973_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_13979_, _13978_, _13977_);
  and (_13980_, _13979_, _13975_);
  and (_13981_, _13976_, _12236_);
  or (_40863_, _13981_, _13980_);
  or (_13982_, _13973_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_13983_, _13982_, _13977_);
  or (_13984_, _13974_, _13494_);
  and (_13985_, _13984_, _13983_);
  and (_13986_, _13976_, _12443_);
  or (_40864_, _13986_, _13985_);
  or (_13987_, _13973_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_13988_, _13987_, _13977_);
  or (_13989_, _13974_, _12645_);
  and (_13990_, _13989_, _13988_);
  and (_13991_, _13976_, _12651_);
  or (_40865_, _13991_, _13990_);
  or (_13992_, _13973_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_13993_, _13992_, _13977_);
  or (_13994_, _13974_, _13506_);
  and (_13995_, _13994_, _13993_);
  and (_13996_, _13976_, _12857_);
  or (_40866_, _13996_, _13995_);
  or (_13997_, _13973_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_13998_, _13997_, _13977_);
  or (_13999_, _13974_, _13513_);
  and (_14000_, _13999_, _13998_);
  and (_14001_, _13976_, _13065_);
  or (_40868_, _14001_, _14000_);
  or (_14002_, _13973_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_14003_, _14002_, _13977_);
  or (_14004_, _13974_, _13518_);
  and (_14005_, _14004_, _14003_);
  and (_14006_, _13976_, _13264_);
  or (_40869_, _14006_, _14005_);
  or (_14007_, _13973_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_14008_, _14007_, _13977_);
  or (_14009_, _13974_, _13527_);
  and (_14010_, _14009_, _14008_);
  and (_14011_, _13976_, _13469_);
  or (_40870_, _14011_, _14010_);
  or (_14012_, _13973_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_14013_, _14012_, _13977_);
  or (_14014_, _13974_, _06980_);
  and (_14015_, _14014_, _14013_);
  and (_14016_, _13976_, _07006_);
  or (_40871_, _14016_, _14015_);
  and (_14017_, _12448_, _05413_);
  not (_14018_, _14017_);
  or (_14019_, _14018_, _13484_);
  and (_14020_, _05402_, _04838_);
  not (_14021_, _14020_);
  or (_14022_, _14017_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_14023_, _14022_, _14021_);
  and (_14024_, _14023_, _14019_);
  and (_14025_, _14020_, _12236_);
  or (_40875_, _14025_, _14024_);
  and (_14026_, _12040_, _05388_);
  or (_14027_, _14026_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_14028_, _14027_, _14021_);
  or (_14029_, _14018_, _13494_);
  and (_14030_, _14029_, _14028_);
  and (_14031_, _14020_, _12443_);
  or (_40876_, _14031_, _14030_);
  or (_14032_, _14026_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_14033_, _14032_, _14021_);
  or (_14034_, _14018_, _12645_);
  and (_14035_, _14034_, _14033_);
  and (_14036_, _14020_, _12651_);
  or (_40877_, _14036_, _14035_);
  or (_14037_, _14026_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_14038_, _14037_, _14021_);
  or (_14039_, _14018_, _13506_);
  and (_14040_, _14039_, _14038_);
  and (_14041_, _14020_, _12857_);
  or (_40879_, _14041_, _14040_);
  or (_14042_, _14018_, _13513_);
  or (_14043_, _14026_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_14044_, _14043_, _14021_);
  and (_14045_, _14044_, _14042_);
  and (_14046_, _14020_, _13065_);
  or (_40880_, _14046_, _14045_);
  or (_14047_, _14018_, _13518_);
  or (_14048_, _14017_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_14049_, _14048_, _14021_);
  and (_14050_, _14049_, _14047_);
  and (_14051_, _14020_, _13264_);
  or (_40881_, _14051_, _14050_);
  or (_14052_, _14026_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_14053_, _14052_, _14021_);
  or (_14054_, _14018_, _13527_);
  and (_14055_, _14054_, _14053_);
  and (_14056_, _14020_, _13469_);
  or (_40882_, _14056_, _14055_);
  or (_14057_, _14026_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_14058_, _14057_, _14021_);
  or (_14059_, _14018_, _06980_);
  and (_14060_, _14059_, _14058_);
  and (_14061_, _14020_, _07006_);
  or (_40883_, _14061_, _14060_);
  and (_14062_, _13476_, _05413_);
  not (_14063_, _14062_);
  or (_14064_, _14063_, _13484_);
  and (_14065_, _05402_, _05123_);
  not (_14066_, _14065_);
  or (_14067_, _14062_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_14068_, _14067_, _14066_);
  and (_14069_, _14068_, _14064_);
  and (_14070_, _14065_, _12236_);
  or (_40887_, _14070_, _14069_);
  and (_14071_, _13708_, _05388_);
  or (_14072_, _14071_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_14073_, _14072_, _14066_);
  not (_14074_, _14071_);
  or (_14075_, _14074_, _12437_);
  and (_14076_, _14075_, _14073_);
  and (_14077_, _14065_, _12443_);
  or (_40888_, _14077_, _14076_);
  or (_14078_, _14071_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_14079_, _14078_, _14066_);
  or (_14080_, _14063_, _12645_);
  and (_14081_, _14080_, _14079_);
  and (_14082_, _14065_, _12651_);
  or (_40890_, _14082_, _14081_);
  or (_14083_, _14071_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_14084_, _14083_, _14066_);
  or (_14085_, _14074_, _12851_);
  and (_14086_, _14085_, _14084_);
  and (_14087_, _14065_, _12857_);
  or (_40891_, _14087_, _14086_);
  or (_14088_, _14071_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_14089_, _14088_, _14066_);
  or (_14090_, _14074_, _13059_);
  and (_14091_, _14090_, _14089_);
  and (_14092_, _14065_, _13065_);
  or (_40892_, _14092_, _14091_);
  or (_14093_, _14063_, _13518_);
  or (_14094_, _14062_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_14095_, _14094_, _14066_);
  and (_14096_, _14095_, _14093_);
  and (_14097_, _14065_, _13264_);
  or (_40893_, _14097_, _14096_);
  or (_14098_, _14071_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_14099_, _14098_, _14066_);
  or (_14100_, _14074_, _13463_);
  and (_14101_, _14100_, _14099_);
  and (_14102_, _14065_, _13469_);
  or (_40894_, _14102_, _14101_);
  or (_14103_, _14071_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_14104_, _14103_, _14066_);
  or (_14105_, _14063_, _06980_);
  and (_14106_, _14105_, _14104_);
  and (_14107_, _14065_, _07006_);
  or (_40896_, _14107_, _14106_);
  and (_14108_, _13557_, _05413_);
  not (_14109_, _14108_);
  or (_14110_, _14109_, _13484_);
  and (_14111_, _06162_, _05402_);
  not (_14112_, _14111_);
  or (_14113_, _14108_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_14114_, _14113_, _14112_);
  and (_14115_, _14114_, _14110_);
  and (_14116_, _14111_, _12236_);
  or (_40899_, _14116_, _14115_);
  and (_14117_, _13537_, _05388_);
  or (_14118_, _14117_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_14119_, _14118_, _14112_);
  not (_14120_, _14117_);
  or (_14121_, _14120_, _12437_);
  and (_14122_, _14121_, _14119_);
  and (_14123_, _14111_, _12443_);
  or (_40900_, _14123_, _14122_);
  or (_14124_, _14117_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_14125_, _14124_, _14112_);
  or (_14126_, _14109_, _12645_);
  and (_14127_, _14126_, _14125_);
  and (_14128_, _14111_, _12651_);
  or (_40902_, _14128_, _14127_);
  or (_14129_, _14117_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_14130_, _14129_, _14112_);
  or (_14131_, _14120_, _12851_);
  and (_14132_, _14131_, _14130_);
  and (_14133_, _14111_, _12857_);
  or (_40903_, _14133_, _14132_);
  or (_14134_, _14117_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_14135_, _14134_, _14112_);
  or (_14136_, _14120_, _13059_);
  and (_14137_, _14136_, _14135_);
  and (_14138_, _14111_, _13065_);
  or (_40904_, _14138_, _14137_);
  or (_14139_, _14117_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_14140_, _14139_, _14112_);
  or (_14141_, _14120_, _13258_);
  and (_14142_, _14141_, _14140_);
  and (_14143_, _14111_, _13264_);
  or (_40905_, _14143_, _14142_);
  or (_14144_, _14117_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_14145_, _14144_, _14112_);
  or (_14146_, _14120_, _13463_);
  and (_14147_, _14146_, _14145_);
  and (_14148_, _14111_, _13469_);
  or (_40906_, _14148_, _14147_);
  or (_14149_, _14117_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_14150_, _14149_, _14112_);
  or (_14151_, _14109_, _06980_);
  and (_14152_, _14151_, _14150_);
  and (_14153_, _14111_, _07006_);
  or (_40908_, _14153_, _14152_);
  or (_14154_, _13484_, _05415_);
  or (_14155_, _05414_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_14156_, _14155_, _05404_);
  and (_14157_, _14156_, _14154_);
  and (_14158_, _12236_, _05403_);
  or (_40911_, _14158_, _14157_);
  or (_14159_, _05389_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_14160_, _14159_, _05404_);
  not (_14161_, _05389_);
  or (_14162_, _12437_, _14161_);
  and (_14163_, _14162_, _14160_);
  and (_14164_, _12443_, _05403_);
  or (_40912_, _14164_, _14163_);
  or (_14165_, _05389_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_14166_, _14165_, _05404_);
  or (_14167_, _12645_, _05415_);
  and (_14168_, _14167_, _14166_);
  and (_14169_, _12651_, _05403_);
  or (_40914_, _14169_, _14168_);
  or (_14170_, _05389_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_14171_, _14170_, _05404_);
  or (_14172_, _12851_, _14161_);
  and (_14173_, _14172_, _14171_);
  and (_14174_, _12857_, _05403_);
  or (_40915_, _14174_, _14173_);
  or (_14175_, _05389_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_14176_, _14175_, _05404_);
  or (_14177_, _13059_, _14161_);
  and (_14178_, _14177_, _14176_);
  and (_14179_, _13065_, _05403_);
  or (_40916_, _14179_, _14178_);
  or (_14180_, _05389_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_14181_, _14180_, _05404_);
  or (_14182_, _13258_, _14161_);
  and (_14183_, _14182_, _14181_);
  and (_14184_, _13264_, _05403_);
  or (_40917_, _14184_, _14183_);
  or (_14185_, _05389_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_14186_, _14185_, _05404_);
  or (_14187_, _13463_, _14161_);
  and (_14188_, _14187_, _14186_);
  and (_14189_, _13469_, _05403_);
  or (_40918_, _14189_, _14188_);
  nor (_14190_, _43152_, _07054_);
  nand (_14191_, _08753_, _05440_);
  nor (_14192_, _05440_, _07054_);
  nor (_14193_, _14192_, _04785_);
  nand (_14194_, _14193_, _14191_);
  and (_14195_, _05440_, _06479_);
  or (_14196_, _14195_, _14192_);
  or (_14197_, _14196_, _04778_);
  nor (_14198_, _12164_, _07937_);
  or (_14199_, _14198_, _14192_);
  and (_14200_, _14199_, _03455_);
  and (_14201_, _05440_, _04700_);
  or (_14202_, _14201_, _14192_);
  or (_14203_, _14202_, _04733_);
  and (_14204_, _05716_, _05440_);
  or (_14205_, _14204_, _14192_);
  or (_14206_, _14205_, _04722_);
  and (_14207_, _05440_, \oc8051_golden_model_1.ACC [0]);
  or (_14208_, _14207_, _14192_);
  and (_14209_, _14208_, _04707_);
  nor (_14210_, _04707_, _07054_);
  or (_14211_, _14210_, _03850_);
  or (_14212_, _14211_, _14209_);
  and (_14213_, _14212_, _03764_);
  and (_14214_, _14213_, _14206_);
  nor (_14215_, _06088_, _07054_);
  and (_14216_, _12064_, _06088_);
  or (_14217_, _14216_, _14215_);
  and (_14218_, _14217_, _03763_);
  or (_14219_, _14218_, _14214_);
  or (_14220_, _14219_, _03848_);
  and (_14221_, _14220_, _14203_);
  or (_14222_, _14221_, _03854_);
  or (_14223_, _14208_, _03855_);
  and (_14224_, _14223_, _03760_);
  and (_14225_, _14224_, _14222_);
  and (_14226_, _14192_, _03759_);
  or (_14227_, _14226_, _03752_);
  or (_14228_, _14227_, _14225_);
  or (_14229_, _14205_, _03753_);
  and (_14230_, _14229_, _14228_);
  or (_14231_, _14230_, _07399_);
  nor (_14232_, _07876_, _07874_);
  nor (_14233_, _14232_, _07877_);
  or (_14234_, _14233_, _07405_);
  and (_14235_, _14234_, _03747_);
  and (_14236_, _14235_, _14231_);
  nand (_14237_, _05432_, _08297_);
  or (_14238_, _14215_, _14237_);
  and (_14239_, _14238_, _03746_);
  and (_14240_, _14239_, _14217_);
  or (_14241_, _14240_, _07927_);
  or (_14242_, _14241_, _14236_);
  and (_14243_, _06962_, _05440_);
  or (_14244_, _14192_, _03738_);
  or (_14245_, _14244_, _14243_);
  or (_14246_, _14202_, _07925_);
  and (_14247_, _14246_, _03820_);
  and (_14248_, _14247_, _14245_);
  and (_14249_, _14248_, _14242_);
  or (_14250_, _14249_, _14200_);
  and (_14251_, _14250_, _07011_);
  nand (_14252_, _07364_, _03498_);
  nor (_14253_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_14254_, _14253_, _07855_);
  or (_14255_, _07364_, _14254_);
  and (_14256_, _14255_, _07010_);
  and (_14257_, _14256_, _14252_);
  or (_14258_, _14257_, _03903_);
  or (_14259_, _14258_, _14251_);
  and (_14260_, _14259_, _14197_);
  or (_14261_, _14260_, _03897_);
  and (_14262_, _12178_, _05440_);
  or (_14263_, _14192_, _04790_);
  or (_14264_, _14263_, _14262_);
  and (_14265_, _14264_, _04792_);
  and (_14266_, _14265_, _14261_);
  nor (_14267_, _10488_, _07937_);
  or (_14268_, _14267_, _14192_);
  and (_14269_, _14191_, _04018_);
  and (_14270_, _14269_, _14268_);
  or (_14271_, _14270_, _14266_);
  and (_14272_, _14271_, _03909_);
  nand (_14273_, _14196_, _03908_);
  nor (_14274_, _14273_, _14204_);
  or (_14275_, _14274_, _04027_);
  or (_14276_, _14275_, _14272_);
  and (_14277_, _14276_, _14194_);
  or (_14278_, _14277_, _03914_);
  nor (_14279_, _12177_, _07937_);
  or (_14280_, _14192_, _06567_);
  or (_14281_, _14280_, _14279_);
  and (_14282_, _14281_, _06572_);
  and (_14283_, _14282_, _14278_);
  and (_14284_, _14268_, _04011_);
  or (_14285_, _14284_, _03773_);
  or (_14286_, _14285_, _14283_);
  or (_14287_, _14205_, _03774_);
  and (_14288_, _14287_, _14286_);
  or (_14289_, _14288_, _03374_);
  or (_14290_, _14192_, _03375_);
  and (_14291_, _14290_, _14289_);
  or (_14292_, _14291_, _03772_);
  or (_14293_, _14205_, _04060_);
  and (_14294_, _14293_, _43152_);
  and (_14295_, _14294_, _14292_);
  or (_14296_, _14295_, _14190_);
  and (_43376_, _14296_, _41894_);
  nor (_14297_, _43152_, _07015_);
  nor (_14298_, _05440_, _07015_);
  nor (_14299_, _08751_, _07937_);
  or (_14300_, _14299_, _14298_);
  or (_14301_, _14300_, _06572_);
  nand (_14302_, _05440_, _04595_);
  or (_14303_, _05440_, \oc8051_golden_model_1.B [1]);
  and (_14304_, _14303_, _03903_);
  and (_14305_, _14304_, _14302_);
  nor (_14306_, _06088_, _07015_);
  and (_14307_, _12252_, _06088_);
  or (_14308_, _14307_, _14306_);
  and (_14309_, _14308_, _03759_);
  and (_14310_, _05440_, _04900_);
  or (_14311_, _14310_, _14298_);
  or (_14312_, _14311_, _04733_);
  and (_14313_, _12262_, _05440_);
  not (_14314_, _14313_);
  and (_14315_, _14314_, _14303_);
  or (_14316_, _14315_, _04722_);
  and (_14317_, _05440_, \oc8051_golden_model_1.ACC [1]);
  or (_14318_, _14317_, _14298_);
  and (_14319_, _14318_, _04707_);
  nor (_14320_, _04707_, _07015_);
  or (_14321_, _14320_, _03850_);
  or (_14322_, _14321_, _14319_);
  and (_14323_, _14322_, _03764_);
  and (_14324_, _14323_, _14316_);
  and (_14325_, _12249_, _06088_);
  or (_14326_, _14325_, _14306_);
  and (_14327_, _14326_, _03763_);
  or (_14328_, _14327_, _03848_);
  or (_14329_, _14328_, _14324_);
  and (_14330_, _14329_, _14312_);
  or (_14331_, _14330_, _03854_);
  or (_14332_, _14318_, _03855_);
  and (_14333_, _14332_, _03760_);
  and (_14334_, _14333_, _14331_);
  or (_14335_, _14334_, _14309_);
  and (_14336_, _14335_, _03753_);
  and (_14337_, _14325_, _12248_);
  or (_14338_, _14337_, _14306_);
  and (_14339_, _14338_, _03752_);
  or (_14340_, _14339_, _07399_);
  or (_14341_, _14340_, _14336_);
  nor (_14342_, _07879_, _07823_);
  nor (_14343_, _14342_, _07880_);
  or (_14344_, _14343_, _07405_);
  and (_14345_, _14344_, _03747_);
  and (_14346_, _14345_, _14341_);
  nor (_14347_, _12293_, _07915_);
  or (_14348_, _14347_, _14306_);
  and (_14349_, _14348_, _03746_);
  or (_14350_, _14349_, _07927_);
  or (_14351_, _14350_, _14346_);
  and (_14352_, _06961_, _05440_);
  or (_14353_, _14298_, _03738_);
  or (_14354_, _14353_, _14352_);
  or (_14355_, _14311_, _07925_);
  and (_14356_, _14355_, _03820_);
  and (_14357_, _14356_, _14354_);
  and (_14358_, _14357_, _14351_);
  nand (_14359_, _12352_, _05440_);
  and (_14360_, _14303_, _03455_);
  and (_14361_, _14360_, _14359_);
  or (_14362_, _14361_, _07010_);
  or (_14363_, _14362_, _14358_);
  and (_14364_, _07364_, _07310_);
  nor (_14365_, _07359_, _07358_);
  or (_14366_, _14365_, _07360_);
  nor (_14367_, _14366_, _07364_);
  or (_14368_, _14367_, _14364_);
  or (_14369_, _14368_, _07011_);
  and (_14370_, _14369_, _04778_);
  and (_14371_, _14370_, _14363_);
  or (_14372_, _14371_, _14305_);
  and (_14373_, _14372_, _04790_);
  or (_14374_, _12366_, _07937_);
  and (_14375_, _14303_, _03897_);
  and (_14376_, _14375_, _14374_);
  or (_14377_, _14376_, _04018_);
  or (_14378_, _14377_, _14373_);
  nand (_14379_, _08750_, _05440_);
  and (_14380_, _14379_, _14300_);
  or (_14381_, _14380_, _04792_);
  and (_14382_, _14381_, _03909_);
  and (_14383_, _14382_, _14378_);
  or (_14384_, _12244_, _07937_);
  and (_14385_, _14303_, _03908_);
  and (_14386_, _14385_, _14384_);
  or (_14387_, _14386_, _04027_);
  or (_14388_, _14387_, _14383_);
  nor (_14389_, _14298_, _04785_);
  nand (_14390_, _14389_, _14379_);
  and (_14391_, _14390_, _06567_);
  and (_14392_, _14391_, _14388_);
  or (_14393_, _14302_, _08366_);
  and (_14394_, _14303_, _03914_);
  and (_14395_, _14394_, _14393_);
  or (_14396_, _14395_, _04011_);
  or (_14397_, _14396_, _14392_);
  and (_14398_, _14397_, _14301_);
  or (_14399_, _14398_, _03773_);
  or (_14400_, _14315_, _03774_);
  and (_14401_, _14400_, _03375_);
  and (_14402_, _14401_, _14399_);
  and (_14403_, _14308_, _03374_);
  or (_14404_, _14403_, _03772_);
  or (_14405_, _14404_, _14402_);
  or (_14406_, _14298_, _04060_);
  or (_14407_, _14406_, _14313_);
  and (_14408_, _14407_, _43152_);
  and (_14409_, _14408_, _14405_);
  or (_14410_, _14409_, _14297_);
  and (_43377_, _14410_, _41894_);
  nor (_14411_, _43152_, _07027_);
  nor (_14412_, _05440_, _07027_);
  and (_14413_, _05440_, _06495_);
  or (_14414_, _14413_, _14412_);
  or (_14415_, _14414_, _04778_);
  nor (_14416_, _12572_, _07937_);
  or (_14417_, _14416_, _14412_);
  and (_14418_, _14417_, _03455_);
  nor (_14419_, _06088_, _07027_);
  and (_14420_, _12467_, _06088_);
  or (_14421_, _14420_, _14419_);
  and (_14422_, _14421_, _03759_);
  and (_14423_, _05440_, _05307_);
  or (_14424_, _14423_, _14412_);
  or (_14425_, _14424_, _04733_);
  nor (_14426_, _12471_, _07937_);
  or (_14427_, _14426_, _14412_);
  or (_14428_, _14427_, _04722_);
  and (_14429_, _05440_, \oc8051_golden_model_1.ACC [2]);
  or (_14430_, _14429_, _14412_);
  and (_14431_, _14430_, _04707_);
  nor (_14432_, _04707_, _07027_);
  or (_14433_, _14432_, _03850_);
  or (_14434_, _14433_, _14431_);
  and (_14435_, _14434_, _03764_);
  and (_14436_, _14435_, _14428_);
  and (_14437_, _12464_, _06088_);
  or (_14438_, _14437_, _14419_);
  and (_14439_, _14438_, _03763_);
  or (_14440_, _14439_, _03848_);
  or (_14441_, _14440_, _14436_);
  and (_14442_, _14441_, _14425_);
  or (_14443_, _14442_, _03854_);
  or (_14444_, _14430_, _03855_);
  and (_14445_, _14444_, _03760_);
  and (_14446_, _14445_, _14443_);
  or (_14447_, _14446_, _14422_);
  and (_14448_, _14447_, _03753_);
  and (_14449_, _14437_, _12463_);
  or (_14450_, _14449_, _14419_);
  and (_14451_, _14450_, _03752_);
  or (_14452_, _14451_, _07399_);
  or (_14453_, _14452_, _14448_);
  or (_14454_, _07881_, _07779_);
  and (_14455_, _14454_, _07882_);
  or (_14456_, _14455_, _07405_);
  and (_14457_, _14456_, _03747_);
  and (_14458_, _14457_, _14453_);
  nor (_14459_, _12514_, _07915_);
  or (_14460_, _14459_, _14419_);
  and (_14461_, _14460_, _03746_);
  or (_14462_, _14461_, _07927_);
  or (_14463_, _14462_, _14458_);
  and (_14464_, _06965_, _05440_);
  or (_14465_, _14412_, _03738_);
  or (_14466_, _14465_, _14464_);
  or (_14467_, _14424_, _07925_);
  and (_14468_, _14467_, _03820_);
  and (_14469_, _14468_, _14466_);
  and (_14470_, _14469_, _14463_);
  or (_14471_, _14470_, _14418_);
  and (_14472_, _14471_, _07011_);
  nor (_14473_, _07360_, _07311_);
  not (_14474_, _14473_);
  and (_14475_, _14474_, _07303_);
  nor (_14476_, _14474_, _07303_);
  nor (_14477_, _14476_, _14475_);
  or (_14478_, _14477_, _07364_);
  nand (_14479_, _07364_, _07300_);
  and (_14480_, _14479_, _07010_);
  and (_14481_, _14480_, _14478_);
  or (_14482_, _14481_, _03903_);
  or (_14483_, _14482_, _14472_);
  and (_14484_, _14483_, _14415_);
  or (_14485_, _14484_, _03897_);
  and (_14486_, _12586_, _05440_);
  or (_14487_, _14412_, _04790_);
  or (_14488_, _14487_, _14486_);
  and (_14489_, _14488_, _04792_);
  and (_14490_, _14489_, _14485_);
  and (_14491_, _08748_, _05440_);
  or (_14492_, _14491_, _14412_);
  and (_14493_, _14492_, _04018_);
  or (_14494_, _14493_, _14490_);
  and (_14495_, _14494_, _03909_);
  or (_14496_, _14412_, _05765_);
  and (_14497_, _14414_, _03908_);
  and (_14498_, _14497_, _14496_);
  or (_14499_, _14498_, _14495_);
  and (_14500_, _14499_, _04785_);
  and (_14501_, _14430_, _04027_);
  and (_14502_, _14501_, _14496_);
  or (_14503_, _14502_, _03914_);
  or (_14504_, _14503_, _14500_);
  nor (_14505_, _12585_, _07937_);
  or (_14506_, _14412_, _06567_);
  or (_14507_, _14506_, _14505_);
  and (_14508_, _14507_, _06572_);
  and (_14509_, _14508_, _14504_);
  nor (_14510_, _08747_, _07937_);
  or (_14511_, _14510_, _14412_);
  and (_14512_, _14511_, _04011_);
  or (_14513_, _14512_, _03773_);
  or (_14514_, _14513_, _14509_);
  or (_14515_, _14427_, _03774_);
  and (_14516_, _14515_, _03375_);
  and (_14517_, _14516_, _14514_);
  and (_14518_, _14421_, _03374_);
  or (_14519_, _14518_, _03772_);
  or (_14520_, _14519_, _14517_);
  and (_14521_, _12642_, _05440_);
  or (_14522_, _14412_, _04060_);
  or (_14523_, _14522_, _14521_);
  and (_14524_, _14523_, _43152_);
  and (_14525_, _14524_, _14520_);
  or (_14526_, _14525_, _14411_);
  and (_43378_, _14526_, _41894_);
  nor (_14527_, _43152_, _07028_);
  nor (_14528_, _05440_, _07028_);
  and (_14529_, _05440_, _06345_);
  or (_14530_, _14529_, _14528_);
  or (_14531_, _14530_, _04778_);
  nor (_14532_, _12775_, _07937_);
  or (_14533_, _14532_, _14528_);
  and (_14534_, _14533_, _03455_);
  nor (_14535_, _06088_, _07028_);
  and (_14536_, _12674_, _06088_);
  or (_14537_, _14536_, _14535_);
  or (_14538_, _14535_, _12673_);
  and (_14539_, _14538_, _14537_);
  or (_14540_, _14539_, _03753_);
  nor (_14541_, _12681_, _07937_);
  or (_14542_, _14541_, _14528_);
  or (_14543_, _14542_, _04722_);
  and (_14544_, _05440_, \oc8051_golden_model_1.ACC [3]);
  or (_14545_, _14544_, _14528_);
  and (_14546_, _14545_, _04707_);
  nor (_14547_, _04707_, _07028_);
  or (_14548_, _14547_, _03850_);
  or (_14549_, _14548_, _14546_);
  and (_14550_, _14549_, _03764_);
  and (_14551_, _14550_, _14543_);
  and (_14552_, _14537_, _03763_);
  or (_14553_, _14552_, _03848_);
  or (_14554_, _14553_, _14551_);
  and (_14555_, _05440_, _05119_);
  or (_14556_, _14555_, _14528_);
  or (_14557_, _14556_, _04733_);
  and (_14558_, _14557_, _14554_);
  or (_14559_, _14558_, _03854_);
  or (_14560_, _14545_, _03855_);
  and (_14561_, _14560_, _03760_);
  and (_14562_, _14561_, _14559_);
  and (_14563_, _12667_, _06088_);
  or (_14564_, _14563_, _14535_);
  and (_14565_, _14564_, _03759_);
  or (_14566_, _14565_, _03752_);
  or (_14567_, _14566_, _14562_);
  and (_14568_, _14567_, _14540_);
  or (_14569_, _14568_, _07399_);
  nor (_14570_, _07884_, _07722_);
  nor (_14571_, _14570_, _07885_);
  or (_14572_, _14571_, _07405_);
  and (_14573_, _14572_, _03747_);
  and (_14574_, _14573_, _14569_);
  nor (_14575_, _12668_, _07915_);
  or (_14576_, _14575_, _14535_);
  and (_14577_, _14576_, _03746_);
  or (_14578_, _14577_, _07927_);
  or (_14579_, _14578_, _14574_);
  and (_14580_, _06964_, _05440_);
  or (_14581_, _14528_, _03738_);
  or (_14582_, _14581_, _14580_);
  or (_14583_, _14556_, _07925_);
  and (_14584_, _14583_, _03820_);
  and (_14585_, _14584_, _14582_);
  and (_14586_, _14585_, _14579_);
  or (_14587_, _14586_, _14534_);
  and (_14588_, _14587_, _07011_);
  nand (_14589_, _07364_, _07291_);
  nor (_14590_, _14475_, _07302_);
  nor (_14591_, _14590_, _07294_);
  and (_14592_, _14590_, _07294_);
  or (_14593_, _14592_, _14591_);
  or (_14594_, _14593_, _07364_);
  and (_14595_, _14594_, _07010_);
  and (_14596_, _14595_, _14589_);
  or (_14597_, _14596_, _03903_);
  or (_14598_, _14597_, _14588_);
  and (_14599_, _14598_, _14531_);
  or (_14600_, _14599_, _03897_);
  and (_14601_, _12789_, _05440_);
  or (_14602_, _14528_, _04790_);
  or (_14603_, _14602_, _14601_);
  and (_14604_, _14603_, _04792_);
  and (_14605_, _14604_, _14600_);
  and (_14606_, _10491_, _05440_);
  or (_14607_, _14606_, _14528_);
  and (_14608_, _14607_, _04018_);
  or (_14609_, _14608_, _14605_);
  and (_14610_, _14609_, _03909_);
  or (_14611_, _14528_, _05622_);
  and (_14612_, _14530_, _03908_);
  and (_14613_, _14612_, _14611_);
  or (_14614_, _14613_, _14610_);
  and (_14615_, _14614_, _04785_);
  and (_14616_, _14545_, _04027_);
  and (_14617_, _14616_, _14611_);
  or (_14618_, _14617_, _03914_);
  or (_14619_, _14618_, _14615_);
  nor (_14620_, _12788_, _07937_);
  or (_14621_, _14528_, _06567_);
  or (_14622_, _14621_, _14620_);
  and (_14623_, _14622_, _06572_);
  and (_14624_, _14623_, _14619_);
  nor (_14625_, _08742_, _07937_);
  or (_14626_, _14625_, _14528_);
  and (_14627_, _14626_, _04011_);
  or (_14628_, _14627_, _03773_);
  or (_14629_, _14628_, _14624_);
  or (_14630_, _14542_, _03774_);
  and (_14631_, _14630_, _03375_);
  and (_14632_, _14631_, _14629_);
  and (_14633_, _14564_, _03374_);
  or (_14634_, _14633_, _03772_);
  or (_14635_, _14634_, _14632_);
  and (_14636_, _12848_, _05440_);
  or (_14637_, _14528_, _04060_);
  or (_14638_, _14637_, _14636_);
  and (_14639_, _14638_, _43152_);
  and (_14640_, _14639_, _14635_);
  or (_14641_, _14640_, _14527_);
  and (_43379_, _14641_, _41894_);
  nor (_14642_, _43152_, _07029_);
  nor (_14643_, _05440_, _07029_);
  and (_14644_, _06456_, _05440_);
  or (_14645_, _14644_, _14643_);
  or (_14646_, _14645_, _04778_);
  nor (_14647_, _12982_, _07937_);
  or (_14648_, _14647_, _14643_);
  and (_14649_, _14648_, _03455_);
  nor (_14650_, _06088_, _07029_);
  and (_14651_, _12870_, _06088_);
  or (_14652_, _14651_, _14650_);
  and (_14653_, _14652_, _03759_);
  nor (_14654_, _12891_, _07937_);
  or (_14655_, _14654_, _14643_);
  or (_14656_, _14655_, _04722_);
  and (_14657_, _05440_, \oc8051_golden_model_1.ACC [4]);
  or (_14658_, _14657_, _14643_);
  and (_14659_, _14658_, _04707_);
  nor (_14660_, _04707_, _07029_);
  or (_14661_, _14660_, _03850_);
  or (_14662_, _14661_, _14659_);
  and (_14663_, _14662_, _03764_);
  and (_14664_, _14663_, _14656_);
  and (_14665_, _12875_, _06088_);
  or (_14666_, _14665_, _14650_);
  and (_14667_, _14666_, _03763_);
  or (_14668_, _14667_, _03848_);
  or (_14669_, _14668_, _14664_);
  and (_14670_, _05950_, _05440_);
  or (_14671_, _14670_, _14643_);
  or (_14672_, _14671_, _04733_);
  and (_14673_, _14672_, _14669_);
  or (_14674_, _14673_, _03854_);
  or (_14675_, _14658_, _03855_);
  and (_14676_, _14675_, _03760_);
  and (_14677_, _14676_, _14674_);
  or (_14678_, _14677_, _14653_);
  and (_14679_, _14678_, _03753_);
  or (_14680_, _14650_, _12874_);
  and (_14681_, _14680_, _03752_);
  and (_14682_, _14681_, _14666_);
  or (_14683_, _14682_, _07399_);
  or (_14684_, _14683_, _14679_);
  or (_14685_, _07888_, _07886_);
  and (_14686_, _14685_, _07889_);
  or (_14687_, _14686_, _07405_);
  and (_14688_, _14687_, _03747_);
  and (_14689_, _14688_, _14684_);
  nor (_14690_, _12872_, _07915_);
  or (_14691_, _14690_, _14650_);
  and (_14692_, _14691_, _03746_);
  or (_14693_, _14692_, _07927_);
  or (_14694_, _14693_, _14689_);
  and (_14695_, _06969_, _05440_);
  or (_14696_, _14643_, _03738_);
  or (_14697_, _14696_, _14695_);
  or (_14698_, _14671_, _07925_);
  and (_14699_, _14698_, _03820_);
  and (_14700_, _14699_, _14697_);
  and (_14701_, _14700_, _14694_);
  or (_14702_, _14701_, _14649_);
  and (_14703_, _14702_, _07011_);
  nor (_14704_, _14590_, _07293_);
  or (_14705_, _14704_, _07292_);
  nand (_14706_, _14705_, _07334_);
  or (_14707_, _14705_, _07334_);
  and (_14708_, _14707_, _14706_);
  or (_14709_, _14708_, _07364_);
  nand (_14710_, _07364_, _07331_);
  and (_14711_, _14710_, _07010_);
  and (_14712_, _14711_, _14709_);
  or (_14713_, _14712_, _03903_);
  or (_14714_, _14713_, _14703_);
  and (_14715_, _14714_, _14646_);
  or (_14716_, _14715_, _03897_);
  and (_14717_, _12997_, _05440_);
  or (_14718_, _14643_, _04790_);
  or (_14719_, _14718_, _14717_);
  and (_14720_, _14719_, _04792_);
  and (_14721_, _14720_, _14716_);
  and (_14722_, _08741_, _05440_);
  or (_14723_, _14722_, _14643_);
  and (_14724_, _14723_, _04018_);
  or (_14725_, _14724_, _14721_);
  and (_14726_, _14725_, _03909_);
  or (_14727_, _14643_, _08336_);
  and (_14728_, _14645_, _03908_);
  and (_14729_, _14728_, _14727_);
  or (_14730_, _14729_, _14726_);
  and (_14731_, _14730_, _04785_);
  and (_14732_, _14658_, _04027_);
  and (_14733_, _14732_, _14727_);
  or (_14734_, _14733_, _03914_);
  or (_14735_, _14734_, _14731_);
  nor (_14736_, _12996_, _07937_);
  or (_14737_, _14643_, _06567_);
  or (_14738_, _14737_, _14736_);
  and (_14739_, _14738_, _06572_);
  and (_14740_, _14739_, _14735_);
  nor (_14741_, _08740_, _07937_);
  or (_14742_, _14741_, _14643_);
  and (_14743_, _14742_, _04011_);
  or (_14744_, _14743_, _03773_);
  or (_14745_, _14744_, _14740_);
  or (_14746_, _14655_, _03774_);
  and (_14747_, _14746_, _03375_);
  and (_14748_, _14747_, _14745_);
  and (_14749_, _14652_, _03374_);
  or (_14750_, _14749_, _03772_);
  or (_14751_, _14750_, _14748_);
  and (_14752_, _13056_, _05440_);
  or (_14753_, _14643_, _04060_);
  or (_14754_, _14753_, _14752_);
  and (_14755_, _14754_, _43152_);
  and (_14756_, _14755_, _14751_);
  or (_14757_, _14756_, _14642_);
  and (_43380_, _14757_, _41894_);
  nor (_14758_, _43152_, _07030_);
  nor (_14759_, _05440_, _07030_);
  nor (_14760_, _13182_, _07937_);
  or (_14761_, _14760_, _14759_);
  and (_14762_, _14761_, _03455_);
  nor (_14763_, _06088_, _07030_);
  and (_14764_, _13071_, _06088_);
  or (_14765_, _14764_, _14763_);
  and (_14766_, _14765_, _03759_);
  nor (_14767_, _13090_, _07937_);
  or (_14768_, _14767_, _14759_);
  or (_14769_, _14768_, _04722_);
  and (_14770_, _05440_, \oc8051_golden_model_1.ACC [5]);
  or (_14771_, _14770_, _14759_);
  and (_14772_, _14771_, _04707_);
  nor (_14773_, _04707_, _07030_);
  or (_14774_, _14773_, _03850_);
  or (_14775_, _14774_, _14772_);
  and (_14776_, _14775_, _03764_);
  and (_14777_, _14776_, _14769_);
  and (_14778_, _13094_, _06088_);
  or (_14779_, _14778_, _14763_);
  and (_14780_, _14779_, _03763_);
  or (_14781_, _14780_, _03848_);
  or (_14782_, _14781_, _14777_);
  and (_14783_, _05857_, _05440_);
  or (_14784_, _14783_, _14759_);
  or (_14785_, _14784_, _04733_);
  and (_14786_, _14785_, _14782_);
  or (_14787_, _14786_, _03854_);
  or (_14788_, _14771_, _03855_);
  and (_14789_, _14788_, _03760_);
  and (_14790_, _14789_, _14787_);
  or (_14791_, _14790_, _14766_);
  and (_14792_, _14791_, _03753_);
  or (_14793_, _14763_, _13109_);
  and (_14794_, _14793_, _03752_);
  and (_14795_, _14794_, _14779_);
  or (_14796_, _14795_, _07399_);
  or (_14797_, _14796_, _14792_);
  nor (_14798_, _07891_, _07597_);
  nor (_14799_, _14798_, _07892_);
  or (_14800_, _14799_, _07405_);
  and (_14801_, _14800_, _03747_);
  and (_14802_, _14801_, _14797_);
  nor (_14803_, _13073_, _07915_);
  or (_14804_, _14803_, _14763_);
  and (_14805_, _14804_, _03746_);
  or (_14806_, _14805_, _07927_);
  or (_14807_, _14806_, _14802_);
  and (_14808_, _06968_, _05440_);
  or (_14809_, _14759_, _03738_);
  or (_14810_, _14809_, _14808_);
  or (_14811_, _14784_, _07925_);
  and (_14812_, _14811_, _03820_);
  and (_14813_, _14812_, _14810_);
  and (_14814_, _14813_, _14807_);
  or (_14815_, _14814_, _14762_);
  and (_14816_, _14815_, _07011_);
  not (_14817_, _07341_);
  and (_14818_, _07364_, _07010_);
  and (_14819_, _14818_, _14817_);
  not (_14820_, _07333_);
  and (_14821_, _14706_, _14820_);
  nor (_14822_, _14821_, _07344_);
  and (_14823_, _14821_, _07344_);
  or (_14824_, _14823_, _14822_);
  nor (_14825_, _07364_, _07011_);
  and (_14826_, _14825_, _14824_);
  or (_14827_, _14826_, _14819_);
  or (_14828_, _14827_, _14816_);
  and (_14829_, _14828_, _04778_);
  and (_14830_, _06447_, _05440_);
  or (_14831_, _14830_, _14759_);
  and (_14832_, _14831_, _03903_);
  or (_14833_, _14832_, _03897_);
  or (_14834_, _14833_, _14829_);
  and (_14835_, _13196_, _05440_);
  or (_14836_, _14835_, _14759_);
  or (_14837_, _14836_, _04790_);
  and (_14838_, _14837_, _04792_);
  and (_14839_, _14838_, _14834_);
  and (_14840_, _10493_, _05440_);
  or (_14841_, _14840_, _14759_);
  and (_14842_, _14841_, _04018_);
  or (_14843_, _14842_, _14839_);
  and (_14844_, _14843_, _03909_);
  or (_14845_, _14759_, _08335_);
  and (_14846_, _14831_, _03908_);
  and (_14847_, _14846_, _14845_);
  or (_14848_, _14847_, _14844_);
  and (_14849_, _14848_, _04785_);
  and (_14850_, _14771_, _04027_);
  and (_14851_, _14850_, _14845_);
  or (_14852_, _14851_, _03914_);
  or (_14853_, _14852_, _14849_);
  nor (_14854_, _13195_, _07937_);
  or (_14855_, _14759_, _06567_);
  or (_14856_, _14855_, _14854_);
  and (_14857_, _14856_, _06572_);
  and (_14858_, _14857_, _14853_);
  nor (_14859_, _08738_, _07937_);
  or (_14860_, _14859_, _14759_);
  and (_14861_, _14860_, _04011_);
  or (_14862_, _14861_, _03773_);
  or (_14863_, _14862_, _14858_);
  or (_14864_, _14768_, _03774_);
  and (_14865_, _14864_, _03375_);
  and (_14866_, _14865_, _14863_);
  and (_14867_, _14765_, _03374_);
  or (_14868_, _14867_, _03772_);
  or (_14869_, _14868_, _14866_);
  and (_14870_, _13255_, _05440_);
  or (_14871_, _14759_, _04060_);
  or (_14872_, _14871_, _14870_);
  and (_14873_, _14872_, _43152_);
  and (_14874_, _14873_, _14869_);
  or (_14875_, _14874_, _14758_);
  and (_43381_, _14875_, _41894_);
  nor (_14876_, _43152_, _07275_);
  nor (_14877_, _05440_, _07275_);
  and (_14878_, _13394_, _05440_);
  or (_14879_, _14878_, _14877_);
  or (_14880_, _14879_, _04778_);
  nor (_14881_, _13387_, _07937_);
  or (_14882_, _14881_, _14877_);
  and (_14883_, _14882_, _03455_);
  nor (_14884_, _06088_, _07275_);
  and (_14885_, _13277_, _06088_);
  or (_14886_, _14885_, _14884_);
  and (_14887_, _14886_, _03759_);
  nor (_14888_, _13293_, _07937_);
  or (_14889_, _14888_, _14877_);
  or (_14890_, _14889_, _04722_);
  and (_14891_, _05440_, \oc8051_golden_model_1.ACC [6]);
  or (_14892_, _14891_, _14877_);
  and (_14893_, _14892_, _04707_);
  nor (_14894_, _04707_, _07275_);
  or (_14895_, _14894_, _03850_);
  or (_14896_, _14895_, _14893_);
  and (_14897_, _14896_, _03764_);
  and (_14898_, _14897_, _14890_);
  and (_14899_, _13297_, _06088_);
  or (_14900_, _14899_, _14884_);
  and (_14901_, _14900_, _03763_);
  or (_14902_, _14901_, _03848_);
  or (_14903_, _14902_, _14898_);
  and (_14904_, _06065_, _05440_);
  or (_14905_, _14904_, _14877_);
  or (_14906_, _14905_, _04733_);
  and (_14907_, _14906_, _14903_);
  or (_14908_, _14907_, _03854_);
  or (_14909_, _14892_, _03855_);
  and (_14910_, _14909_, _03760_);
  and (_14911_, _14910_, _14908_);
  or (_14912_, _14911_, _14887_);
  and (_14913_, _14912_, _03753_);
  or (_14914_, _14884_, _13312_);
  and (_14915_, _14900_, _03752_);
  and (_14916_, _14915_, _14914_);
  or (_14917_, _14916_, _07399_);
  or (_14918_, _14917_, _14913_);
  nor (_14919_, _07904_, _07893_);
  nor (_14920_, _14919_, _07905_);
  or (_14921_, _14920_, _07405_);
  and (_14922_, _14921_, _03747_);
  and (_14923_, _14922_, _14918_);
  nor (_14924_, _13279_, _07915_);
  or (_14925_, _14924_, _14884_);
  and (_14926_, _14925_, _03746_);
  or (_14927_, _14926_, _07927_);
  or (_14928_, _14927_, _14923_);
  and (_14929_, _06641_, _05440_);
  or (_14930_, _14877_, _03738_);
  or (_14931_, _14930_, _14929_);
  or (_14932_, _14905_, _07925_);
  and (_14933_, _14932_, _03820_);
  and (_14934_, _14933_, _14931_);
  and (_14935_, _14934_, _14928_);
  or (_14936_, _14935_, _14883_);
  and (_14937_, _14936_, _07011_);
  nor (_14938_, _14821_, _07342_);
  or (_14939_, _14938_, _07343_);
  and (_14940_, _14939_, _07324_);
  nor (_14941_, _14939_, _07324_);
  or (_14942_, _14941_, _14940_);
  or (_14943_, _14942_, _07364_);
  and (_14944_, _07281_, _07010_);
  or (_14945_, _14944_, _14825_);
  and (_14946_, _14945_, _14943_);
  or (_14947_, _14946_, _03903_);
  or (_14948_, _14947_, _14937_);
  and (_14949_, _14948_, _14880_);
  or (_14950_, _14949_, _03897_);
  and (_14951_, _13402_, _05440_);
  or (_14952_, _14951_, _14877_);
  or (_14953_, _14952_, _04790_);
  and (_14954_, _14953_, _04792_);
  and (_14955_, _14954_, _14950_);
  and (_14956_, _08736_, _05440_);
  or (_14957_, _14956_, _14877_);
  and (_14958_, _14957_, _04018_);
  or (_14959_, _14958_, _14955_);
  and (_14960_, _14959_, _03909_);
  or (_14961_, _14877_, _08322_);
  and (_14962_, _14879_, _03908_);
  and (_14963_, _14962_, _14961_);
  or (_14964_, _14963_, _14960_);
  and (_14965_, _14964_, _04785_);
  and (_14966_, _14892_, _04027_);
  and (_14967_, _14966_, _14961_);
  or (_14968_, _14967_, _03914_);
  or (_14969_, _14968_, _14965_);
  nor (_14970_, _13401_, _07937_);
  or (_14971_, _14877_, _06567_);
  or (_14972_, _14971_, _14970_);
  and (_14973_, _14972_, _06572_);
  and (_14974_, _14973_, _14969_);
  nor (_14975_, _08735_, _07937_);
  or (_14976_, _14975_, _14877_);
  and (_14977_, _14976_, _04011_);
  or (_14978_, _14977_, _03773_);
  or (_14979_, _14978_, _14974_);
  or (_14980_, _14889_, _03774_);
  and (_14981_, _14980_, _03375_);
  and (_14982_, _14981_, _14979_);
  and (_14983_, _14886_, _03374_);
  or (_14984_, _14983_, _03772_);
  or (_14985_, _14984_, _14982_);
  nor (_14986_, _13460_, _07937_);
  or (_14987_, _14877_, _04060_);
  or (_14988_, _14987_, _14986_);
  and (_14989_, _14988_, _43152_);
  and (_14990_, _14989_, _14985_);
  or (_14991_, _14990_, _14876_);
  and (_43382_, _14991_, _41894_);
  nor (_14992_, _43152_, _03498_);
  and (_14993_, _08820_, \oc8051_golden_model_1.ACC [1]);
  nand (_14994_, _08772_, _06554_);
  and (_14995_, _06733_, _03498_);
  nor (_14996_, _14995_, _08714_);
  or (_14997_, _14996_, _10058_);
  nand (_14998_, _08657_, _08297_);
  nor (_14999_, _08373_, _03498_);
  nor (_15000_, _14999_, _08374_);
  nand (_15001_, _15000_, _04022_);
  and (_15002_, _15001_, _08659_);
  nor (_15003_, _05429_, _03498_);
  nor (_15004_, _12177_, _08479_);
  nor (_15005_, _15004_, _15003_);
  nand (_15006_, _15005_, _03914_);
  nand (_15007_, _08573_, _14995_);
  and (_15008_, _08115_, _03392_);
  nor (_15009_, _04700_, \oc8051_golden_model_1.ACC [0]);
  nor (_15010_, _07919_, _04420_);
  nand (_15011_, _15010_, _15009_);
  or (_15012_, _08753_, _04026_);
  and (_15013_, _15012_, _08557_);
  and (_15014_, _08122_, _08022_);
  and (_15015_, _12178_, _05429_);
  nor (_15016_, _15015_, _15003_);
  nand (_15017_, _15016_, _03897_);
  not (_15018_, _10087_);
  nor (_15019_, _08094_, _03498_);
  nor (_15020_, _15019_, _08134_);
  nand (_15021_, _15020_, _08248_);
  and (_15022_, _15021_, _15018_);
  or (_15023_, _08157_, _04700_);
  nor (_15024_, _08159_, _04716_);
  or (_15025_, _15024_, _06962_);
  and (_15026_, _08169_, _04700_);
  or (_15027_, _04263_, \oc8051_golden_model_1.ACC [0]);
  nand (_15028_, _04263_, \oc8051_golden_model_1.ACC [0]);
  nand (_15029_, _15028_, _15027_);
  nor (_15030_, _15029_, _08169_);
  or (_15031_, _15030_, _08159_);
  or (_15032_, _15031_, _15026_);
  and (_15033_, _15032_, _03436_);
  or (_15034_, _15033_, _04716_);
  and (_15035_, _15034_, _04722_);
  and (_15036_, _15035_, _15025_);
  and (_15037_, _05716_, _05429_);
  nor (_15038_, _15037_, _15003_);
  nor (_15039_, _15038_, _04722_);
  or (_15040_, _15039_, _03763_);
  or (_15041_, _15040_, _15036_);
  nor (_15042_, _06096_, _03498_);
  and (_15043_, _12064_, _06096_);
  nor (_15044_, _15043_, _15042_);
  nand (_15045_, _15044_, _03763_);
  and (_15046_, _15045_, _04733_);
  and (_15047_, _15046_, _15041_);
  and (_15048_, _05429_, _04700_);
  nor (_15049_, _15048_, _15003_);
  nor (_15050_, _15049_, _04733_);
  or (_15051_, _15050_, _08212_);
  or (_15052_, _15051_, _15047_);
  and (_15053_, _15052_, _15023_);
  or (_15054_, _15053_, _04738_);
  or (_15055_, _06962_, _04739_);
  and (_15056_, _15055_, _03855_);
  and (_15057_, _15056_, _15054_);
  nor (_15058_, _05716_, _03855_);
  or (_15059_, _15058_, _08224_);
  or (_15060_, _15059_, _15057_);
  nand (_15061_, _08224_, _07090_);
  and (_15062_, _15061_, _15060_);
  or (_15063_, _15062_, _03759_);
  or (_15064_, _15003_, _03760_);
  and (_15065_, _15064_, _03753_);
  and (_15066_, _15065_, _15063_);
  nor (_15067_, _15038_, _03753_);
  or (_15068_, _15067_, _07399_);
  or (_15069_, _15068_, _15066_);
  not (_15070_, _07855_);
  and (_15071_, _07399_, _15070_);
  nor (_15072_, _15071_, _08148_);
  and (_15073_, _15072_, _11878_);
  and (_15074_, _15073_, _15069_);
  or (_15075_, _15074_, _15022_);
  nor (_15076_, _08299_, _03498_);
  nor (_15077_, _15076_, _08300_);
  nand (_15078_, _15077_, _04330_);
  and (_15079_, _15078_, _15075_);
  or (_15080_, _15079_, _03883_);
  nand (_15081_, _15000_, _03883_);
  and (_15082_, _15081_, _08321_);
  and (_15083_, _15082_, _15080_);
  nor (_15084_, _08441_, _03498_);
  nor (_15085_, _08442_, _15084_);
  nor (_15086_, _15085_, _08321_);
  or (_15087_, _15086_, _03425_);
  or (_15088_, _15087_, _15083_);
  nand (_15089_, _03715_, _03425_);
  and (_15090_, _15089_, _03747_);
  and (_15091_, _15090_, _15088_);
  nor (_15092_, _12104_, _08465_);
  or (_15093_, _15092_, _15042_);
  and (_15094_, _15093_, _03746_);
  or (_15095_, _15094_, _07927_);
  or (_15096_, _15095_, _15091_);
  and (_15097_, _06962_, _05429_);
  nor (_15098_, _15097_, _15003_);
  nand (_15099_, _15098_, _03737_);
  nand (_15100_, _15049_, _08474_);
  and (_15101_, _15100_, _03820_);
  and (_15102_, _15101_, _15099_);
  and (_15103_, _15102_, _15096_);
  nor (_15104_, _12164_, _08479_);
  nor (_15105_, _15104_, _15003_);
  nor (_15106_, _15105_, _03820_);
  or (_15107_, _15106_, _07010_);
  or (_15108_, _15107_, _15103_);
  nor (_15109_, _14818_, _03469_);
  and (_15110_, _15109_, _15108_);
  nor (_15111_, _03715_, _03479_);
  or (_15112_, _15111_, _03903_);
  or (_15113_, _15112_, _15110_);
  and (_15114_, _05429_, _06479_);
  nor (_15115_, _15114_, _15003_);
  nand (_15116_, _15115_, _03903_);
  and (_15117_, _15116_, _08493_);
  and (_15118_, _15117_, _15113_);
  nor (_15119_, _08493_, _03715_);
  or (_15120_, _15119_, _08503_);
  or (_15121_, _15120_, _15118_);
  nor (_15122_, _15009_, _08022_);
  or (_15123_, _08502_, _15122_);
  and (_15124_, _15123_, _08514_);
  and (_15125_, _15124_, _15121_);
  and (_15126_, _08515_, _15122_);
  or (_15127_, _15126_, _08519_);
  or (_15128_, _15127_, _15125_);
  or (_15129_, _14996_, _08520_);
  and (_15130_, _15129_, _15128_);
  or (_15131_, _15130_, _04016_);
  nand (_15132_, _10489_, _04016_);
  and (_15133_, _15132_, _08531_);
  and (_15134_, _15133_, _15131_);
  and (_15135_, _08530_, _10507_);
  or (_15136_, _15135_, _03897_);
  or (_15137_, _15136_, _15134_);
  and (_15138_, _15137_, _15017_);
  or (_15139_, _15138_, _04018_);
  or (_15140_, _15003_, _04792_);
  and (_15141_, _15140_, _08121_);
  and (_15142_, _15141_, _15139_);
  or (_15143_, _15142_, _15014_);
  and (_15144_, _15143_, _08548_);
  and (_15145_, _08547_, _08714_);
  or (_15146_, _15145_, _04025_);
  or (_15147_, _15146_, _15144_);
  and (_15148_, _15147_, _15013_);
  and (_15149_, _08553_, _08793_);
  or (_15150_, _15149_, _15148_);
  and (_15151_, _15150_, _03909_);
  nor (_15152_, _15115_, _15037_);
  and (_15153_, _15152_, _03908_);
  or (_15154_, _15153_, _15010_);
  or (_15155_, _15154_, _15151_);
  and (_15156_, _15155_, _15011_);
  or (_15157_, _15156_, _15008_);
  and (_15158_, _03831_, _03392_);
  not (_15159_, _15158_);
  nand (_15160_, _15008_, _15009_);
  and (_15161_, _15160_, _15159_);
  and (_15162_, _15161_, _15157_);
  nor (_15163_, _15009_, _15159_);
  or (_15164_, _15163_, _08573_);
  or (_15165_, _15164_, _15162_);
  and (_15166_, _15165_, _15007_);
  or (_15167_, _15166_, _04013_);
  nand (_15168_, _10488_, _04013_);
  and (_15169_, _15168_, _08583_);
  and (_15170_, _15169_, _15167_);
  nor (_15171_, _08583_, _10506_);
  or (_15172_, _15171_, _03914_);
  or (_15173_, _15172_, _15170_);
  and (_15174_, _15173_, _15006_);
  or (_15175_, _15174_, _08590_);
  nor (_15176_, _08597_, _15020_);
  or (_15177_, _15176_, _10061_);
  and (_15178_, _15177_, _15175_);
  nor (_15179_, _08599_, _15077_);
  or (_15180_, _15179_, _04022_);
  or (_15181_, _15180_, _15178_);
  and (_15182_, _15181_, _15002_);
  nor (_15183_, _08659_, _15085_);
  or (_15184_, _15183_, _08657_);
  or (_15185_, _15184_, _15182_);
  and (_15186_, _15185_, _14998_);
  or (_15187_, _15186_, _04206_);
  not (_15188_, _04206_);
  or (_15189_, _15122_, _15188_);
  nor (_15190_, _04621_, _04215_);
  and (_15191_, _15190_, _11983_);
  and (_15192_, _15191_, _11987_);
  and (_15193_, _15192_, _15189_);
  and (_15194_, _15193_, _15187_);
  not (_15195_, _15192_);
  and (_15196_, _15195_, _15122_);
  or (_15197_, _15196_, _08691_);
  or (_15198_, _15197_, _15194_);
  and (_15199_, _15198_, _14997_);
  or (_15200_, _15199_, _03779_);
  not (_15201_, _08733_);
  nand (_15202_, _10489_, _03779_);
  and (_15203_, _15202_, _15201_);
  and (_15204_, _15203_, _15200_);
  and (_15205_, _08733_, _10507_);
  or (_15206_, _15205_, _08772_);
  or (_15207_, _15206_, _15204_);
  and (_15208_, _15207_, _14994_);
  or (_15209_, _15208_, _03773_);
  nand (_15210_, _15038_, _03773_);
  and (_15211_, _15210_, _08816_);
  and (_15212_, _15211_, _15209_);
  and (_15213_, _08815_, _03498_);
  or (_15214_, _15213_, _15212_);
  and (_15215_, _15214_, _12016_);
  or (_15216_, _15215_, _14993_);
  and (_15217_, _15216_, _03375_);
  and (_15218_, _15003_, _03374_);
  or (_15219_, _15218_, _03772_);
  or (_15220_, _15219_, _15217_);
  nand (_15221_, _15038_, _03772_);
  and (_15222_, _15221_, _08838_);
  and (_15223_, _15222_, _15220_);
  nor (_15224_, _08844_, _03498_);
  nor (_15225_, _15224_, _10965_);
  or (_15226_, _15225_, _15223_);
  nand (_15227_, _08844_, _03474_);
  and (_15228_, _15227_, _43152_);
  and (_15229_, _15228_, _15226_);
  or (_15230_, _15229_, _14992_);
  and (_43383_, _15230_, _41894_);
  nor (_15231_, _43152_, _03474_);
  nand (_15232_, _08772_, _03498_);
  nor (_15233_, _08714_, _08713_);
  nor (_15234_, _15233_, _08715_);
  or (_15235_, _15234_, _10058_);
  and (_15236_, _08668_, _08666_);
  nor (_15237_, _15236_, _08669_);
  or (_15238_, _15237_, _08659_);
  nand (_15239_, _08573_, _08712_);
  nand (_15240_, _15010_, _08020_);
  and (_15241_, _08122_, _08019_);
  nor (_15242_, _05429_, _03474_);
  and (_15243_, _12366_, _05429_);
  nor (_15244_, _15243_, _15242_);
  nand (_15245_, _15244_, _03897_);
  and (_15246_, \oc8051_golden_model_1.PSW [7], _03498_);
  and (_15247_, _08297_, \oc8051_golden_model_1.ACC [0]);
  not (_15248_, _15247_);
  and (_15249_, _15248_, _06962_);
  nor (_15250_, _15249_, _15246_);
  and (_15251_, _15250_, _08713_);
  nor (_15252_, _15250_, _08713_);
  or (_15253_, _15252_, _15251_);
  or (_15254_, _15253_, _08248_);
  or (_15255_, _08157_, _04900_);
  or (_15256_, _15024_, _06961_);
  and (_15257_, _08169_, _04900_);
  or (_15258_, _04263_, \oc8051_golden_model_1.ACC [1]);
  nand (_15259_, _04263_, \oc8051_golden_model_1.ACC [1]);
  nand (_15260_, _15259_, _15258_);
  nor (_15261_, _15260_, _08169_);
  or (_15262_, _15261_, _08159_);
  or (_15263_, _15262_, _15257_);
  and (_15264_, _15263_, _03436_);
  or (_15265_, _15264_, _04716_);
  and (_15266_, _15265_, _15256_);
  or (_15267_, _15266_, _03850_);
  nor (_15268_, _05429_, \oc8051_golden_model_1.ACC [1]);
  and (_15269_, _12262_, _05429_);
  nor (_15270_, _15269_, _15268_);
  or (_15271_, _15270_, _04722_);
  and (_15272_, _15271_, _15267_);
  or (_15273_, _15272_, _08179_);
  nor (_15274_, _08186_, \oc8051_golden_model_1.PSW [6]);
  nor (_15275_, _15274_, \oc8051_golden_model_1.ACC [1]);
  and (_15276_, _15274_, \oc8051_golden_model_1.ACC [1]);
  nor (_15277_, _15276_, _15275_);
  nand (_15278_, _15277_, _08179_);
  and (_15279_, _15278_, _03856_);
  and (_15280_, _15279_, _15273_);
  nor (_15281_, _06096_, _03474_);
  and (_15282_, _12249_, _06096_);
  nor (_15283_, _15282_, _15281_);
  nor (_15284_, _15283_, _03764_);
  and (_15285_, _05429_, _04900_);
  nor (_15286_, _15285_, _15242_);
  nor (_15287_, _15286_, _04733_);
  or (_15288_, _15287_, _08212_);
  or (_15289_, _15288_, _15284_);
  or (_15290_, _15289_, _15280_);
  and (_15291_, _15290_, _15255_);
  or (_15292_, _15291_, _04738_);
  or (_15293_, _06961_, _04739_);
  and (_15294_, _15293_, _03855_);
  and (_15295_, _15294_, _15292_);
  nor (_15296_, _05669_, _03855_);
  or (_15297_, _15296_, _08224_);
  or (_15298_, _15297_, _15295_);
  nand (_15299_, _08224_, _07084_);
  and (_15300_, _15299_, _15298_);
  or (_15301_, _15300_, _03759_);
  and (_15302_, _12252_, _06096_);
  nor (_15303_, _15302_, _15281_);
  nand (_15304_, _15303_, _03759_);
  and (_15305_, _15304_, _03753_);
  and (_15306_, _15305_, _15301_);
  and (_15307_, _15282_, _12248_);
  nor (_15308_, _15307_, _15281_);
  nor (_15309_, _15308_, _03753_);
  or (_15310_, _15309_, _07399_);
  or (_15311_, _15310_, _15306_);
  and (_15312_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_15313_, _15312_, _07306_);
  nor (_15314_, _15313_, _07856_);
  or (_15315_, _15314_, _07405_);
  and (_15316_, _15315_, _08153_);
  and (_15317_, _15316_, _15311_);
  and (_15318_, _15248_, _04700_);
  nor (_15319_, _15318_, _15246_);
  and (_15320_, _15319_, _08021_);
  nor (_15321_, _15319_, _08021_);
  or (_15322_, _15321_, _15320_);
  or (_15323_, _15322_, _04330_);
  and (_15324_, _15323_, _15018_);
  or (_15325_, _15324_, _15317_);
  and (_15326_, _15325_, _15254_);
  or (_15327_, _15326_, _03883_);
  nor (_15328_, _15247_, _05716_);
  nor (_15329_, _15328_, _15246_);
  and (_15330_, _15329_, _08752_);
  nor (_15331_, _15329_, _08752_);
  or (_15332_, _15331_, _15330_);
  or (_15333_, _15332_, _03888_);
  and (_15334_, _15333_, _08321_);
  and (_15335_, _15334_, _15327_);
  nor (_15336_, _15247_, _03715_);
  nor (_15337_, _15336_, _15246_);
  and (_15338_, _15337_, _08792_);
  nor (_15339_, _15337_, _08792_);
  nor (_15340_, _15339_, _15338_);
  nor (_15341_, _15340_, _08321_);
  or (_15342_, _15341_, _03425_);
  or (_15343_, _15342_, _15335_);
  nand (_15344_, _04563_, _03425_);
  and (_15345_, _15344_, _03747_);
  and (_15346_, _15345_, _15343_);
  nor (_15347_, _12293_, _08465_);
  nor (_15348_, _15347_, _15281_);
  nor (_15349_, _15348_, _03747_);
  or (_15350_, _15349_, _07927_);
  or (_15351_, _15350_, _15346_);
  and (_15352_, _06961_, _05429_);
  nor (_15353_, _15352_, _15242_);
  nand (_15354_, _15353_, _03737_);
  nand (_15355_, _15286_, _08474_);
  and (_15356_, _15355_, _03820_);
  and (_15357_, _15356_, _15354_);
  and (_15358_, _15357_, _15351_);
  nor (_15359_, _12352_, _08479_);
  nor (_15360_, _15359_, _15242_);
  nor (_15361_, _15360_, _03820_);
  or (_15362_, _15361_, _07010_);
  or (_15363_, _15362_, _15358_);
  or (_15364_, _07269_, _07011_);
  and (_15365_, _15364_, _03479_);
  and (_15366_, _15365_, _15363_);
  nor (_15367_, _04563_, _03479_);
  or (_15368_, _15367_, _03903_);
  or (_15369_, _15368_, _15366_);
  and (_15370_, _05429_, _04595_);
  nor (_15371_, _15370_, _15268_);
  or (_15372_, _15371_, _04778_);
  and (_15373_, _15372_, _08493_);
  and (_15374_, _15373_, _15369_);
  nor (_15375_, _08493_, _04563_);
  or (_15376_, _15375_, _08503_);
  or (_15377_, _15376_, _15374_);
  or (_15378_, _08502_, _08021_);
  and (_15379_, _15378_, _08508_);
  and (_15380_, _15379_, _15377_);
  not (_15381_, _08508_);
  and (_15382_, _15381_, _08021_);
  or (_15383_, _15382_, _08512_);
  or (_15384_, _15383_, _15380_);
  or (_15385_, _08513_, _08021_);
  and (_15386_, _15385_, _08520_);
  and (_15387_, _15386_, _15384_);
  and (_15388_, _08713_, _08519_);
  or (_15389_, _15388_, _04016_);
  or (_15390_, _15389_, _15387_);
  or (_15391_, _08752_, _04017_);
  and (_15392_, _15391_, _08531_);
  and (_15393_, _15392_, _15390_);
  and (_15394_, _08530_, _08792_);
  or (_15395_, _15394_, _03897_);
  or (_15396_, _15395_, _15393_);
  and (_15397_, _15396_, _15245_);
  or (_15398_, _15397_, _04018_);
  or (_15399_, _15242_, _04792_);
  and (_15400_, _15399_, _08121_);
  and (_15401_, _15400_, _15398_);
  or (_15402_, _15401_, _15241_);
  and (_15403_, _15402_, _08548_);
  and (_15404_, _08547_, _08711_);
  or (_15405_, _15404_, _04025_);
  or (_15406_, _15405_, _15403_);
  or (_15407_, _08750_, _04026_);
  and (_15408_, _15407_, _08557_);
  and (_15409_, _15408_, _15406_);
  and (_15410_, _08553_, _08790_);
  or (_15411_, _15410_, _15409_);
  and (_15412_, _15411_, _03909_);
  and (_15413_, _12244_, _05429_);
  nor (_15414_, _15413_, _15242_);
  nor (_15415_, _15414_, _03909_);
  or (_15416_, _15415_, _15010_);
  or (_15417_, _15416_, _15412_);
  and (_15418_, _15417_, _15240_);
  or (_15419_, _15418_, _15008_);
  nand (_15420_, _07922_, _03392_);
  nor (_15421_, _08020_, _15158_);
  or (_15422_, _15421_, _15420_);
  and (_15423_, _15422_, _15419_);
  nor (_15424_, _08020_, _15159_);
  or (_15425_, _15424_, _08573_);
  or (_15426_, _15425_, _15423_);
  and (_15427_, _15426_, _15239_);
  or (_15428_, _15427_, _04013_);
  nand (_15429_, _08751_, _04013_);
  and (_15430_, _15429_, _08583_);
  and (_15431_, _15430_, _15428_);
  nor (_15432_, _08583_, _08791_);
  or (_15433_, _15432_, _03914_);
  or (_15434_, _15433_, _15431_);
  nor (_15435_, _12365_, _08479_);
  or (_15436_, _15435_, _15242_);
  or (_15437_, _15436_, _06567_);
  and (_15438_, _15437_, _08119_);
  and (_15439_, _15438_, _15434_);
  and (_15440_, _08096_, _08092_);
  nor (_15441_, _15440_, _08097_);
  or (_15442_, _15441_, _08597_);
  and (_15443_, _15442_, _10688_);
  or (_15444_, _15443_, _15439_);
  and (_15445_, _08608_, _08606_);
  nor (_15446_, _15445_, _08609_);
  or (_15447_, _15446_, _08599_);
  and (_15448_, _15447_, _04023_);
  and (_15449_, _15448_, _15444_);
  and (_15450_, _08638_, _08636_);
  nor (_15451_, _15450_, _08639_);
  and (_15452_, _15451_, _04022_);
  or (_15453_, _15452_, _08627_);
  or (_15454_, _15453_, _15449_);
  and (_15455_, _15454_, _15238_);
  or (_15456_, _15455_, _08657_);
  nand (_15457_, _08657_, _03498_);
  and (_15458_, _15457_, _07999_);
  and (_15459_, _15458_, _15456_);
  not (_15460_, _07999_);
  nor (_15461_, _08022_, _08021_);
  nor (_15462_, _15461_, _08023_);
  and (_15463_, _15462_, _15460_);
  or (_15464_, _15463_, _08691_);
  or (_15465_, _15464_, _15459_);
  and (_15466_, _15465_, _15235_);
  or (_15467_, _15466_, _03779_);
  nor (_15468_, _08753_, _08752_);
  nor (_15469_, _15468_, _08754_);
  or (_15470_, _15469_, _04140_);
  and (_15471_, _15470_, _15201_);
  and (_15472_, _15471_, _15467_);
  nor (_15473_, _08793_, _08792_);
  nor (_15474_, _15473_, _08794_);
  and (_15475_, _15474_, _08733_);
  or (_15476_, _15475_, _08772_);
  or (_15477_, _15476_, _15472_);
  and (_15478_, _15477_, _15232_);
  or (_15479_, _15478_, _03773_);
  or (_15480_, _15270_, _03774_);
  and (_15481_, _15480_, _08816_);
  and (_15482_, _15481_, _15479_);
  nor (_15483_, _08845_, _08821_);
  nor (_15484_, _15483_, _08816_);
  or (_15485_, _15484_, _08820_);
  or (_15486_, _15485_, _15482_);
  nand (_15487_, _08820_, _07190_);
  and (_15488_, _15487_, _03375_);
  and (_15489_, _15488_, _15486_);
  nor (_15490_, _15303_, _03375_);
  or (_15491_, _15490_, _03772_);
  or (_15492_, _15491_, _15489_);
  nor (_15493_, _15269_, _15242_);
  nand (_15494_, _15493_, _03772_);
  and (_15495_, _15494_, _08838_);
  and (_15496_, _15495_, _15492_);
  nor (_15497_, _15483_, _08844_);
  nor (_15498_, _15497_, _10965_);
  or (_15499_, _15498_, _15496_);
  nand (_15500_, _08844_, _07190_);
  and (_15501_, _15500_, _43152_);
  and (_15502_, _15501_, _15499_);
  or (_15503_, _15502_, _15231_);
  and (_43384_, _15503_, _41894_);
  nor (_15504_, _43152_, _07190_);
  nand (_15505_, _08772_, _03474_);
  and (_15506_, _08640_, _08364_);
  nor (_15507_, _15506_, _08641_);
  or (_15508_, _15507_, _04023_);
  and (_15509_, _15508_, _08659_);
  nand (_15510_, _08573_, _08708_);
  nand (_15511_, _15010_, _08016_);
  and (_15512_, _08115_, _03387_);
  not (_15513_, _08153_);
  or (_15514_, _08157_, _05307_);
  or (_15515_, _15024_, _06965_);
  and (_15516_, _08169_, _05307_);
  or (_15517_, _04263_, \oc8051_golden_model_1.ACC [2]);
  nand (_15518_, _04263_, \oc8051_golden_model_1.ACC [2]);
  nand (_15519_, _15518_, _15517_);
  nor (_15520_, _15519_, _08169_);
  or (_15521_, _15520_, _08159_);
  or (_15522_, _15521_, _15516_);
  and (_15523_, _15522_, _03436_);
  or (_15524_, _15523_, _04716_);
  and (_15525_, _15524_, _15515_);
  and (_15526_, _15525_, _04722_);
  nor (_15527_, _05429_, _07190_);
  nor (_15528_, _12471_, _08479_);
  nor (_15529_, _15528_, _15527_);
  nor (_15530_, _15529_, _04722_);
  or (_15531_, _15530_, _08179_);
  or (_15532_, _15531_, _15526_);
  nand (_15533_, _15274_, \oc8051_golden_model_1.ACC [2]);
  and (_15534_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_15535_, _15534_, _08185_);
  or (_15536_, _15535_, _15274_);
  and (_15537_, _15536_, _15533_);
  nand (_15538_, _15537_, _08179_);
  and (_15539_, _15538_, _03856_);
  and (_15540_, _15539_, _15532_);
  nor (_15541_, _06096_, _07190_);
  and (_15542_, _12464_, _06096_);
  nor (_15543_, _15542_, _15541_);
  nor (_15544_, _15543_, _03764_);
  and (_15545_, _05429_, _05307_);
  nor (_15546_, _15545_, _15527_);
  nor (_15547_, _15546_, _04733_);
  or (_15548_, _15547_, _08212_);
  or (_15549_, _15548_, _15544_);
  or (_15550_, _15549_, _15540_);
  and (_15551_, _15550_, _15514_);
  or (_15552_, _15551_, _04738_);
  or (_15553_, _06965_, _04739_);
  and (_15554_, _15553_, _03855_);
  and (_15555_, _15554_, _15552_);
  nor (_15556_, _05764_, _03855_);
  or (_15557_, _15556_, _08224_);
  or (_15558_, _15557_, _15555_);
  nand (_15559_, _08224_, _07036_);
  and (_15560_, _15559_, _15558_);
  or (_15561_, _15560_, _03759_);
  and (_15562_, _12467_, _06096_);
  nor (_15563_, _15562_, _15541_);
  nand (_15564_, _15563_, _03759_);
  and (_15565_, _15564_, _03753_);
  and (_15566_, _15565_, _15561_);
  and (_15567_, _15542_, _12463_);
  nor (_15568_, _15567_, _15541_);
  nor (_15569_, _15568_, _03753_);
  or (_15570_, _15569_, _07399_);
  or (_15571_, _15570_, _15566_);
  nor (_15572_, _07858_, _07856_);
  nor (_15573_, _15572_, _07859_);
  or (_15574_, _15573_, _07405_);
  and (_15575_, _15574_, _15571_);
  or (_15576_, _15575_, _15513_);
  nor (_15577_, _04900_, _03474_);
  and (_15578_, _04700_, _03498_);
  nor (_15579_, _15578_, _08021_);
  nor (_15580_, _15579_, _15577_);
  nor (_15581_, _15580_, _08017_);
  and (_15582_, _15580_, _08017_);
  nor (_15583_, _15582_, _15581_);
  nor (_15584_, _15122_, _08021_);
  not (_15585_, _15584_);
  or (_15586_, _15585_, _15583_);
  and (_15587_, _15586_, \oc8051_golden_model_1.PSW [7]);
  nor (_15588_, _15583_, \oc8051_golden_model_1.PSW [7]);
  or (_15589_, _15588_, _15587_);
  nand (_15590_, _15585_, _15583_);
  and (_15591_, _15590_, _15589_);
  nand (_15592_, _15591_, _15513_);
  and (_15593_, _15592_, _08248_);
  and (_15594_, _15593_, _15576_);
  and (_15595_, _06688_, \oc8051_golden_model_1.ACC [1]);
  and (_15596_, _06962_, _03498_);
  nor (_15597_, _15596_, _08713_);
  nor (_15598_, _15597_, _15595_);
  nor (_15599_, _08709_, _15598_);
  and (_15600_, _08709_, _15598_);
  nor (_15601_, _15600_, _15599_);
  nor (_15602_, _14996_, _08713_);
  not (_15603_, _15602_);
  or (_15604_, _15603_, _15601_);
  and (_15605_, _15604_, \oc8051_golden_model_1.PSW [7]);
  nor (_15606_, _15601_, \oc8051_golden_model_1.PSW [7]);
  or (_15607_, _15606_, _15605_);
  nand (_15608_, _15603_, _15601_);
  and (_15609_, _15608_, _15607_);
  nor (_15610_, _15609_, _08248_);
  or (_15611_, _15610_, _10086_);
  or (_15612_, _15611_, _15594_);
  and (_15613_, _05669_, \oc8051_golden_model_1.ACC [1]);
  nor (_15614_, _05716_, \oc8051_golden_model_1.ACC [0]);
  nor (_15615_, _11803_, _15614_);
  nor (_15616_, _15615_, _15613_);
  nor (_15617_, _08748_, _15616_);
  and (_15618_, _08748_, _15616_);
  nor (_15619_, _15618_, _15617_);
  not (_15620_, _15619_);
  and (_15621_, _10490_, \oc8051_golden_model_1.PSW [7]);
  and (_15622_, _15621_, _15620_);
  nor (_15623_, _15621_, _15620_);
  nor (_15624_, _15623_, _15622_);
  nand (_15625_, _15624_, _03883_);
  nor (_15626_, _03715_, \oc8051_golden_model_1.ACC [0]);
  nor (_15627_, _15626_, _08792_);
  nor (_15628_, _15627_, _11844_);
  nor (_15629_, _08788_, _15628_);
  and (_15630_, _08788_, _15628_);
  nor (_15631_, _15630_, _15629_);
  not (_15632_, _10508_);
  or (_15633_, _15632_, _15631_);
  and (_15634_, _15633_, \oc8051_golden_model_1.PSW [7]);
  nor (_15635_, _15631_, \oc8051_golden_model_1.PSW [7]);
  or (_15636_, _15635_, _15634_);
  nand (_15637_, _15632_, _15631_);
  and (_15638_, _15637_, _15636_);
  nand (_15639_, _15638_, _08320_);
  and (_15640_, _15639_, _15625_);
  and (_15641_, _15640_, _15612_);
  or (_15642_, _15641_, _03425_);
  nand (_15643_, _04139_, _03425_);
  and (_15644_, _15643_, _03747_);
  and (_15645_, _15644_, _15642_);
  nor (_15646_, _12514_, _08465_);
  nor (_15647_, _15646_, _15541_);
  nor (_15648_, _15647_, _03747_);
  or (_15649_, _15648_, _07927_);
  or (_15650_, _15649_, _15645_);
  and (_15651_, _06965_, _05429_);
  nor (_15652_, _15651_, _15527_);
  nand (_15653_, _15652_, _03737_);
  nand (_15654_, _15546_, _08474_);
  and (_15655_, _15654_, _03820_);
  and (_15656_, _15655_, _15653_);
  and (_15657_, _15656_, _15650_);
  nor (_15658_, _12572_, _08479_);
  nor (_15659_, _15658_, _15527_);
  nor (_15660_, _15659_, _03820_);
  or (_15661_, _15660_, _07010_);
  or (_15662_, _15661_, _15657_);
  or (_15663_, _07204_, _07011_);
  and (_15664_, _15663_, _03479_);
  and (_15665_, _15664_, _15662_);
  nor (_15666_, _04139_, _03479_);
  or (_15667_, _15666_, _03903_);
  or (_15668_, _15667_, _15665_);
  and (_15669_, _05429_, _06495_);
  nor (_15670_, _15669_, _15527_);
  nand (_15671_, _15670_, _03903_);
  and (_15672_, _15671_, _08493_);
  and (_15673_, _15672_, _15668_);
  nor (_15674_, _08493_, _04139_);
  or (_15675_, _15674_, _08503_);
  or (_15676_, _15675_, _15673_);
  or (_15677_, _08502_, _08017_);
  and (_15678_, _03825_, _03404_);
  not (_15679_, _15678_);
  and (_15680_, _15679_, _08508_);
  and (_15681_, _15680_, _15677_);
  and (_15682_, _15681_, _15676_);
  nor (_15683_, _15680_, _08018_);
  or (_15684_, _15683_, _04397_);
  or (_15685_, _15684_, _15682_);
  nand (_15686_, _08018_, _04397_);
  and (_15687_, _15686_, _08520_);
  and (_15688_, _15687_, _15685_);
  and (_15689_, _08709_, _08519_);
  or (_15690_, _15689_, _04016_);
  or (_15691_, _15690_, _15688_);
  or (_15692_, _08748_, _04017_);
  and (_15693_, _15692_, _15691_);
  and (_15694_, _15693_, _08531_);
  and (_15695_, _08530_, _08788_);
  or (_15696_, _15695_, _03897_);
  or (_15697_, _15696_, _15694_);
  and (_15698_, _12586_, _05429_);
  or (_15699_, _15698_, _15527_);
  or (_15700_, _15699_, _04790_);
  and (_15701_, _15700_, _04792_);
  and (_15702_, _15701_, _15697_);
  not (_15703_, _03387_);
  nor (_15704_, _07919_, _15703_);
  and (_15705_, _15527_, _04018_);
  or (_15706_, _15705_, _15704_);
  or (_15707_, _15706_, _15702_);
  not (_15708_, _08015_);
  nand (_15709_, _15704_, _15708_);
  and (_15710_, _15709_, _15707_);
  or (_15711_, _15710_, _15512_);
  nand (_15712_, _15512_, _15708_);
  and (_15713_, _15712_, _15711_);
  or (_15714_, _15713_, _04409_);
  not (_15715_, _04409_);
  or (_15716_, _08015_, _15715_);
  and (_15717_, _15716_, _08548_);
  and (_15718_, _15717_, _15714_);
  and (_15719_, _08547_, _08707_);
  or (_15720_, _15719_, _04025_);
  or (_15721_, _15720_, _15718_);
  or (_15722_, _08746_, _04026_);
  and (_15723_, _15722_, _15721_);
  or (_15724_, _15723_, _08553_);
  or (_15725_, _08557_, _08786_);
  and (_15726_, _15725_, _03909_);
  and (_15727_, _15726_, _15724_);
  or (_15728_, _15670_, _08747_);
  nor (_15729_, _15728_, _03909_);
  or (_15730_, _15729_, _15010_);
  or (_15731_, _15730_, _15727_);
  and (_15732_, _15731_, _15511_);
  or (_15733_, _15732_, _15008_);
  nor (_15734_, _08016_, _15158_);
  or (_15735_, _15734_, _15420_);
  and (_15736_, _15735_, _15733_);
  nor (_15737_, _08016_, _15159_);
  or (_15738_, _15737_, _08573_);
  or (_15739_, _15738_, _15736_);
  and (_15740_, _15739_, _15510_);
  or (_15741_, _15740_, _04013_);
  nand (_15742_, _08747_, _04013_);
  and (_15743_, _15742_, _08583_);
  and (_15744_, _15743_, _15741_);
  nor (_15745_, _08583_, _08787_);
  or (_15746_, _15745_, _03914_);
  or (_15747_, _15746_, _15744_);
  nor (_15748_, _12585_, _08479_);
  nor (_15749_, _15748_, _15527_);
  nand (_15750_, _15749_, _03914_);
  and (_15751_, _15750_, _08119_);
  and (_15752_, _15751_, _15747_);
  and (_15753_, _08098_, _08085_);
  nor (_15754_, _15753_, _08099_);
  and (_15755_, _15754_, _08590_);
  or (_15756_, _15755_, _15752_);
  and (_15757_, _15756_, _08599_);
  and (_15758_, _08610_, _08290_);
  nor (_15759_, _15758_, _08611_);
  and (_15760_, _15759_, _08597_);
  or (_15761_, _15760_, _04022_);
  or (_15762_, _15761_, _15757_);
  and (_15763_, _15762_, _15509_);
  and (_15764_, _08670_, _08433_);
  nor (_15765_, _15764_, _08671_);
  and (_15766_, _15765_, _08627_);
  or (_15767_, _15766_, _08657_);
  or (_15768_, _15767_, _15763_);
  nand (_15769_, _08657_, _03474_);
  and (_15770_, _15769_, _07999_);
  and (_15771_, _15770_, _15768_);
  and (_15772_, _08024_, _08018_);
  nor (_15773_, _15772_, _08025_);
  and (_15774_, _15773_, _15460_);
  or (_15775_, _15774_, _15771_);
  and (_15776_, _15775_, _10058_);
  and (_15777_, _08716_, _08710_);
  nor (_15778_, _15777_, _08717_);
  and (_15779_, _15778_, _08691_);
  or (_15780_, _15779_, _03779_);
  or (_15781_, _15780_, _15776_);
  and (_15782_, _08755_, _08749_);
  nor (_15783_, _15782_, _08756_);
  or (_15784_, _15783_, _04140_);
  and (_15785_, _15784_, _15201_);
  and (_15786_, _15785_, _15781_);
  and (_15787_, _08795_, _08789_);
  nor (_15788_, _15787_, _08796_);
  and (_15789_, _15788_, _08733_);
  or (_15790_, _15789_, _08772_);
  or (_15791_, _15790_, _15786_);
  and (_15792_, _15791_, _15505_);
  or (_15793_, _15792_, _03773_);
  nand (_15794_, _15529_, _03773_);
  and (_15795_, _15794_, _08816_);
  and (_15796_, _15795_, _15793_);
  and (_15797_, _08185_, _03498_);
  nor (_15798_, _08821_, _07190_);
  or (_15799_, _15798_, _15797_);
  and (_15800_, _15799_, _08815_);
  or (_15801_, _15800_, _08820_);
  or (_15802_, _15801_, _15796_);
  nand (_15803_, _08820_, _07184_);
  and (_15804_, _15803_, _03375_);
  and (_15805_, _15804_, _15802_);
  nor (_15806_, _15563_, _03375_);
  or (_15807_, _15806_, _03772_);
  or (_15808_, _15807_, _15805_);
  and (_15809_, _12642_, _05429_);
  nor (_15810_, _15809_, _15527_);
  nand (_15811_, _15810_, _03772_);
  and (_15812_, _15811_, _08838_);
  and (_15813_, _15812_, _15808_);
  and (_15814_, _08845_, \oc8051_golden_model_1.ACC [2]);
  nor (_15815_, _08845_, \oc8051_golden_model_1.ACC [2]);
  nor (_15816_, _15815_, _15814_);
  nor (_15817_, _15816_, _08844_);
  nor (_15818_, _15817_, _10965_);
  or (_15819_, _15818_, _15813_);
  nand (_15820_, _08844_, _07184_);
  and (_15821_, _15820_, _43152_);
  and (_15822_, _15821_, _15819_);
  or (_15823_, _15822_, _15504_);
  and (_43385_, _15823_, _41894_);
  nor (_15824_, _43152_, _07184_);
  nor (_15825_, _08014_, _08013_);
  nor (_15826_, _15825_, _08026_);
  and (_15827_, _15825_, _08026_);
  nor (_15828_, _15827_, _15826_);
  nand (_15829_, _15828_, _15460_);
  nor (_15830_, _05429_, _07184_);
  nor (_15831_, _12788_, _08479_);
  nor (_15832_, _15831_, _15830_);
  nor (_15833_, _15832_, _06567_);
  nand (_15834_, _08568_, _08014_);
  and (_15835_, _12789_, _05429_);
  nor (_15836_, _15835_, _15830_);
  nand (_15837_, _15836_, _03897_);
  nor (_15838_, _08493_, _03678_);
  and (_15839_, _06824_, \oc8051_golden_model_1.ACC [2]);
  nor (_15840_, _15599_, _15839_);
  nor (_15841_, _08706_, _08705_);
  nor (_15842_, _15841_, _15840_);
  and (_15843_, _15841_, _15840_);
  nor (_15844_, _15843_, _15842_);
  and (_15845_, _15844_, \oc8051_golden_model_1.PSW [7]);
  nor (_15846_, _15844_, \oc8051_golden_model_1.PSW [7]);
  nor (_15847_, _15846_, _15845_);
  and (_15848_, _15847_, _15605_);
  nor (_15849_, _15847_, _15605_);
  or (_15850_, _15849_, _15848_);
  nand (_15851_, _15850_, _04330_);
  nor (_15852_, _07861_, _07859_);
  nor (_15853_, _15852_, _07862_);
  and (_15854_, _15853_, _07399_);
  nor (_15855_, _06096_, _07184_);
  and (_15856_, _12674_, _06096_);
  and (_15857_, _15856_, _12673_);
  nor (_15858_, _15857_, _15855_);
  nor (_15859_, _15858_, _03753_);
  or (_15860_, _08157_, _05119_);
  or (_15861_, _10400_, _05119_);
  nor (_15862_, _04263_, _07184_);
  and (_15863_, _04263_, _07184_);
  or (_15864_, _15863_, _15862_);
  or (_15865_, _15864_, _08169_);
  and (_15866_, _15865_, _08160_);
  and (_15867_, _15866_, _15861_);
  and (_15868_, _15867_, _04717_);
  or (_15869_, _15868_, _06964_);
  or (_15870_, _15867_, _08159_);
  and (_15871_, _15870_, _03436_);
  or (_15872_, _15871_, _04716_);
  and (_15873_, _15872_, _04722_);
  and (_15874_, _15873_, _15869_);
  nor (_15875_, _12681_, _08479_);
  nor (_15876_, _15875_, _15830_);
  nor (_15877_, _15876_, _04722_);
  or (_15878_, _15877_, _08179_);
  or (_15879_, _15878_, _15874_);
  not (_15880_, \oc8051_golden_model_1.PSW [6]);
  nor (_15881_, _08185_, _15880_);
  nor (_15882_, _15881_, \oc8051_golden_model_1.ACC [3]);
  or (_15883_, _15882_, _08186_);
  nand (_15884_, _15883_, _08179_);
  and (_15885_, _15884_, _15879_);
  or (_15886_, _15885_, _03763_);
  nor (_15887_, _15856_, _15855_);
  nand (_15888_, _15887_, _03763_);
  and (_15889_, _15888_, _04733_);
  and (_15890_, _15889_, _15886_);
  and (_15891_, _05429_, _05119_);
  nor (_15892_, _15891_, _15830_);
  nor (_15893_, _15892_, _04733_);
  or (_15894_, _15893_, _08212_);
  or (_15895_, _15894_, _15890_);
  and (_15896_, _15895_, _15860_);
  or (_15897_, _15896_, _04738_);
  or (_15898_, _06964_, _04739_);
  and (_15899_, _15898_, _03855_);
  and (_15900_, _15899_, _15897_);
  nor (_15901_, _05621_, _03855_);
  or (_15902_, _15901_, _08224_);
  or (_15903_, _15902_, _15900_);
  nand (_15904_, _08224_, _06554_);
  and (_15905_, _15904_, _15903_);
  or (_15906_, _15905_, _03759_);
  and (_15907_, _12667_, _06096_);
  nor (_15908_, _15907_, _15855_);
  nand (_15909_, _15908_, _03759_);
  and (_15910_, _15909_, _03753_);
  and (_15911_, _15910_, _15906_);
  or (_15912_, _15911_, _15859_);
  and (_15913_, _15912_, _07405_);
  or (_15914_, _15913_, _11880_);
  or (_15915_, _15914_, _15854_);
  nor (_15916_, _05307_, _07190_);
  nor (_15917_, _15581_, _15916_);
  nor (_15918_, _15917_, _15825_);
  and (_15919_, _15917_, _15825_);
  nor (_15920_, _15919_, _15918_);
  and (_15921_, _15920_, \oc8051_golden_model_1.PSW [7]);
  nor (_15922_, _15920_, \oc8051_golden_model_1.PSW [7]);
  nor (_15923_, _15922_, _15921_);
  and (_15924_, _15923_, _15587_);
  nor (_15925_, _15923_, _15587_);
  or (_15926_, _15925_, _15924_);
  nand (_15927_, _15926_, _11880_);
  and (_15928_, _15927_, _11883_);
  and (_15929_, _15928_, _15915_);
  nor (_15930_, _15926_, _11883_);
  or (_15931_, _15930_, _04330_);
  or (_15932_, _15931_, _15929_);
  and (_15933_, _15932_, _15851_);
  or (_15934_, _15933_, _03883_);
  nand (_15935_, _10490_, _15620_);
  and (_15936_, _15935_, \oc8051_golden_model_1.PSW [7]);
  and (_15937_, _05764_, \oc8051_golden_model_1.ACC [2]);
  nor (_15938_, _15617_, _15937_);
  nor (_15939_, _10491_, _15938_);
  and (_15940_, _10491_, _15938_);
  nor (_15941_, _15940_, _15939_);
  and (_15942_, _15941_, \oc8051_golden_model_1.PSW [7]);
  nor (_15943_, _15941_, \oc8051_golden_model_1.PSW [7]);
  nor (_15944_, _15943_, _15942_);
  and (_15945_, _15944_, _15936_);
  nor (_15946_, _15944_, _15936_);
  or (_15947_, _15946_, _15945_);
  nand (_15948_, _15947_, _03883_);
  and (_15949_, _15948_, _08321_);
  and (_15950_, _15949_, _15934_);
  and (_15951_, _04139_, \oc8051_golden_model_1.ACC [2]);
  nor (_15952_, _15629_, _15951_);
  nor (_15953_, _10509_, _15952_);
  and (_15954_, _10509_, _15952_);
  nor (_15955_, _15954_, _15953_);
  and (_15956_, _15955_, \oc8051_golden_model_1.PSW [7]);
  nor (_15957_, _15955_, \oc8051_golden_model_1.PSW [7]);
  nor (_15958_, _15957_, _15956_);
  and (_15959_, _15958_, _15634_);
  nor (_15960_, _15958_, _15634_);
  or (_15961_, _15960_, _15959_);
  nor (_15962_, _15961_, _08321_);
  or (_15963_, _15962_, _03425_);
  or (_15964_, _15963_, _15950_);
  nand (_15965_, _03678_, _03425_);
  and (_15966_, _15965_, _03747_);
  and (_15967_, _15966_, _15964_);
  nor (_15968_, _12668_, _08465_);
  nor (_15969_, _15968_, _15855_);
  nor (_15970_, _15969_, _03747_);
  or (_15971_, _15970_, _07927_);
  or (_15972_, _15971_, _15967_);
  and (_15973_, _06964_, _05429_);
  nor (_15974_, _15973_, _15830_);
  nand (_15975_, _15974_, _03737_);
  nand (_15976_, _15892_, _08474_);
  and (_15977_, _15976_, _03820_);
  and (_15978_, _15977_, _15975_);
  and (_15979_, _15978_, _15972_);
  nor (_15980_, _12775_, _08479_);
  nor (_15981_, _15980_, _15830_);
  nor (_15982_, _15981_, _03820_);
  or (_15983_, _15982_, _07010_);
  or (_15984_, _15983_, _15979_);
  or (_15985_, _07151_, _07011_);
  and (_15986_, _15985_, _03479_);
  and (_15987_, _15986_, _15984_);
  nor (_15988_, _03678_, _03479_);
  or (_15989_, _15988_, _03903_);
  or (_15990_, _15989_, _15987_);
  and (_15991_, _05429_, _06345_);
  nor (_15992_, _15991_, _15830_);
  nand (_15993_, _15992_, _03903_);
  and (_15994_, _15993_, _08493_);
  and (_15995_, _15994_, _15990_);
  or (_15996_, _15995_, _15838_);
  and (_15997_, _08508_, _08502_);
  nor (_15998_, _15678_, _04397_);
  and (_15999_, _15998_, _15997_);
  and (_16000_, _15999_, _15996_);
  not (_16001_, _15999_);
  and (_16002_, _16001_, _15825_);
  or (_16003_, _16002_, _16000_);
  and (_16004_, _16003_, _08520_);
  and (_16005_, _15841_, _08519_);
  or (_16006_, _16005_, _04016_);
  or (_16007_, _16006_, _16004_);
  or (_16008_, _10491_, _04017_);
  and (_16009_, _16008_, _08531_);
  and (_16010_, _16009_, _16007_);
  and (_16011_, _08530_, _10509_);
  or (_16012_, _16011_, _03897_);
  or (_16013_, _16012_, _16010_);
  and (_16014_, _16013_, _15837_);
  or (_16015_, _16014_, _04018_);
  or (_16016_, _15830_, _04792_);
  and (_16017_, _16016_, _04186_);
  and (_16018_, _16017_, _16015_);
  nand (_16019_, _03729_, _03387_);
  not (_16020_, _04186_);
  nand (_16021_, _08013_, _16020_);
  nand (_16022_, _16021_, _16019_);
  or (_16023_, _16022_, _16018_);
  and (_16024_, _03719_, _03387_);
  not (_16025_, _16024_);
  or (_16026_, _08013_, _16019_);
  and (_16027_, _16026_, _16025_);
  and (_16028_, _16027_, _16023_);
  and (_16029_, _16024_, _08013_);
  or (_16030_, _16029_, _08547_);
  or (_16031_, _16030_, _16028_);
  or (_16032_, _08548_, _08705_);
  and (_16033_, _16032_, _16031_);
  or (_16034_, _16033_, _04025_);
  or (_16035_, _08744_, _04026_);
  and (_16036_, _16035_, _08557_);
  and (_16037_, _16036_, _16034_);
  and (_16038_, _08553_, _08784_);
  or (_16039_, _16038_, _16037_);
  and (_16040_, _16039_, _03909_);
  or (_16041_, _15992_, _08742_);
  nor (_16042_, _16041_, _03909_);
  or (_16043_, _16042_, _08563_);
  or (_16044_, _16043_, _16040_);
  nand (_16045_, _08563_, _08014_);
  and (_16046_, _16045_, _08567_);
  and (_16047_, _16046_, _16044_);
  and (_16048_, _08569_, _08014_);
  nor (_16049_, _16048_, _08570_);
  or (_16050_, _16049_, _16047_);
  and (_16051_, _16050_, _15834_);
  or (_16052_, _16051_, _08573_);
  nand (_16053_, _08573_, _08706_);
  and (_16054_, _16053_, _04014_);
  and (_16055_, _16054_, _16052_);
  nand (_16056_, _08583_, _08742_);
  and (_16057_, _16056_, _08582_);
  or (_16058_, _16057_, _16055_);
  nand (_16059_, _08580_, _08785_);
  and (_16060_, _16059_, _06567_);
  and (_16061_, _16060_, _16058_);
  or (_16062_, _16061_, _15833_);
  and (_16063_, _16062_, _08119_);
  and (_16064_, _08100_, _08079_);
  nor (_16065_, _16064_, _08101_);
  and (_16066_, _16065_, _08590_);
  or (_16067_, _16066_, _08597_);
  or (_16068_, _16067_, _16063_);
  and (_16069_, _08612_, _08285_);
  nor (_16070_, _16069_, _08613_);
  or (_16071_, _16070_, _08599_);
  and (_16072_, _16071_, _04023_);
  and (_16073_, _16072_, _16068_);
  and (_16074_, _08642_, _08358_);
  nor (_16075_, _16074_, _08643_);
  and (_16076_, _16075_, _04022_);
  or (_16077_, _16076_, _08627_);
  or (_16078_, _16077_, _16073_);
  and (_16079_, _08672_, _08428_);
  nor (_16080_, _16079_, _08673_);
  or (_16081_, _16080_, _08659_);
  and (_16082_, _16081_, _08658_);
  and (_16083_, _16082_, _16078_);
  nand (_16084_, _08657_, \oc8051_golden_model_1.ACC [2]);
  nand (_16085_, _16084_, _07999_);
  or (_16087_, _16085_, _16083_);
  and (_16088_, _16087_, _15829_);
  or (_16089_, _16088_, _08691_);
  nor (_16090_, _08718_, _15841_);
  and (_16091_, _08718_, _15841_);
  nor (_16092_, _16091_, _16090_);
  nand (_16093_, _16092_, _08691_);
  and (_16094_, _16093_, _04140_);
  and (_16095_, _16094_, _16089_);
  nor (_16096_, _08757_, _10491_);
  and (_16098_, _08757_, _10491_);
  nor (_16099_, _16098_, _16096_);
  nand (_16100_, _16099_, _15201_);
  and (_16101_, _16100_, _10057_);
  or (_16102_, _16101_, _16095_);
  nor (_16103_, _08797_, _10509_);
  and (_16104_, _08797_, _10509_);
  nor (_16105_, _16104_, _16103_);
  nand (_16106_, _16105_, _08733_);
  and (_16107_, _16106_, _08773_);
  and (_16109_, _16107_, _16102_);
  and (_16110_, _08772_, \oc8051_golden_model_1.ACC [2]);
  or (_16111_, _16110_, _03773_);
  or (_16112_, _16111_, _16109_);
  nand (_16113_, _15876_, _03773_);
  and (_16114_, _16113_, _08816_);
  and (_16115_, _16114_, _16112_);
  nor (_16116_, _15797_, _07184_);
  or (_16117_, _16116_, _08822_);
  and (_16118_, _16117_, _08815_);
  or (_16120_, _16118_, _08820_);
  or (_16121_, _16120_, _16115_);
  nand (_16122_, _08820_, _07090_);
  and (_16123_, _16122_, _03375_);
  and (_16124_, _16123_, _16121_);
  nor (_16125_, _15908_, _03375_);
  or (_16126_, _16125_, _03772_);
  or (_16127_, _16126_, _16124_);
  and (_16128_, _12848_, _05429_);
  nor (_16129_, _16128_, _15830_);
  nand (_16131_, _16129_, _03772_);
  and (_16132_, _16131_, _08838_);
  and (_16133_, _16132_, _16127_);
  or (_16134_, _15814_, \oc8051_golden_model_1.ACC [3]);
  and (_16135_, _16134_, _08846_);
  and (_16136_, _16135_, _08837_);
  or (_16137_, _16136_, _08844_);
  or (_16138_, _16137_, _16133_);
  nand (_16139_, _08844_, _07090_);
  and (_16140_, _16139_, _43152_);
  and (_16142_, _16140_, _16138_);
  or (_16143_, _16142_, _15824_);
  and (_43386_, _16143_, _41894_);
  nor (_16144_, _43152_, _07090_);
  nand (_16145_, _08772_, _07184_);
  nor (_16146_, _08614_, _08277_);
  nor (_16147_, _16146_, _08615_);
  or (_16148_, _16147_, _08599_);
  nand (_16149_, _08580_, _08782_);
  nor (_16150_, _05429_, _07090_);
  and (_16152_, _12997_, _05429_);
  nor (_16153_, _16152_, _16150_);
  nand (_16154_, _16153_, _03897_);
  or (_16155_, _08704_, _08520_);
  or (_16156_, _08502_, _08012_);
  or (_16157_, _08157_, _05950_);
  or (_16158_, _10400_, _05950_);
  nor (_16159_, _04263_, _07090_);
  and (_16160_, _04263_, _07090_);
  or (_16161_, _16160_, _16159_);
  or (_16163_, _16161_, _08169_);
  and (_16164_, _16163_, _08160_);
  and (_16165_, _16164_, _16158_);
  and (_16166_, _08159_, _06969_);
  or (_16167_, _16166_, _16165_);
  and (_16168_, _16167_, _08163_);
  nor (_16169_, _12891_, _08479_);
  nor (_16170_, _16169_, _16150_);
  nor (_16171_, _16170_, _04722_);
  or (_16172_, _16171_, _08179_);
  or (_16174_, _16172_, _16168_);
  nor (_16175_, _08186_, \oc8051_golden_model_1.ACC [4]);
  or (_16176_, _16175_, _08192_);
  nand (_16177_, _16176_, _08179_);
  and (_16178_, _16177_, _03856_);
  and (_16179_, _16178_, _16174_);
  nor (_16180_, _06096_, _07090_);
  and (_16181_, _12875_, _06096_);
  nor (_16182_, _16181_, _16180_);
  nor (_16183_, _16182_, _03764_);
  and (_16185_, _05950_, _05429_);
  nor (_16186_, _16185_, _16150_);
  nor (_16187_, _16186_, _04733_);
  or (_16188_, _16187_, _08212_);
  or (_16189_, _16188_, _16183_);
  or (_16190_, _16189_, _16179_);
  and (_16191_, _16190_, _16157_);
  or (_16192_, _16191_, _04738_);
  or (_16193_, _06969_, _04739_);
  and (_16194_, _16193_, _03855_);
  and (_16196_, _16194_, _16192_);
  nor (_16197_, _05953_, _03855_);
  or (_16198_, _16197_, _08224_);
  or (_16199_, _16198_, _16196_);
  nand (_16200_, _08224_, _03498_);
  and (_16201_, _16200_, _16199_);
  or (_16202_, _16201_, _03759_);
  and (_16203_, _12870_, _06096_);
  nor (_16204_, _16203_, _16180_);
  nand (_16205_, _16204_, _03759_);
  and (_16207_, _16205_, _03753_);
  and (_16208_, _16207_, _16202_);
  and (_16209_, _16181_, _12874_);
  nor (_16210_, _16209_, _16180_);
  nor (_16211_, _16210_, _03753_);
  or (_16212_, _16211_, _07399_);
  or (_16213_, _16212_, _16208_);
  nor (_16214_, _07864_, _07862_);
  nor (_16215_, _16214_, _07865_);
  or (_16216_, _16215_, _07405_);
  and (_16218_, _16216_, _16213_);
  or (_16219_, _16218_, _15513_);
  or (_16220_, _15924_, _15921_);
  and (_16221_, _05119_, _07184_);
  or (_16222_, _05119_, _07184_);
  and (_16223_, _15917_, _16222_);
  or (_16224_, _16223_, _16221_);
  nor (_16225_, _16224_, _08012_);
  and (_16226_, _16224_, _08012_);
  nor (_16227_, _16226_, _16225_);
  and (_16229_, _16227_, \oc8051_golden_model_1.PSW [7]);
  nor (_16230_, _16227_, \oc8051_golden_model_1.PSW [7]);
  nor (_16231_, _16230_, _16229_);
  and (_16232_, _16231_, _16220_);
  nor (_16233_, _16231_, _16220_);
  nor (_16234_, _16233_, _16232_);
  or (_16235_, _16234_, _08153_);
  and (_16236_, _16235_, _16219_);
  or (_16237_, _16236_, _04330_);
  or (_16238_, _15848_, _15845_);
  and (_16240_, _06964_, _07184_);
  or (_16241_, _06964_, _07184_);
  and (_16242_, _16241_, _15840_);
  or (_16243_, _16242_, _16240_);
  nor (_16244_, _08704_, _16243_);
  and (_16245_, _08704_, _16243_);
  nor (_16246_, _16245_, _16244_);
  and (_16247_, _16246_, \oc8051_golden_model_1.PSW [7]);
  nor (_16248_, _16246_, \oc8051_golden_model_1.PSW [7]);
  nor (_16249_, _16248_, _16247_);
  and (_16251_, _16249_, _16238_);
  nor (_16252_, _16249_, _16238_);
  nor (_16253_, _16252_, _16251_);
  or (_16254_, _16253_, _08248_);
  and (_16255_, _16254_, _16237_);
  or (_16256_, _16255_, _03883_);
  or (_16257_, _15945_, _15942_);
  or (_16258_, _15938_, _11820_);
  and (_16259_, _16258_, _11819_);
  nor (_16260_, _08741_, _16259_);
  and (_16261_, _08741_, _16259_);
  nor (_16262_, _16261_, _16260_);
  and (_16263_, _16262_, \oc8051_golden_model_1.PSW [7]);
  nor (_16264_, _16262_, \oc8051_golden_model_1.PSW [7]);
  nor (_16265_, _16264_, _16263_);
  and (_16266_, _16265_, _16257_);
  nor (_16267_, _16265_, _16257_);
  nor (_16268_, _16267_, _16266_);
  or (_16269_, _16268_, _03888_);
  and (_16270_, _16269_, _08321_);
  and (_16272_, _16270_, _16256_);
  or (_16273_, _15959_, _15956_);
  or (_16274_, _15952_, _11850_);
  and (_16275_, _16274_, _11849_);
  nor (_16276_, _08783_, _16275_);
  and (_16277_, _08783_, _16275_);
  nor (_16278_, _16277_, _16276_);
  and (_16279_, _16278_, \oc8051_golden_model_1.PSW [7]);
  nor (_16280_, _16278_, \oc8051_golden_model_1.PSW [7]);
  nor (_16281_, _16280_, _16279_);
  and (_16283_, _16281_, _16273_);
  nor (_16284_, _16281_, _16273_);
  nor (_16285_, _16284_, _16283_);
  and (_16286_, _16285_, _08320_);
  or (_16287_, _16286_, _03425_);
  or (_16288_, _16287_, _16272_);
  nand (_16289_, _04526_, _03425_);
  and (_16290_, _16289_, _03747_);
  and (_16291_, _16290_, _16288_);
  nor (_16292_, _12872_, _08465_);
  nor (_16294_, _16292_, _16180_);
  nor (_16295_, _16294_, _03747_);
  or (_16296_, _16295_, _07927_);
  or (_16297_, _16296_, _16291_);
  and (_16298_, _06969_, _05429_);
  nor (_16299_, _16298_, _16150_);
  nand (_16300_, _16299_, _03737_);
  nand (_16301_, _16186_, _08474_);
  and (_16302_, _16301_, _03820_);
  and (_16303_, _16302_, _16300_);
  and (_16305_, _16303_, _16297_);
  nor (_16306_, _12982_, _08479_);
  nor (_16307_, _16306_, _16150_);
  nor (_16308_, _16307_, _03820_);
  or (_16309_, _16308_, _07010_);
  or (_16310_, _16309_, _16305_);
  or (_16311_, _07099_, _07011_);
  and (_16312_, _16311_, _03479_);
  and (_16313_, _16312_, _16310_);
  nor (_16314_, _04526_, _03479_);
  or (_16316_, _16314_, _03903_);
  or (_16317_, _16316_, _16313_);
  and (_16318_, _06456_, _05429_);
  nor (_16319_, _16318_, _16150_);
  nand (_16320_, _16319_, _03903_);
  and (_16321_, _16320_, _08493_);
  and (_16322_, _16321_, _16317_);
  nor (_16323_, _08493_, _04526_);
  or (_16324_, _16323_, _08503_);
  or (_16325_, _16324_, _16322_);
  and (_16327_, _16325_, _16156_);
  or (_16328_, _16327_, _04400_);
  not (_16329_, _04400_);
  or (_16330_, _08012_, _16329_);
  nor (_16331_, _08506_, _04394_);
  nand (_16332_, _16331_, _15679_);
  nor (_16333_, _16332_, _04397_);
  and (_16334_, _16333_, _16330_);
  and (_16335_, _16334_, _16328_);
  not (_16336_, _16333_);
  and (_16338_, _16336_, _08012_);
  or (_16339_, _16338_, _08519_);
  or (_16340_, _16339_, _16335_);
  and (_16341_, _16340_, _16155_);
  or (_16342_, _16341_, _04016_);
  or (_16343_, _08741_, _04017_);
  and (_16344_, _16343_, _08531_);
  and (_16345_, _16344_, _16342_);
  and (_16346_, _08530_, _08783_);
  or (_16347_, _16346_, _03897_);
  or (_16349_, _16347_, _16345_);
  and (_16350_, _16349_, _16154_);
  or (_16351_, _16350_, _04018_);
  or (_16352_, _16150_, _04792_);
  and (_16353_, _16352_, _04186_);
  and (_16354_, _16353_, _16351_);
  and (_16355_, _03728_, _03387_);
  or (_16356_, _16355_, _08010_);
  and (_16357_, _16356_, _08122_);
  or (_16358_, _16357_, _16354_);
  not (_16360_, _16355_);
  or (_16361_, _16360_, _08010_);
  and (_16362_, _16361_, _08548_);
  and (_16363_, _16362_, _16358_);
  and (_16364_, _08547_, _08702_);
  or (_16365_, _16364_, _16363_);
  and (_16366_, _16365_, _04026_);
  and (_16367_, _08739_, _04025_);
  or (_16368_, _16367_, _08553_);
  or (_16369_, _16368_, _16366_);
  or (_16371_, _08557_, _08781_);
  and (_16372_, _16371_, _03909_);
  and (_16373_, _16372_, _16369_);
  not (_16374_, _10071_);
  or (_16375_, _16319_, _08740_);
  nor (_16376_, _16375_, _03909_);
  or (_16377_, _16376_, _16374_);
  or (_16378_, _16377_, _16373_);
  nand (_16379_, _16374_, _08011_);
  and (_16380_, _16379_, _08569_);
  and (_16382_, _16380_, _16378_);
  nor (_16383_, _08569_, _08011_);
  or (_16384_, _16383_, _08573_);
  or (_16385_, _16384_, _16382_);
  nand (_16386_, _08573_, _08703_);
  and (_16387_, _16386_, _04014_);
  and (_16388_, _16387_, _16385_);
  nand (_16389_, _08583_, _08740_);
  and (_16390_, _16389_, _08582_);
  or (_16391_, _16390_, _16388_);
  and (_16393_, _16391_, _16149_);
  or (_16394_, _16393_, _03914_);
  nor (_16395_, _12996_, _08479_);
  nor (_16396_, _16395_, _16150_);
  nand (_16397_, _16396_, _03914_);
  and (_16398_, _16397_, _08119_);
  and (_16399_, _16398_, _16394_);
  nor (_16400_, _08102_, _08071_);
  nor (_16401_, _16400_, _08103_);
  and (_16402_, _16401_, _08590_);
  or (_16404_, _16402_, _08597_);
  or (_16405_, _16404_, _16399_);
  and (_16406_, _16405_, _16148_);
  or (_16407_, _16406_, _04022_);
  nor (_16408_, _08644_, _08351_);
  nor (_16409_, _16408_, _08645_);
  or (_16410_, _16409_, _04023_);
  and (_16411_, _16410_, _08659_);
  and (_16412_, _16411_, _16407_);
  nor (_16413_, _08674_, _08422_);
  nor (_16415_, _16413_, _08675_);
  and (_16416_, _16415_, _08627_);
  or (_16417_, _16416_, _08657_);
  or (_16418_, _16417_, _16412_);
  nand (_16419_, _08657_, _07184_);
  and (_16420_, _16419_, _07999_);
  and (_16421_, _16420_, _16418_);
  nor (_16422_, _08028_, _08012_);
  nor (_16423_, _16422_, _08029_);
  and (_16424_, _16423_, _15460_);
  or (_16426_, _16424_, _16421_);
  and (_16427_, _16426_, _10058_);
  nor (_16428_, _08720_, _08704_);
  nor (_16429_, _16428_, _08721_);
  and (_16430_, _16429_, _08691_);
  or (_16431_, _16430_, _03779_);
  or (_16432_, _16431_, _16427_);
  nor (_16433_, _08759_, _08741_);
  nor (_16434_, _16433_, _08760_);
  or (_16435_, _16434_, _04140_);
  and (_16437_, _16435_, _15201_);
  and (_16438_, _16437_, _16432_);
  nor (_16439_, _08799_, _08783_);
  nor (_16440_, _16439_, _08800_);
  and (_16441_, _16440_, _08733_);
  or (_16442_, _16441_, _08772_);
  or (_16443_, _16442_, _16438_);
  and (_16444_, _16443_, _16145_);
  or (_16445_, _16444_, _03773_);
  nand (_16446_, _16170_, _03773_);
  and (_16448_, _16446_, _08816_);
  and (_16449_, _16448_, _16445_);
  and (_16450_, _08822_, _07090_);
  nor (_16451_, _08822_, _07090_);
  nor (_16452_, _16451_, _16450_);
  not (_16453_, _16452_);
  nor (_16454_, _16453_, _08820_);
  nor (_16455_, _16454_, _10943_);
  or (_16456_, _16455_, _16449_);
  nand (_16457_, _08820_, _07084_);
  and (_16460_, _16457_, _03375_);
  and (_16461_, _16460_, _16456_);
  nor (_16462_, _16204_, _03375_);
  or (_16463_, _16462_, _03772_);
  or (_16464_, _16463_, _16461_);
  and (_16465_, _13056_, _05429_);
  nor (_16466_, _16465_, _16150_);
  nand (_16467_, _16466_, _03772_);
  and (_16468_, _16467_, _08838_);
  and (_16469_, _16468_, _16464_);
  and (_16471_, _08846_, _07090_);
  nor (_16472_, _16471_, _08847_);
  nor (_16473_, _16472_, _08844_);
  nor (_16474_, _16473_, _10965_);
  or (_16475_, _16474_, _16469_);
  nand (_16476_, _08844_, _07084_);
  and (_16477_, _16476_, _43152_);
  and (_16478_, _16477_, _16475_);
  or (_16479_, _16478_, _16144_);
  and (_43387_, _16479_, _41894_);
  nor (_16481_, _43152_, _07084_);
  and (_16482_, _08030_, _08009_);
  nor (_16483_, _16482_, _08031_);
  or (_16484_, _16483_, _07999_);
  and (_16485_, _08104_, _08062_);
  nor (_16486_, _16485_, _08105_);
  or (_16487_, _16486_, _08119_);
  nor (_16488_, _08569_, _08007_);
  or (_16489_, _16488_, _08573_);
  not (_16490_, _08006_);
  and (_16492_, _16019_, _04186_);
  nor (_16493_, _16492_, _16490_);
  nor (_16494_, _05429_, _07084_);
  and (_16495_, _13196_, _05429_);
  nor (_16496_, _16495_, _16494_);
  nand (_16497_, _16496_, _03897_);
  or (_16498_, _08700_, _08520_);
  nor (_16499_, _08493_, _04093_);
  and (_16500_, _06918_, \oc8051_golden_model_1.ACC [4]);
  nor (_16501_, _16244_, _16500_);
  nor (_16503_, _08700_, _16501_);
  and (_16504_, _08700_, _16501_);
  nor (_16505_, _16504_, _16503_);
  and (_16506_, _16505_, \oc8051_golden_model_1.PSW [7]);
  nor (_16507_, _16505_, \oc8051_golden_model_1.PSW [7]);
  nor (_16508_, _16507_, _16506_);
  nor (_16509_, _16251_, _16247_);
  not (_16510_, _16509_);
  and (_16511_, _16510_, _16508_);
  nor (_16512_, _16510_, _16508_);
  nor (_16514_, _16512_, _16511_);
  or (_16515_, _16514_, _08248_);
  nor (_16516_, _06096_, _07084_);
  and (_16517_, _13094_, _06096_);
  and (_16518_, _16517_, _13109_);
  nor (_16519_, _16518_, _16516_);
  nor (_16520_, _16519_, _03753_);
  or (_16521_, _08157_, _05857_);
  or (_16522_, _10400_, _05857_);
  nor (_16523_, _04263_, _07084_);
  and (_16525_, _04263_, _07084_);
  or (_16526_, _16525_, _16523_);
  or (_16527_, _16526_, _08169_);
  and (_16528_, _16527_, _08160_);
  and (_16529_, _16528_, _16522_);
  and (_16530_, _08159_, _06968_);
  or (_16531_, _16530_, _16529_);
  and (_16532_, _16531_, _08163_);
  nor (_16533_, _13090_, _08479_);
  nor (_16534_, _16533_, _16494_);
  nor (_16536_, _16534_, _04722_);
  or (_16537_, _16536_, _08179_);
  or (_16538_, _16537_, _16532_);
  and (_16539_, _11762_, _08194_);
  nor (_16540_, _11762_, _08194_);
  nor (_16541_, _16540_, _16539_);
  nand (_16542_, _16541_, _08179_);
  and (_16543_, _16542_, _03856_);
  and (_16544_, _16543_, _16538_);
  nor (_16545_, _16517_, _16516_);
  nor (_16547_, _16545_, _03764_);
  and (_16548_, _05857_, _05429_);
  nor (_16549_, _16548_, _16494_);
  nor (_16550_, _16549_, _04733_);
  or (_16551_, _16550_, _08212_);
  or (_16552_, _16551_, _16547_);
  or (_16553_, _16552_, _16544_);
  and (_16554_, _16553_, _16521_);
  or (_16555_, _16554_, _04738_);
  or (_16556_, _06968_, _04739_);
  and (_16558_, _16556_, _03855_);
  and (_16559_, _16558_, _16555_);
  nor (_16560_, _05859_, _03855_);
  or (_16561_, _16560_, _08224_);
  or (_16562_, _16561_, _16559_);
  nand (_16563_, _08224_, _03474_);
  and (_16564_, _16563_, _16562_);
  or (_16565_, _16564_, _03759_);
  and (_16566_, _13071_, _06096_);
  nor (_16567_, _16566_, _16516_);
  nand (_16569_, _16567_, _03759_);
  and (_16570_, _16569_, _03753_);
  and (_16571_, _16570_, _16565_);
  or (_16572_, _16571_, _16520_);
  and (_16573_, _16572_, _07405_);
  nor (_16574_, _07867_, _07865_);
  nor (_16575_, _16574_, _07868_);
  and (_16576_, _16575_, _07399_);
  or (_16577_, _16576_, _11880_);
  or (_16578_, _16577_, _16573_);
  nor (_16580_, _05950_, _07090_);
  nor (_16581_, _16225_, _16580_);
  nor (_16582_, _16581_, _08009_);
  and (_16583_, _16581_, _08009_);
  nor (_16584_, _16583_, _16582_);
  nor (_16585_, _16584_, _08297_);
  and (_16586_, _16584_, _08297_);
  nor (_16587_, _16586_, _16585_);
  nor (_16588_, _16232_, _16229_);
  not (_16589_, _16588_);
  and (_16591_, _16589_, _16587_);
  nor (_16592_, _16589_, _16587_);
  nor (_16593_, _16592_, _16591_);
  or (_16594_, _16593_, _11879_);
  and (_16595_, _16594_, _11883_);
  and (_16596_, _16595_, _16578_);
  and (_16597_, _16593_, _04335_);
  or (_16598_, _16597_, _04330_);
  or (_16599_, _16598_, _16596_);
  and (_16600_, _16599_, _16515_);
  or (_16602_, _16600_, _03883_);
  and (_16603_, _05953_, \oc8051_golden_model_1.ACC [4]);
  nor (_16604_, _16260_, _16603_);
  nor (_16605_, _10493_, _16604_);
  and (_16606_, _10493_, _16604_);
  nor (_16607_, _16606_, _16605_);
  and (_16608_, _16607_, \oc8051_golden_model_1.PSW [7]);
  nor (_16609_, _16607_, \oc8051_golden_model_1.PSW [7]);
  nor (_16610_, _16609_, _16608_);
  nor (_16611_, _16266_, _16263_);
  not (_16613_, _16611_);
  and (_16614_, _16613_, _16610_);
  nor (_16615_, _16613_, _16610_);
  nor (_16616_, _16615_, _16614_);
  or (_16617_, _16616_, _03888_);
  and (_16618_, _16617_, _08321_);
  and (_16619_, _16618_, _16602_);
  and (_16620_, _04526_, \oc8051_golden_model_1.ACC [4]);
  nor (_16621_, _16276_, _16620_);
  nor (_16622_, _08779_, _16621_);
  and (_16624_, _08779_, _16621_);
  nor (_16625_, _16624_, _16622_);
  and (_16626_, _16625_, \oc8051_golden_model_1.PSW [7]);
  nor (_16627_, _16625_, \oc8051_golden_model_1.PSW [7]);
  nor (_16628_, _16627_, _16626_);
  nor (_16629_, _16283_, _16279_);
  not (_16630_, _16629_);
  and (_16631_, _16630_, _16628_);
  nor (_16632_, _16630_, _16628_);
  nor (_16633_, _16632_, _16631_);
  and (_16635_, _16633_, _08320_);
  or (_16636_, _16635_, _03425_);
  or (_16637_, _16636_, _16619_);
  nand (_16638_, _04093_, _03425_);
  and (_16639_, _16638_, _03747_);
  and (_16640_, _16639_, _16637_);
  nor (_16641_, _13073_, _08465_);
  nor (_16642_, _16641_, _16516_);
  nor (_16643_, _16642_, _03747_);
  or (_16644_, _16643_, _07927_);
  or (_16646_, _16644_, _16640_);
  and (_16647_, _06968_, _05429_);
  nor (_16648_, _16647_, _16494_);
  nand (_16649_, _16648_, _03737_);
  nand (_16650_, _16549_, _08474_);
  and (_16651_, _16650_, _03820_);
  and (_16652_, _16651_, _16649_);
  and (_16653_, _16652_, _16646_);
  nor (_16654_, _13182_, _08479_);
  nor (_16655_, _16654_, _16494_);
  nor (_16657_, _16655_, _03820_);
  or (_16658_, _16657_, _07010_);
  or (_16659_, _16658_, _16653_);
  or (_16660_, _07069_, _07011_);
  and (_16661_, _16660_, _03479_);
  and (_16662_, _16661_, _16659_);
  nor (_16663_, _04093_, _03479_);
  or (_16664_, _16663_, _03903_);
  or (_16665_, _16664_, _16662_);
  and (_16666_, _06447_, _05429_);
  nor (_16668_, _16666_, _16494_);
  nand (_16669_, _16668_, _03903_);
  and (_16670_, _16669_, _08493_);
  and (_16671_, _16670_, _16665_);
  or (_16672_, _16671_, _16499_);
  and (_16673_, _16672_, _08502_);
  and (_16674_, _08503_, _08008_);
  or (_16675_, _16674_, _04400_);
  or (_16676_, _16675_, _16673_);
  nor (_16677_, _08008_, _16329_);
  nor (_16679_, _16677_, _08506_);
  and (_16680_, _16679_, _16676_);
  and (_16681_, _08008_, _08506_);
  or (_16682_, _16681_, _04394_);
  or (_16683_, _16682_, _16680_);
  or (_16684_, _08008_, _04395_);
  and (_16685_, _16684_, _15998_);
  and (_16686_, _16685_, _16683_);
  not (_16687_, _15998_);
  and (_16688_, _16687_, _08008_);
  or (_16690_, _16688_, _08519_);
  or (_16691_, _16690_, _16686_);
  and (_16692_, _16691_, _16498_);
  or (_16693_, _16692_, _04016_);
  or (_16694_, _10493_, _04017_);
  and (_16695_, _16694_, _08531_);
  and (_16696_, _16695_, _16693_);
  and (_16697_, _08530_, _08779_);
  or (_16698_, _16697_, _03897_);
  or (_16699_, _16698_, _16696_);
  and (_16701_, _16699_, _16497_);
  or (_16702_, _16701_, _04018_);
  or (_16703_, _16494_, _04792_);
  and (_16704_, _16703_, _16492_);
  and (_16705_, _16704_, _16702_);
  or (_16706_, _16705_, _16493_);
  and (_16707_, _16706_, _16025_);
  and (_16708_, _16024_, _08006_);
  or (_16709_, _16708_, _16707_);
  and (_16710_, _16709_, _08548_);
  and (_16712_, _08547_, _08698_);
  or (_16713_, _16712_, _04025_);
  or (_16714_, _16713_, _16710_);
  or (_16715_, _08737_, _04026_);
  and (_16716_, _16715_, _08557_);
  and (_16717_, _16716_, _16714_);
  and (_16718_, _08553_, _08777_);
  or (_16719_, _16718_, _16717_);
  and (_16720_, _16719_, _03909_);
  or (_16721_, _16668_, _08738_);
  nor (_16723_, _16721_, _03909_);
  or (_16724_, _16723_, _08563_);
  or (_16725_, _16724_, _16720_);
  nand (_16726_, _08563_, _08007_);
  and (_16727_, _16726_, _08567_);
  and (_16728_, _16727_, _16725_);
  nor (_16729_, _08007_, _08567_);
  or (_16730_, _16729_, _16728_);
  and (_16731_, _16730_, _08569_);
  or (_16732_, _16731_, _16489_);
  nand (_16734_, _08573_, _08699_);
  and (_16735_, _16734_, _04014_);
  and (_16736_, _16735_, _16732_);
  nand (_16737_, _08583_, _08738_);
  and (_16738_, _16737_, _08582_);
  or (_16739_, _16738_, _16736_);
  nand (_16740_, _08580_, _08778_);
  and (_16741_, _16740_, _06567_);
  and (_16742_, _16741_, _16739_);
  nor (_16743_, _13195_, _08479_);
  nor (_16745_, _16743_, _16494_);
  nor (_16746_, _16745_, _06567_);
  or (_16747_, _16746_, _08590_);
  or (_16748_, _16747_, _16742_);
  and (_16749_, _16748_, _16487_);
  or (_16750_, _16749_, _08597_);
  and (_16751_, _08616_, _08274_);
  nor (_16752_, _16751_, _08617_);
  or (_16753_, _16752_, _08599_);
  and (_16754_, _16753_, _04023_);
  and (_16756_, _16754_, _16750_);
  and (_16757_, _08646_, _08348_);
  nor (_16758_, _16757_, _08647_);
  and (_16759_, _16758_, _04022_);
  or (_16760_, _16759_, _08627_);
  or (_16761_, _16760_, _16756_);
  and (_16762_, _08676_, _08416_);
  nor (_16763_, _16762_, _08677_);
  or (_16764_, _16763_, _08659_);
  and (_16765_, _16764_, _08658_);
  and (_16767_, _16765_, _16761_);
  nand (_16768_, _08657_, \oc8051_golden_model_1.ACC [4]);
  nand (_16769_, _16768_, _07999_);
  or (_16770_, _16769_, _16767_);
  and (_16771_, _16770_, _16484_);
  or (_16772_, _16771_, _08691_);
  and (_16773_, _08722_, _08701_);
  nor (_16774_, _16773_, _08723_);
  or (_16775_, _16774_, _10058_);
  and (_16776_, _16775_, _04140_);
  and (_16778_, _16776_, _16772_);
  nor (_16779_, _08761_, _10493_);
  and (_16780_, _08761_, _10493_);
  or (_16781_, _16780_, _16779_);
  or (_16782_, _16781_, _08733_);
  and (_16783_, _16782_, _10057_);
  or (_16784_, _16783_, _16778_);
  and (_16785_, _08801_, _08780_);
  nor (_16786_, _16785_, _08802_);
  or (_16787_, _16786_, _15201_);
  and (_16789_, _16787_, _08773_);
  and (_16790_, _16789_, _16784_);
  and (_16791_, _08772_, \oc8051_golden_model_1.ACC [4]);
  or (_16792_, _16791_, _03773_);
  or (_16793_, _16792_, _16790_);
  nand (_16794_, _16534_, _03773_);
  and (_16795_, _16794_, _08816_);
  and (_16796_, _16795_, _16793_);
  nor (_16797_, _16450_, _07084_);
  or (_16798_, _16797_, _08823_);
  and (_16800_, _16798_, _08815_);
  or (_16801_, _16800_, _08820_);
  or (_16802_, _16801_, _16796_);
  nand (_16803_, _08820_, _07036_);
  and (_16804_, _16803_, _03375_);
  and (_16805_, _16804_, _16802_);
  nor (_16806_, _16567_, _03375_);
  or (_16807_, _16806_, _03772_);
  or (_16808_, _16807_, _16805_);
  and (_16809_, _13255_, _05429_);
  nor (_16811_, _16809_, _16494_);
  nand (_16812_, _16811_, _03772_);
  and (_16813_, _16812_, _08838_);
  and (_16814_, _16813_, _16808_);
  nor (_16815_, _08847_, \oc8051_golden_model_1.ACC [5]);
  nor (_16816_, _16815_, _08848_);
  and (_16817_, _16816_, _08837_);
  or (_16818_, _16817_, _08844_);
  or (_16819_, _16818_, _16814_);
  nand (_16820_, _08844_, _07036_);
  and (_16822_, _16820_, _43152_);
  and (_16823_, _16822_, _16819_);
  or (_16824_, _16823_, _16481_);
  and (_43390_, _16824_, _41894_);
  nor (_16825_, _43152_, _07036_);
  nand (_16826_, _08772_, _07084_);
  nor (_16827_, _08618_, _08311_);
  nor (_16828_, _16827_, _08619_);
  or (_16829_, _16828_, _08599_);
  nand (_16830_, _08573_, _08696_);
  nor (_16832_, _08004_, _15158_);
  or (_16833_, _16832_, _15420_);
  nor (_16834_, _05429_, _07036_);
  and (_16835_, _13394_, _05429_);
  nor (_16836_, _16835_, _16834_);
  or (_16837_, _16836_, _08735_);
  nor (_16838_, _16837_, _03909_);
  and (_16839_, _13402_, _05429_);
  nor (_16840_, _16839_, _16834_);
  nand (_16841_, _16840_, _03897_);
  and (_16843_, _04760_, _03404_);
  and (_16844_, _16843_, _08697_);
  not (_16845_, _16843_);
  not (_16846_, _08005_);
  nor (_16847_, _04396_, _04204_);
  and (_16848_, _16847_, _16331_);
  nor (_16849_, _16848_, _16846_);
  or (_16850_, _06968_, _07084_);
  and (_16851_, _06968_, _07084_);
  or (_16852_, _16501_, _16851_);
  and (_16854_, _16852_, _16850_);
  nor (_16855_, _16854_, _08697_);
  and (_16856_, _16854_, _08697_);
  nor (_16857_, _16856_, _16855_);
  nor (_16858_, _16511_, _16506_);
  and (_16859_, _16858_, \oc8051_golden_model_1.PSW [7]);
  nor (_16860_, _16859_, _16857_);
  and (_16861_, _16859_, _16857_);
  nor (_16862_, _16861_, _16860_);
  and (_16863_, _16862_, _04330_);
  or (_16865_, _08157_, _06065_);
  or (_16866_, _10400_, _06065_);
  nor (_16867_, _04263_, _07036_);
  and (_16868_, _04263_, _07036_);
  or (_16869_, _16868_, _16867_);
  or (_16870_, _16869_, _08169_);
  and (_16871_, _16870_, _08160_);
  and (_16872_, _16871_, _16866_);
  and (_16873_, _08159_, _06641_);
  or (_16874_, _16873_, _16872_);
  and (_16876_, _16874_, _08163_);
  nor (_16877_, _13293_, _08479_);
  nor (_16878_, _16877_, _16834_);
  nor (_16879_, _16878_, _04722_);
  or (_16880_, _16879_, _08179_);
  or (_16881_, _16880_, _16876_);
  not (_16882_, _08196_);
  nor (_16883_, _16540_, _16882_);
  and (_16884_, _11761_, _08197_);
  nor (_16885_, _16884_, _16883_);
  nand (_16887_, _16885_, _08179_);
  and (_16888_, _16887_, _03856_);
  and (_16889_, _16888_, _16881_);
  nor (_16890_, _06096_, _07036_);
  and (_16891_, _13297_, _06096_);
  nor (_16892_, _16891_, _16890_);
  nor (_16893_, _16892_, _03764_);
  and (_16894_, _06065_, _05429_);
  nor (_16895_, _16894_, _16834_);
  nor (_16896_, _16895_, _04733_);
  or (_16898_, _16896_, _08212_);
  or (_16899_, _16898_, _16893_);
  or (_16900_, _16899_, _16889_);
  and (_16901_, _16900_, _16865_);
  or (_16902_, _16901_, _04738_);
  or (_16903_, _06641_, _04739_);
  and (_16904_, _16903_, _03855_);
  and (_16905_, _16904_, _16902_);
  nor (_16906_, _06068_, _03855_);
  or (_16907_, _16906_, _08224_);
  or (_16909_, _16907_, _16905_);
  nand (_16910_, _08224_, _07190_);
  and (_16911_, _16910_, _16909_);
  or (_16912_, _16911_, _03759_);
  and (_16913_, _13277_, _06096_);
  nor (_16914_, _16913_, _16890_);
  nand (_16915_, _16914_, _03759_);
  and (_16916_, _16915_, _03753_);
  and (_16917_, _16916_, _16912_);
  and (_16918_, _16891_, _13312_);
  nor (_16920_, _16918_, _16890_);
  nor (_16921_, _16920_, _03753_);
  or (_16922_, _16921_, _07399_);
  or (_16923_, _16922_, _16917_);
  nor (_16924_, _07870_, _07868_);
  nor (_16925_, _16924_, _07871_);
  or (_16926_, _16925_, _07405_);
  and (_16927_, _16926_, _16923_);
  or (_16928_, _16927_, _15513_);
  or (_16929_, _05857_, _07084_);
  and (_16931_, _05857_, _07084_);
  or (_16932_, _16581_, _16931_);
  and (_16933_, _16932_, _16929_);
  nor (_16934_, _16933_, _08005_);
  and (_16935_, _16933_, _08005_);
  nor (_16936_, _16935_, _16934_);
  nor (_16937_, _16591_, _16585_);
  and (_16938_, _16937_, \oc8051_golden_model_1.PSW [7]);
  nor (_16939_, _16938_, _16936_);
  and (_16940_, _16938_, _16936_);
  nor (_16942_, _16940_, _16939_);
  or (_16943_, _16942_, _08153_);
  and (_16944_, _16943_, _08248_);
  and (_16945_, _16944_, _16928_);
  or (_16946_, _16945_, _03883_);
  or (_16947_, _16946_, _16863_);
  or (_16948_, _16604_, _11813_);
  and (_16949_, _16948_, _11812_);
  nor (_16950_, _08736_, _16949_);
  and (_16951_, _08736_, _16949_);
  nor (_16953_, _16951_, _16950_);
  nor (_16954_, _16614_, _16608_);
  and (_16955_, _16954_, \oc8051_golden_model_1.PSW [7]);
  or (_16956_, _16955_, _16953_);
  nand (_16957_, _16955_, _16953_);
  and (_16958_, _16957_, _16956_);
  or (_16959_, _16958_, _03888_);
  and (_16960_, _16959_, _08321_);
  and (_16961_, _16960_, _16947_);
  or (_16962_, _16621_, _11837_);
  and (_16964_, _16962_, _11836_);
  nor (_16965_, _16964_, _08776_);
  and (_16966_, _16964_, _08776_);
  nor (_16967_, _16966_, _16965_);
  nor (_16968_, _16631_, _16626_);
  and (_16969_, _16968_, \oc8051_golden_model_1.PSW [7]);
  or (_16970_, _16969_, _16967_);
  nand (_16971_, _16969_, _16967_);
  and (_16972_, _16971_, _16970_);
  and (_16973_, _16972_, _08320_);
  or (_16975_, _16973_, _03425_);
  or (_16976_, _16975_, _16961_);
  nand (_16977_, _03810_, _03425_);
  and (_16978_, _16977_, _03747_);
  and (_16979_, _16978_, _16976_);
  nor (_16980_, _13279_, _08465_);
  nor (_16981_, _16980_, _16890_);
  nor (_16982_, _16981_, _03747_);
  or (_16983_, _16982_, _07927_);
  or (_16984_, _16983_, _16979_);
  and (_16986_, _06641_, _05429_);
  nor (_16987_, _16986_, _16834_);
  nand (_16988_, _16987_, _03737_);
  nand (_16989_, _16895_, _08474_);
  and (_16990_, _16989_, _03820_);
  and (_16991_, _16990_, _16988_);
  and (_16992_, _16991_, _16984_);
  nor (_16993_, _13387_, _08479_);
  nor (_16994_, _16993_, _16834_);
  nor (_16995_, _16994_, _03820_);
  or (_16997_, _16995_, _07010_);
  or (_16998_, _16997_, _16992_);
  not (_16999_, _07037_);
  and (_17000_, _07041_, _16999_);
  or (_17001_, _17000_, _07011_);
  and (_17002_, _17001_, _03479_);
  and (_17003_, _17002_, _16998_);
  nor (_17004_, _03810_, _03479_);
  or (_17005_, _17004_, _03903_);
  or (_17006_, _17005_, _17003_);
  nand (_17008_, _16836_, _03903_);
  and (_17009_, _17008_, _08493_);
  and (_17010_, _17009_, _17006_);
  and (_17011_, _03910_, _03404_);
  nor (_17012_, _08493_, _03810_);
  or (_17013_, _17012_, _17011_);
  or (_17014_, _17013_, _17010_);
  nand (_17015_, _16846_, _17011_);
  and (_17016_, _17015_, _16848_);
  and (_17017_, _17016_, _17014_);
  or (_17019_, _17017_, _16849_);
  and (_17020_, _17019_, _15998_);
  and (_17021_, _16687_, _08005_);
  or (_17022_, _17021_, _17020_);
  and (_17023_, _17022_, _16845_);
  nor (_17024_, _17023_, _16844_);
  nor (_17025_, _17024_, _04401_);
  and (_17026_, _08697_, _04401_);
  or (_17027_, _17026_, _04016_);
  or (_17028_, _17027_, _17025_);
  or (_17030_, _08736_, _04017_);
  and (_17031_, _17030_, _08531_);
  and (_17032_, _17031_, _17028_);
  and (_17033_, _08530_, _08776_);
  or (_17034_, _17033_, _03897_);
  or (_17035_, _17034_, _17032_);
  and (_17036_, _17035_, _16841_);
  or (_17037_, _17036_, _04018_);
  or (_17038_, _16834_, _04792_);
  and (_17039_, _17038_, _08121_);
  and (_17041_, _17039_, _17037_);
  and (_17042_, _08122_, _08003_);
  or (_17043_, _17042_, _08547_);
  or (_17044_, _17043_, _17041_);
  or (_17045_, _08548_, _08695_);
  and (_17046_, _17045_, _04026_);
  and (_17047_, _17046_, _17044_);
  or (_17048_, _08553_, _08734_);
  and (_17049_, _17048_, _10659_);
  or (_17050_, _17049_, _17047_);
  or (_17052_, _08557_, _08774_);
  and (_17053_, _17052_, _03909_);
  and (_17054_, _17053_, _17050_);
  nor (_17055_, _17054_, _16838_);
  nor (_17056_, _17055_, _15010_);
  not (_17057_, _15010_);
  nor (_17058_, _17057_, _08004_);
  or (_17059_, _17058_, _15008_);
  or (_17060_, _17059_, _17056_);
  and (_17061_, _17060_, _16833_);
  nor (_17063_, _08004_, _15159_);
  or (_17064_, _17063_, _08573_);
  or (_17065_, _17064_, _17061_);
  and (_17066_, _17065_, _16830_);
  or (_17067_, _17066_, _04013_);
  nand (_17068_, _08735_, _04013_);
  and (_17069_, _17068_, _08583_);
  and (_17070_, _17069_, _17067_);
  nor (_17071_, _08583_, _08775_);
  or (_17072_, _17071_, _03914_);
  or (_17074_, _17072_, _17070_);
  nor (_17075_, _13401_, _08479_);
  nor (_17076_, _17075_, _16834_);
  nand (_17077_, _17076_, _03914_);
  and (_17078_, _17077_, _08119_);
  and (_17079_, _17078_, _17074_);
  nor (_17080_, _08106_, _08054_);
  nor (_17081_, _17080_, _08107_);
  and (_17082_, _17081_, _08590_);
  or (_17083_, _17082_, _08597_);
  or (_17085_, _17083_, _17079_);
  and (_17086_, _17085_, _16829_);
  or (_17087_, _17086_, _04022_);
  nor (_17088_, _08648_, _08385_);
  nor (_17089_, _17088_, _08649_);
  or (_17090_, _17089_, _04023_);
  and (_17091_, _17090_, _08659_);
  and (_17092_, _17091_, _17087_);
  and (_17093_, _08678_, _08411_);
  nor (_17094_, _17093_, _08679_);
  and (_17096_, _17094_, _08627_);
  or (_17097_, _17096_, _08657_);
  or (_17098_, _17097_, _17092_);
  nand (_17099_, _08657_, _07084_);
  and (_17100_, _17099_, _07999_);
  and (_17101_, _17100_, _17098_);
  nor (_17102_, _08032_, _08005_);
  nor (_17103_, _17102_, _08033_);
  and (_17104_, _17103_, _15460_);
  or (_17105_, _17104_, _17101_);
  and (_17107_, _17105_, _10058_);
  nor (_17108_, _08724_, _08697_);
  nor (_17109_, _17108_, _08725_);
  and (_17110_, _17109_, _08691_);
  or (_17111_, _17110_, _03779_);
  or (_17112_, _17111_, _17107_);
  nor (_17113_, _08763_, _08736_);
  nor (_17114_, _17113_, _08764_);
  or (_17115_, _17114_, _04140_);
  and (_17116_, _17115_, _15201_);
  and (_17118_, _17116_, _17112_);
  nor (_17119_, _08803_, _08776_);
  nor (_17120_, _17119_, _08804_);
  and (_17121_, _17120_, _08733_);
  or (_17122_, _17121_, _08772_);
  or (_17123_, _17122_, _17118_);
  and (_17124_, _17123_, _16826_);
  or (_17125_, _17124_, _03773_);
  nand (_17126_, _16878_, _03773_);
  and (_17127_, _17126_, _08816_);
  and (_17129_, _17127_, _17125_);
  nor (_17130_, _08823_, _07036_);
  or (_17131_, _17130_, _08824_);
  and (_17132_, _17131_, _08815_);
  or (_17133_, _17132_, _08820_);
  or (_17134_, _17133_, _17129_);
  nand (_17135_, _08820_, _06554_);
  and (_17136_, _17135_, _03375_);
  and (_17137_, _17136_, _17134_);
  nor (_17138_, _16914_, _03375_);
  or (_17140_, _17138_, _03772_);
  or (_17141_, _17140_, _17137_);
  nor (_17142_, _13460_, _08479_);
  nor (_17143_, _17142_, _16834_);
  nand (_17144_, _17143_, _03772_);
  and (_17145_, _17144_, _08838_);
  and (_17146_, _17145_, _17141_);
  nor (_17147_, _08848_, \oc8051_golden_model_1.ACC [6]);
  nor (_17148_, _17147_, _08849_);
  and (_17149_, _17148_, _08837_);
  or (_17151_, _17149_, _08844_);
  or (_17152_, _17151_, _17146_);
  nand (_17153_, _08844_, _06554_);
  and (_17154_, _17153_, _43152_);
  and (_17155_, _17154_, _17152_);
  or (_17156_, _17155_, _16825_);
  and (_43391_, _17156_, _41894_);
  not (_17157_, _04144_);
  not (_17158_, \oc8051_golden_model_1.SBUF [0]);
  nor (_17159_, _05491_, _17158_);
  and (_17161_, _05716_, _05491_);
  nor (_17162_, _17161_, _17159_);
  and (_17163_, _17162_, _17157_);
  nand (_17164_, _08753_, _05491_);
  nor (_17165_, _17159_, _04785_);
  and (_17166_, _17165_, _17164_);
  and (_17167_, _06962_, _05491_);
  nor (_17168_, _17159_, _03738_);
  not (_17169_, _17168_);
  nor (_17170_, _17169_, _17167_);
  and (_17171_, _05491_, _04700_);
  nor (_17172_, _17171_, _17159_);
  and (_17173_, _17172_, _08474_);
  and (_17174_, _05491_, \oc8051_golden_model_1.ACC [0]);
  nor (_17175_, _17174_, _17159_);
  nor (_17176_, _17175_, _04708_);
  nor (_17177_, _04707_, _17158_);
  or (_17178_, _17177_, _17176_);
  and (_17179_, _17178_, _04722_);
  nor (_17180_, _17162_, _04722_);
  or (_17183_, _17180_, _17179_);
  and (_17184_, _17183_, _04733_);
  nor (_17185_, _17172_, _04733_);
  nor (_17186_, _17185_, _17184_);
  nor (_17187_, _17186_, _03854_);
  nor (_17188_, _17175_, _03855_);
  or (_17189_, _17188_, _07927_);
  nor (_17190_, _17189_, _17187_);
  nor (_17191_, _17190_, _17173_);
  not (_17192_, _17191_);
  nor (_17193_, _17192_, _17170_);
  and (_17194_, _17193_, _03820_);
  nor (_17195_, _12164_, _08897_);
  nor (_17196_, _17195_, _17159_);
  nor (_17197_, _17196_, _03820_);
  or (_17198_, _17197_, _17194_);
  and (_17199_, _17198_, _04778_);
  and (_17200_, _05491_, _06479_);
  nor (_17201_, _17200_, _17159_);
  nor (_17202_, _17201_, _04778_);
  or (_17205_, _17202_, _17199_);
  and (_17206_, _17205_, _04790_);
  and (_17207_, _12178_, _05491_);
  nor (_17208_, _17207_, _17159_);
  nor (_17209_, _17208_, _04790_);
  or (_17210_, _17209_, _17206_);
  and (_17211_, _17210_, _04792_);
  nor (_17212_, _10488_, _08897_);
  nor (_17213_, _17212_, _17159_);
  nand (_17214_, _17164_, _04018_);
  nor (_17216_, _17214_, _17213_);
  nor (_17217_, _17216_, _17211_);
  nor (_17218_, _17217_, _03908_);
  nor (_17219_, _17201_, _03909_);
  not (_17220_, _17219_);
  nor (_17221_, _17220_, _17161_);
  nor (_17222_, _17221_, _04027_);
  not (_17223_, _17222_);
  nor (_17224_, _17223_, _17218_);
  nor (_17225_, _17224_, _17166_);
  and (_17227_, _17225_, _06567_);
  nor (_17228_, _12177_, _08897_);
  nor (_17229_, _17228_, _17159_);
  nor (_17230_, _17229_, _06567_);
  or (_17231_, _17230_, _17227_);
  and (_17232_, _17231_, _06572_);
  nor (_17233_, _17213_, _06572_);
  nor (_17234_, _17233_, _17157_);
  not (_17235_, _17234_);
  nor (_17236_, _17235_, _17232_);
  nor (_17238_, _17236_, _17163_);
  or (_17239_, _17238_, _43156_);
  or (_17240_, _43152_, \oc8051_golden_model_1.SBUF [0]);
  and (_17241_, _17240_, _41894_);
  and (_43392_, _17241_, _17239_);
  and (_17242_, _05491_, _04595_);
  not (_17243_, _17242_);
  nor (_17244_, _05491_, \oc8051_golden_model_1.SBUF [1]);
  nor (_17245_, _17244_, _04778_);
  and (_17246_, _17245_, _17243_);
  and (_17248_, _06961_, _05491_);
  not (_17249_, \oc8051_golden_model_1.SBUF [1]);
  nor (_17250_, _05491_, _17249_);
  nor (_17251_, _17250_, _03738_);
  not (_17252_, _17251_);
  nor (_17253_, _17252_, _17248_);
  not (_17254_, _17253_);
  and (_17255_, _05491_, \oc8051_golden_model_1.ACC [1]);
  nor (_17256_, _17255_, _17250_);
  nor (_17257_, _17256_, _04708_);
  nor (_17259_, _04707_, _17249_);
  or (_17260_, _17259_, _17257_);
  and (_17261_, _17260_, _04722_);
  and (_17262_, _12262_, _05491_);
  nor (_17263_, _17262_, _17244_);
  and (_17264_, _17263_, _03850_);
  or (_17265_, _17264_, _17261_);
  and (_17266_, _17265_, _04733_);
  and (_17267_, _05491_, _04900_);
  nor (_17268_, _17267_, _17250_);
  nor (_17270_, _17268_, _04733_);
  nor (_17271_, _17270_, _17266_);
  nor (_17272_, _17271_, _03854_);
  nor (_17273_, _17256_, _03855_);
  or (_17274_, _17273_, _07927_);
  or (_17275_, _17274_, _17272_);
  and (_17276_, _17268_, _08474_);
  nor (_17277_, _17276_, _03455_);
  and (_17278_, _17277_, _17275_);
  and (_17279_, _17278_, _17254_);
  and (_17281_, _12352_, _05491_);
  or (_17282_, _17281_, _03820_);
  nor (_17283_, _17282_, _17244_);
  nor (_17284_, _17283_, _17279_);
  nor (_17285_, _17284_, _03903_);
  nor (_17286_, _17285_, _17246_);
  nor (_17287_, _17286_, _03897_);
  and (_17288_, _12366_, _05491_);
  or (_17289_, _17288_, _17250_);
  and (_17290_, _17289_, _03897_);
  nor (_17292_, _17290_, _17287_);
  nor (_17293_, _17292_, _04018_);
  nor (_17294_, _08751_, _08897_);
  nor (_17295_, _17294_, _17250_);
  and (_17296_, _08750_, _05491_);
  nor (_17297_, _17296_, _17295_);
  and (_17298_, _17297_, _04018_);
  or (_17299_, _17298_, _17293_);
  and (_17300_, _17299_, _03909_);
  and (_17301_, _12244_, _05491_);
  or (_17303_, _17301_, _17250_);
  and (_17304_, _17303_, _03908_);
  or (_17305_, _17304_, _17300_);
  and (_17306_, _17305_, _04785_);
  nor (_17307_, _17296_, _17250_);
  nor (_17308_, _17307_, _04785_);
  or (_17309_, _17308_, _17306_);
  and (_17310_, _17309_, _06567_);
  nor (_17311_, _12365_, _08897_);
  or (_17312_, _17311_, _17250_);
  and (_17314_, _17312_, _03914_);
  or (_17315_, _17314_, _17310_);
  and (_17316_, _17315_, _06572_);
  nor (_17317_, _17295_, _06572_);
  or (_17318_, _17317_, _17316_);
  nor (_17319_, _17318_, _03773_);
  nor (_17320_, _17263_, _03774_);
  or (_17321_, _17320_, _03772_);
  nor (_17322_, _17321_, _17319_);
  nor (_17323_, _17262_, _17250_);
  nor (_17325_, _17323_, _04060_);
  or (_17326_, _17325_, _17322_);
  or (_17327_, _17326_, _43156_);
  or (_17328_, _43152_, \oc8051_golden_model_1.SBUF [1]);
  and (_17329_, _17328_, _41894_);
  and (_43395_, _17329_, _17327_);
  and (_17330_, _06965_, _05491_);
  not (_17331_, \oc8051_golden_model_1.SBUF [2]);
  nor (_17332_, _05491_, _17331_);
  nor (_17333_, _17332_, _03738_);
  not (_17335_, _17333_);
  nor (_17336_, _17335_, _17330_);
  not (_17337_, _17336_);
  and (_17338_, _05491_, _05307_);
  nor (_17339_, _17338_, _17332_);
  and (_17340_, _17339_, _08474_);
  and (_17341_, _05491_, \oc8051_golden_model_1.ACC [2]);
  nor (_17342_, _17341_, _17332_);
  nor (_17343_, _17342_, _04708_);
  nor (_17344_, _04707_, _17331_);
  or (_17346_, _17344_, _17343_);
  and (_17347_, _17346_, _04722_);
  nor (_17348_, _12471_, _08897_);
  nor (_17349_, _17348_, _17332_);
  nor (_17350_, _17349_, _04722_);
  or (_17351_, _17350_, _17347_);
  and (_17352_, _17351_, _04733_);
  nor (_17353_, _17339_, _04733_);
  nor (_17354_, _17353_, _17352_);
  nor (_17355_, _17354_, _03854_);
  nor (_17357_, _17342_, _03855_);
  or (_17358_, _17357_, _07927_);
  nor (_17359_, _17358_, _17355_);
  nor (_17360_, _17359_, _17340_);
  and (_17361_, _17360_, _17337_);
  and (_17362_, _17361_, _03820_);
  nor (_17363_, _12572_, _08897_);
  nor (_17364_, _17363_, _17332_);
  nor (_17365_, _17364_, _03820_);
  or (_17366_, _17365_, _17362_);
  and (_17368_, _17366_, _04778_);
  and (_17369_, _05491_, _06495_);
  nor (_17370_, _17369_, _17332_);
  nor (_17371_, _17370_, _04778_);
  or (_17372_, _17371_, _17368_);
  and (_17373_, _17372_, _04790_);
  and (_17374_, _12586_, _05491_);
  nor (_17375_, _17374_, _17332_);
  nor (_17376_, _17375_, _04790_);
  or (_17377_, _17376_, _17373_);
  and (_17379_, _17377_, _04792_);
  and (_17380_, _08748_, _05491_);
  nor (_17381_, _17380_, _17332_);
  nor (_17382_, _17381_, _04792_);
  nor (_17383_, _17382_, _17379_);
  nor (_17384_, _17383_, _03908_);
  nor (_17385_, _17332_, _05765_);
  not (_17386_, _17385_);
  nor (_17387_, _17370_, _03909_);
  and (_17388_, _17387_, _17386_);
  nor (_17390_, _17388_, _17384_);
  nor (_17391_, _17390_, _04027_);
  nor (_17392_, _17342_, _04785_);
  and (_17393_, _17392_, _17386_);
  or (_17394_, _17393_, _17391_);
  and (_17395_, _17394_, _06567_);
  nor (_17396_, _12585_, _08897_);
  nor (_17397_, _17396_, _17332_);
  nor (_17398_, _17397_, _06567_);
  or (_17399_, _17398_, _17395_);
  and (_17401_, _17399_, _06572_);
  nor (_17402_, _08747_, _08897_);
  nor (_17403_, _17402_, _17332_);
  nor (_17404_, _17403_, _06572_);
  or (_17405_, _17404_, _03773_);
  nor (_17406_, _17405_, _17401_);
  and (_17407_, _17349_, _03773_);
  or (_17408_, _17407_, _03772_);
  nor (_17409_, _17408_, _17406_);
  and (_17410_, _12642_, _05491_);
  nor (_17412_, _17410_, _17332_);
  nor (_17413_, _17412_, _04060_);
  or (_17414_, _17413_, _17409_);
  or (_17415_, _17414_, _43156_);
  or (_17416_, _43152_, \oc8051_golden_model_1.SBUF [2]);
  and (_17417_, _17416_, _41894_);
  and (_43396_, _17417_, _17415_);
  not (_17418_, \oc8051_golden_model_1.SBUF [3]);
  nor (_17419_, _05491_, _17418_);
  and (_17420_, _05491_, \oc8051_golden_model_1.ACC [3]);
  nor (_17422_, _17420_, _17419_);
  nor (_17423_, _17422_, _04708_);
  nor (_17424_, _04707_, _17418_);
  or (_17425_, _17424_, _17423_);
  and (_17426_, _17425_, _04722_);
  nor (_17427_, _12681_, _08897_);
  nor (_17428_, _17427_, _17419_);
  nor (_17429_, _17428_, _04722_);
  or (_17430_, _17429_, _17426_);
  and (_17431_, _17430_, _04733_);
  and (_17433_, _05491_, _05119_);
  nor (_17434_, _17433_, _17419_);
  nor (_17435_, _17434_, _04733_);
  nor (_17436_, _17435_, _17431_);
  nor (_17437_, _17436_, _03854_);
  nor (_17438_, _17422_, _03855_);
  or (_17439_, _17438_, _07927_);
  or (_17440_, _17439_, _17437_);
  and (_17441_, _06964_, _05491_);
  nor (_17442_, _17419_, _03738_);
  not (_17444_, _17442_);
  nor (_17445_, _17444_, _17441_);
  and (_17446_, _17434_, _08474_);
  or (_17447_, _17446_, _03455_);
  nor (_17448_, _17447_, _17445_);
  and (_17449_, _17448_, _17440_);
  nor (_17450_, _12775_, _08897_);
  nor (_17451_, _17450_, _17419_);
  nor (_17452_, _17451_, _03820_);
  or (_17453_, _17452_, _17449_);
  and (_17455_, _17453_, _04778_);
  and (_17456_, _05491_, _06345_);
  nor (_17457_, _17456_, _17419_);
  nor (_17458_, _17457_, _04778_);
  or (_17459_, _17458_, _17455_);
  nor (_17460_, _17459_, _03897_);
  and (_17461_, _12789_, _05491_);
  or (_17462_, _17419_, _04790_);
  nor (_17463_, _17462_, _17461_);
  or (_17464_, _17463_, _04018_);
  nor (_17466_, _17464_, _17460_);
  and (_17467_, _10491_, _05491_);
  nor (_17468_, _17467_, _17419_);
  nor (_17469_, _17468_, _04792_);
  nor (_17470_, _17469_, _17466_);
  nor (_17471_, _17470_, _03908_);
  nor (_17472_, _17419_, _05622_);
  not (_17473_, _17472_);
  nor (_17474_, _17457_, _03909_);
  and (_17475_, _17474_, _17473_);
  nor (_17477_, _17475_, _17471_);
  nor (_17478_, _17477_, _04027_);
  nor (_17479_, _17422_, _04785_);
  and (_17480_, _17479_, _17473_);
  or (_17481_, _17480_, _17478_);
  and (_17482_, _17481_, _06567_);
  nor (_17483_, _12788_, _08897_);
  nor (_17484_, _17483_, _17419_);
  nor (_17485_, _17484_, _06567_);
  or (_17486_, _17485_, _17482_);
  and (_17488_, _17486_, _06572_);
  nor (_17489_, _08742_, _08897_);
  nor (_17490_, _17489_, _17419_);
  nor (_17491_, _17490_, _06572_);
  or (_17492_, _17491_, _03773_);
  nor (_17493_, _17492_, _17488_);
  and (_17494_, _17428_, _03773_);
  or (_17495_, _17494_, _03772_);
  nor (_17496_, _17495_, _17493_);
  and (_17497_, _12848_, _05491_);
  nor (_17499_, _17497_, _17419_);
  nor (_17500_, _17499_, _04060_);
  or (_17501_, _17500_, _17496_);
  or (_17502_, _17501_, _43156_);
  or (_17503_, _43152_, \oc8051_golden_model_1.SBUF [3]);
  and (_17504_, _17503_, _41894_);
  and (_43397_, _17504_, _17502_);
  not (_17505_, \oc8051_golden_model_1.SBUF [4]);
  nor (_17506_, _05491_, _17505_);
  and (_17507_, _05491_, \oc8051_golden_model_1.ACC [4]);
  nor (_17509_, _17507_, _17506_);
  nor (_17510_, _17509_, _04708_);
  nor (_17511_, _04707_, _17505_);
  or (_17512_, _17511_, _17510_);
  and (_17513_, _17512_, _04722_);
  nor (_17514_, _12891_, _08897_);
  nor (_17515_, _17514_, _17506_);
  nor (_17516_, _17515_, _04722_);
  or (_17517_, _17516_, _17513_);
  and (_17518_, _17517_, _04733_);
  and (_17520_, _05950_, _05491_);
  nor (_17521_, _17520_, _17506_);
  nor (_17522_, _17521_, _04733_);
  nor (_17523_, _17522_, _17518_);
  nor (_17524_, _17523_, _03854_);
  nor (_17525_, _17509_, _03855_);
  or (_17526_, _17525_, _07927_);
  or (_17527_, _17526_, _17524_);
  and (_17528_, _06969_, _05491_);
  nor (_17529_, _17506_, _03738_);
  not (_17531_, _17529_);
  nor (_17532_, _17531_, _17528_);
  and (_17533_, _17521_, _08474_);
  or (_17534_, _17533_, _03455_);
  nor (_17535_, _17534_, _17532_);
  and (_17536_, _17535_, _17527_);
  nor (_17537_, _12982_, _08897_);
  nor (_17538_, _17537_, _17506_);
  nor (_17539_, _17538_, _03820_);
  or (_17540_, _17539_, _17536_);
  and (_17542_, _17540_, _04778_);
  and (_17543_, _06456_, _05491_);
  nor (_17544_, _17543_, _17506_);
  nor (_17545_, _17544_, _04778_);
  or (_17546_, _17545_, _17542_);
  and (_17547_, _17546_, _04790_);
  and (_17548_, _12997_, _05491_);
  nor (_17549_, _17548_, _17506_);
  nor (_17550_, _17549_, _04790_);
  or (_17551_, _17550_, _17547_);
  and (_17553_, _17551_, _04792_);
  and (_17554_, _08741_, _05491_);
  nor (_17555_, _17554_, _17506_);
  nor (_17556_, _17555_, _04792_);
  nor (_17557_, _17556_, _17553_);
  nor (_17558_, _17557_, _03908_);
  nor (_17559_, _17506_, _08336_);
  not (_17560_, _17559_);
  nor (_17561_, _17544_, _03909_);
  and (_17562_, _17561_, _17560_);
  nor (_17564_, _17562_, _17558_);
  nor (_17565_, _17564_, _04027_);
  nor (_17566_, _17509_, _04785_);
  and (_17567_, _17566_, _17560_);
  or (_17568_, _17567_, _17565_);
  and (_17569_, _17568_, _06567_);
  nor (_17570_, _12996_, _08897_);
  nor (_17571_, _17570_, _17506_);
  nor (_17572_, _17571_, _06567_);
  or (_17573_, _17572_, _17569_);
  and (_17575_, _17573_, _06572_);
  nor (_17576_, _08740_, _08897_);
  nor (_17577_, _17576_, _17506_);
  nor (_17578_, _17577_, _06572_);
  or (_17579_, _17578_, _03773_);
  nor (_17580_, _17579_, _17575_);
  and (_17581_, _17515_, _03773_);
  or (_17582_, _17581_, _03772_);
  nor (_17583_, _17582_, _17580_);
  and (_17584_, _13056_, _05491_);
  nor (_17586_, _17584_, _17506_);
  nor (_17587_, _17586_, _04060_);
  or (_17588_, _17587_, _17583_);
  or (_17589_, _17588_, _43156_);
  or (_17590_, _43152_, \oc8051_golden_model_1.SBUF [4]);
  and (_17591_, _17590_, _41894_);
  and (_43398_, _17591_, _17589_);
  not (_17592_, \oc8051_golden_model_1.SBUF [5]);
  nor (_17593_, _05491_, _17592_);
  and (_17594_, _05491_, \oc8051_golden_model_1.ACC [5]);
  nor (_17596_, _17594_, _17593_);
  nor (_17597_, _17596_, _04708_);
  nor (_17598_, _04707_, _17592_);
  or (_17599_, _17598_, _17597_);
  and (_17600_, _17599_, _04722_);
  nor (_17601_, _13090_, _08897_);
  nor (_17602_, _17601_, _17593_);
  nor (_17603_, _17602_, _04722_);
  or (_17604_, _17603_, _17600_);
  and (_17605_, _17604_, _04733_);
  and (_17607_, _05857_, _05491_);
  nor (_17608_, _17607_, _17593_);
  nor (_17609_, _17608_, _04733_);
  nor (_17610_, _17609_, _17605_);
  nor (_17611_, _17610_, _03854_);
  nor (_17612_, _17596_, _03855_);
  or (_17613_, _17612_, _07927_);
  or (_17614_, _17613_, _17611_);
  and (_17615_, _06968_, _05491_);
  nor (_17616_, _17593_, _03738_);
  not (_17618_, _17616_);
  nor (_17619_, _17618_, _17615_);
  and (_17620_, _17608_, _08474_);
  or (_17621_, _17620_, _03455_);
  nor (_17622_, _17621_, _17619_);
  and (_17623_, _17622_, _17614_);
  nor (_17624_, _13182_, _08897_);
  nor (_17625_, _17624_, _17593_);
  nor (_17626_, _17625_, _03820_);
  or (_17627_, _17626_, _17623_);
  and (_17629_, _17627_, _04778_);
  and (_17630_, _06447_, _05491_);
  nor (_17631_, _17630_, _17593_);
  nor (_17632_, _17631_, _04778_);
  or (_17633_, _17632_, _17629_);
  nor (_17634_, _17633_, _03897_);
  and (_17635_, _13196_, _05491_);
  or (_17636_, _17593_, _04790_);
  nor (_17637_, _17636_, _17635_);
  or (_17638_, _17637_, _04018_);
  nor (_17640_, _17638_, _17634_);
  and (_17641_, _10493_, _05491_);
  nor (_17642_, _17641_, _17593_);
  nor (_17643_, _17642_, _04792_);
  nor (_17644_, _17643_, _17640_);
  nor (_17645_, _17644_, _03908_);
  nor (_17646_, _17593_, _08335_);
  not (_17647_, _17646_);
  nor (_17648_, _17631_, _03909_);
  and (_17649_, _17648_, _17647_);
  nor (_17651_, _17649_, _17645_);
  nor (_17652_, _17651_, _04027_);
  nor (_17653_, _17596_, _04785_);
  and (_17654_, _17653_, _17647_);
  nor (_17655_, _17654_, _03914_);
  not (_17656_, _17655_);
  nor (_17657_, _17656_, _17652_);
  nor (_17658_, _13195_, _08897_);
  or (_17659_, _17593_, _06567_);
  nor (_17660_, _17659_, _17658_);
  or (_17662_, _17660_, _04011_);
  nor (_17663_, _17662_, _17657_);
  nor (_17664_, _08738_, _08897_);
  nor (_17665_, _17664_, _17593_);
  nor (_17666_, _17665_, _06572_);
  nor (_17667_, _17666_, _17663_);
  nor (_17668_, _17667_, _03773_);
  nor (_17669_, _17602_, _03774_);
  or (_17670_, _17669_, _03772_);
  nor (_17671_, _17670_, _17668_);
  and (_17673_, _13255_, _05491_);
  nor (_17674_, _17673_, _17593_);
  and (_17675_, _17674_, _03772_);
  nor (_17676_, _17675_, _17671_);
  or (_17677_, _17676_, _43156_);
  or (_17678_, _43152_, \oc8051_golden_model_1.SBUF [5]);
  and (_17679_, _17678_, _41894_);
  and (_43399_, _17679_, _17677_);
  not (_17680_, \oc8051_golden_model_1.SBUF [6]);
  nor (_17681_, _05491_, _17680_);
  and (_17683_, _05491_, \oc8051_golden_model_1.ACC [6]);
  nor (_17684_, _17683_, _17681_);
  nor (_17685_, _17684_, _04708_);
  nor (_17686_, _04707_, _17680_);
  or (_17687_, _17686_, _17685_);
  and (_17688_, _17687_, _04722_);
  nor (_17689_, _13293_, _08897_);
  nor (_17690_, _17689_, _17681_);
  nor (_17691_, _17690_, _04722_);
  or (_17692_, _17691_, _17688_);
  and (_17694_, _17692_, _04733_);
  and (_17695_, _06065_, _05491_);
  nor (_17696_, _17695_, _17681_);
  nor (_17697_, _17696_, _04733_);
  nor (_17698_, _17697_, _17694_);
  nor (_17699_, _17698_, _03854_);
  nor (_17700_, _17684_, _03855_);
  or (_17701_, _17700_, _07927_);
  or (_17702_, _17701_, _17699_);
  and (_17703_, _06641_, _05491_);
  nor (_17705_, _17681_, _03738_);
  not (_17706_, _17705_);
  nor (_17707_, _17706_, _17703_);
  and (_17708_, _17696_, _08474_);
  or (_17709_, _17708_, _03455_);
  nor (_17710_, _17709_, _17707_);
  and (_17711_, _17710_, _17702_);
  nor (_17712_, _13387_, _08897_);
  nor (_17713_, _17712_, _17681_);
  nor (_17714_, _17713_, _03820_);
  or (_17716_, _17714_, _17711_);
  and (_17717_, _17716_, _04778_);
  and (_17718_, _13394_, _05491_);
  nor (_17719_, _17718_, _17681_);
  nor (_17720_, _17719_, _04778_);
  or (_17721_, _17720_, _17717_);
  and (_17722_, _17721_, _04790_);
  and (_17723_, _13402_, _05491_);
  nor (_17724_, _17723_, _17681_);
  nor (_17725_, _17724_, _04790_);
  or (_17727_, _17725_, _17722_);
  and (_17728_, _17727_, _04792_);
  and (_17729_, _08736_, _05491_);
  nor (_17730_, _17729_, _17681_);
  nor (_17731_, _17730_, _04792_);
  nor (_17732_, _17731_, _17728_);
  nor (_17733_, _17732_, _03908_);
  nor (_17734_, _17681_, _08322_);
  not (_17735_, _17734_);
  nor (_17736_, _17719_, _03909_);
  and (_17738_, _17736_, _17735_);
  nor (_17739_, _17738_, _17733_);
  nor (_17740_, _17739_, _04027_);
  nor (_17741_, _17684_, _04785_);
  and (_17742_, _17741_, _17735_);
  or (_17743_, _17742_, _17740_);
  and (_17744_, _17743_, _06567_);
  nor (_17745_, _13401_, _08897_);
  nor (_17746_, _17745_, _17681_);
  nor (_17747_, _17746_, _06567_);
  or (_17749_, _17747_, _17744_);
  and (_17750_, _17749_, _06572_);
  nor (_17751_, _08735_, _08897_);
  nor (_17752_, _17751_, _17681_);
  nor (_17753_, _17752_, _06572_);
  or (_17754_, _17753_, _03773_);
  nor (_17755_, _17754_, _17750_);
  and (_17756_, _17690_, _03773_);
  or (_17757_, _17756_, _03772_);
  nor (_17758_, _17757_, _17755_);
  nor (_17760_, _13460_, _08897_);
  nor (_17761_, _17760_, _17681_);
  nor (_17762_, _17761_, _04060_);
  or (_17763_, _17762_, _17758_);
  or (_17764_, _17763_, _43156_);
  or (_17765_, _43152_, \oc8051_golden_model_1.SBUF [6]);
  and (_17766_, _17765_, _41894_);
  and (_43400_, _17766_, _17764_);
  not (_17767_, \oc8051_golden_model_1.SCON [0]);
  nor (_17768_, _05465_, _17767_);
  and (_17770_, _05716_, _05465_);
  nor (_17771_, _17770_, _17768_);
  nor (_17772_, _17771_, _04060_);
  and (_17773_, _05465_, \oc8051_golden_model_1.ACC [0]);
  nor (_17774_, _17773_, _17768_);
  nor (_17775_, _17774_, _04708_);
  nor (_17776_, _04707_, _17767_);
  or (_17777_, _17776_, _17775_);
  and (_17778_, _17777_, _04722_);
  nor (_17779_, _17771_, _04722_);
  or (_17781_, _17779_, _17778_);
  and (_17782_, _17781_, _03764_);
  nor (_17783_, _06101_, _17767_);
  and (_17784_, _12064_, _06101_);
  nor (_17785_, _17784_, _17783_);
  nor (_17786_, _17785_, _03764_);
  nor (_17787_, _17786_, _17782_);
  nor (_17788_, _17787_, _03848_);
  and (_17789_, _05465_, _04700_);
  nor (_17790_, _17789_, _17768_);
  nor (_17792_, _17790_, _04733_);
  or (_17793_, _17792_, _17788_);
  and (_17794_, _17793_, _03855_);
  nor (_17795_, _17774_, _03855_);
  or (_17796_, _17795_, _17794_);
  and (_17797_, _17796_, _03760_);
  and (_17798_, _17768_, _03759_);
  or (_17799_, _17798_, _17797_);
  and (_17800_, _17799_, _03753_);
  nor (_17801_, _17771_, _03753_);
  or (_17803_, _17801_, _17800_);
  and (_17804_, _17803_, _03747_);
  nor (_17805_, _17783_, _14237_);
  or (_17806_, _17805_, _03747_);
  nor (_17807_, _17806_, _17785_);
  or (_17808_, _17807_, _07927_);
  or (_17809_, _17808_, _17804_);
  and (_17810_, _06962_, _05465_);
  nor (_17811_, _17768_, _03738_);
  not (_17812_, _17811_);
  nor (_17814_, _17812_, _17810_);
  and (_17815_, _17790_, _08474_);
  or (_17816_, _17815_, _03455_);
  nor (_17817_, _17816_, _17814_);
  and (_17818_, _17817_, _17809_);
  nor (_17819_, _12164_, _09001_);
  nor (_17820_, _17819_, _17768_);
  nor (_17821_, _17820_, _03820_);
  or (_17822_, _17821_, _17818_);
  and (_17823_, _17822_, _04778_);
  and (_17825_, _05465_, _06479_);
  nor (_17826_, _17825_, _17768_);
  nor (_17827_, _17826_, _04778_);
  or (_17828_, _17827_, _17823_);
  and (_17829_, _17828_, _04790_);
  and (_17830_, _12178_, _05465_);
  nor (_17831_, _17830_, _17768_);
  nor (_17832_, _17831_, _04790_);
  or (_17833_, _17832_, _17829_);
  and (_17834_, _17833_, _04792_);
  nor (_17836_, _10488_, _09001_);
  nor (_17837_, _17836_, _17768_);
  not (_17838_, _17837_);
  and (_17839_, _08753_, _05465_);
  nor (_17840_, _17839_, _04792_);
  and (_17841_, _17840_, _17838_);
  nor (_17842_, _17841_, _17834_);
  nor (_17843_, _17842_, _03908_);
  and (_17844_, _12058_, _05465_);
  or (_17845_, _17844_, _17768_);
  and (_17847_, _17845_, _03908_);
  or (_17848_, _17847_, _17843_);
  and (_17849_, _17848_, _04785_);
  nor (_17850_, _17839_, _17768_);
  nor (_17851_, _17850_, _04785_);
  or (_17852_, _17851_, _17849_);
  and (_17853_, _17852_, _06567_);
  nor (_17854_, _12177_, _09001_);
  nor (_17855_, _17854_, _17768_);
  nor (_17856_, _17855_, _06567_);
  or (_17858_, _17856_, _17853_);
  and (_17859_, _17858_, _06572_);
  nor (_17860_, _17837_, _06572_);
  or (_17861_, _17860_, _03773_);
  or (_17862_, _17861_, _17859_);
  nand (_17863_, _17771_, _03773_);
  and (_17864_, _17863_, _17862_);
  nor (_17865_, _17864_, _03374_);
  nor (_17866_, _17768_, _03375_);
  nor (_17867_, _17866_, _17865_);
  and (_17869_, _17867_, _04060_);
  nor (_17870_, _17869_, _17772_);
  nand (_17871_, _17870_, _43152_);
  or (_17872_, _43152_, \oc8051_golden_model_1.SCON [0]);
  and (_17873_, _17872_, _41894_);
  and (_43401_, _17873_, _17871_);
  not (_17874_, \oc8051_golden_model_1.SCON [1]);
  nor (_17875_, _05465_, _17874_);
  and (_17876_, _05465_, \oc8051_golden_model_1.ACC [1]);
  nor (_17877_, _17876_, _17875_);
  nor (_17879_, _17877_, _04708_);
  nor (_17880_, _04707_, _17874_);
  or (_17881_, _17880_, _17879_);
  and (_17882_, _17881_, _04722_);
  nor (_17883_, _05465_, \oc8051_golden_model_1.SCON [1]);
  and (_17884_, _12262_, _05465_);
  nor (_17885_, _17884_, _17883_);
  and (_17886_, _17885_, _03850_);
  or (_17887_, _17886_, _17882_);
  and (_17888_, _17887_, _03764_);
  nor (_17890_, _06101_, _17874_);
  and (_17891_, _12249_, _06101_);
  nor (_17892_, _17891_, _17890_);
  nor (_17893_, _17892_, _03764_);
  or (_17894_, _17893_, _17888_);
  and (_17895_, _17894_, _04733_);
  and (_17896_, _05465_, _04900_);
  nor (_17897_, _17896_, _17875_);
  nor (_17898_, _17897_, _04733_);
  or (_17899_, _17898_, _17895_);
  and (_17901_, _17899_, _03855_);
  nor (_17902_, _17877_, _03855_);
  or (_17903_, _17902_, _17901_);
  and (_17904_, _17903_, _03760_);
  and (_17905_, _12252_, _06101_);
  nor (_17906_, _17905_, _17890_);
  nor (_17907_, _17906_, _03760_);
  or (_17908_, _17907_, _03752_);
  or (_17909_, _17908_, _17904_);
  and (_17910_, _17891_, _12248_);
  or (_17912_, _17890_, _03753_);
  or (_17913_, _17912_, _17910_);
  and (_17914_, _17913_, _03747_);
  and (_17915_, _17914_, _17909_);
  nor (_17916_, _12293_, _08987_);
  nor (_17917_, _17916_, _17890_);
  nor (_17918_, _17917_, _03747_);
  or (_17919_, _17918_, _07927_);
  or (_17920_, _17919_, _17915_);
  and (_17921_, _06961_, _05465_);
  nor (_17923_, _17875_, _03738_);
  not (_17924_, _17923_);
  nor (_17925_, _17924_, _17921_);
  and (_17926_, _17897_, _08474_);
  or (_17927_, _17926_, _03455_);
  nor (_17928_, _17927_, _17925_);
  and (_17929_, _17928_, _17920_);
  nor (_17930_, _12352_, _09001_);
  nor (_17931_, _17930_, _17875_);
  nor (_17932_, _17931_, _03820_);
  nor (_17934_, _17932_, _17929_);
  nor (_17935_, _17934_, _03903_);
  and (_17936_, _05465_, _04595_);
  not (_17937_, _17936_);
  nor (_17938_, _17883_, _04778_);
  and (_17939_, _17938_, _17937_);
  nor (_17940_, _17939_, _17935_);
  nor (_17941_, _17940_, _03897_);
  and (_17942_, _12366_, _05465_);
  or (_17943_, _17942_, _17875_);
  and (_17945_, _17943_, _03897_);
  nor (_17946_, _17945_, _17941_);
  nor (_17947_, _17946_, _04018_);
  nor (_17948_, _08751_, _09001_);
  nor (_17949_, _17948_, _17875_);
  and (_17950_, _08750_, _05465_);
  nor (_17951_, _17950_, _17949_);
  and (_17952_, _17951_, _04018_);
  or (_17953_, _17952_, _17947_);
  and (_17954_, _17953_, _03909_);
  and (_17956_, _12244_, _05465_);
  or (_17957_, _17956_, _17875_);
  and (_17958_, _17957_, _03908_);
  or (_17959_, _17958_, _17954_);
  and (_17960_, _17959_, _04785_);
  nor (_17961_, _17950_, _17875_);
  nor (_17962_, _17961_, _04785_);
  or (_17963_, _17962_, _17960_);
  and (_17964_, _17963_, _06567_);
  and (_17965_, _17936_, _05669_);
  or (_17967_, _17965_, _06567_);
  nor (_17968_, _17967_, _17883_);
  or (_17969_, _17968_, _17964_);
  and (_17970_, _17969_, _06572_);
  nor (_17971_, _17949_, _06572_);
  or (_17972_, _17971_, _17970_);
  and (_17973_, _17972_, _03774_);
  and (_17974_, _17885_, _03773_);
  or (_17975_, _17974_, _17973_);
  and (_17976_, _17975_, _03375_);
  nor (_17978_, _17906_, _03375_);
  or (_17979_, _17978_, _17976_);
  and (_17980_, _17979_, _04060_);
  nor (_17981_, _17884_, _17875_);
  nor (_17982_, _17981_, _04060_);
  or (_17983_, _17982_, _17980_);
  or (_17984_, _17983_, _43156_);
  or (_17985_, _43152_, \oc8051_golden_model_1.SCON [1]);
  and (_17986_, _17985_, _41894_);
  and (_43402_, _17986_, _17984_);
  not (_17988_, \oc8051_golden_model_1.SCON [2]);
  nor (_17989_, _05465_, _17988_);
  and (_17990_, _05465_, \oc8051_golden_model_1.ACC [2]);
  nor (_17991_, _17990_, _17989_);
  nor (_17992_, _17991_, _04708_);
  nor (_17993_, _04707_, _17988_);
  or (_17994_, _17993_, _17992_);
  and (_17995_, _17994_, _04722_);
  nor (_17996_, _12471_, _09001_);
  nor (_17997_, _17996_, _17989_);
  nor (_17999_, _17997_, _04722_);
  or (_18000_, _17999_, _17995_);
  and (_18001_, _18000_, _03764_);
  nor (_18002_, _06101_, _17988_);
  and (_18003_, _12464_, _06101_);
  nor (_18004_, _18003_, _18002_);
  nor (_18005_, _18004_, _03764_);
  or (_18006_, _18005_, _18001_);
  and (_18007_, _18006_, _04733_);
  and (_18008_, _05465_, _05307_);
  nor (_18010_, _18008_, _17989_);
  nor (_18011_, _18010_, _04733_);
  or (_18012_, _18011_, _18007_);
  and (_18013_, _18012_, _03855_);
  nor (_18014_, _17991_, _03855_);
  or (_18015_, _18014_, _18013_);
  and (_18016_, _18015_, _03760_);
  and (_18017_, _12467_, _06101_);
  nor (_18018_, _18017_, _18002_);
  nor (_18019_, _18018_, _03760_);
  or (_18021_, _18019_, _18016_);
  and (_18022_, _18021_, _03753_);
  and (_18023_, _18003_, _12463_);
  or (_18024_, _18023_, _18002_);
  and (_18025_, _18024_, _03752_);
  or (_18026_, _18025_, _18022_);
  and (_18027_, _18026_, _03747_);
  nor (_18028_, _12514_, _08987_);
  nor (_18029_, _18028_, _18002_);
  nor (_18030_, _18029_, _03747_);
  or (_18032_, _18030_, _07927_);
  or (_18033_, _18032_, _18027_);
  and (_18034_, _06965_, _05465_);
  nor (_18035_, _17989_, _03738_);
  not (_18036_, _18035_);
  nor (_18037_, _18036_, _18034_);
  and (_18038_, _18010_, _08474_);
  or (_18039_, _18038_, _03455_);
  nor (_18040_, _18039_, _18037_);
  and (_18041_, _18040_, _18033_);
  nor (_18043_, _12572_, _09001_);
  nor (_18044_, _18043_, _17989_);
  nor (_18045_, _18044_, _03820_);
  or (_18046_, _18045_, _18041_);
  and (_18047_, _18046_, _04778_);
  and (_18048_, _05465_, _06495_);
  nor (_18049_, _18048_, _17989_);
  nor (_18050_, _18049_, _04778_);
  or (_18051_, _18050_, _18047_);
  and (_18052_, _18051_, _04790_);
  and (_18054_, _12586_, _05465_);
  nor (_18055_, _18054_, _17989_);
  nor (_18056_, _18055_, _04790_);
  or (_18057_, _18056_, _18052_);
  and (_18058_, _18057_, _04792_);
  and (_18059_, _08748_, _05465_);
  nor (_18060_, _18059_, _17989_);
  nor (_18061_, _18060_, _04792_);
  nor (_18062_, _18061_, _18058_);
  nor (_18063_, _18062_, _03908_);
  nor (_18065_, _17989_, _05765_);
  not (_18066_, _18065_);
  nor (_18067_, _18049_, _03909_);
  and (_18068_, _18067_, _18066_);
  nor (_18069_, _18068_, _18063_);
  nor (_18070_, _18069_, _04027_);
  nor (_18071_, _17991_, _04785_);
  and (_18072_, _18071_, _18066_);
  or (_18073_, _18072_, _18070_);
  and (_18074_, _18073_, _06567_);
  nor (_18076_, _12585_, _09001_);
  nor (_18077_, _18076_, _17989_);
  nor (_18078_, _18077_, _06567_);
  or (_18079_, _18078_, _18074_);
  and (_18080_, _18079_, _06572_);
  nor (_18081_, _08747_, _09001_);
  nor (_18082_, _18081_, _17989_);
  nor (_18083_, _18082_, _06572_);
  or (_18084_, _18083_, _18080_);
  and (_18085_, _18084_, _03774_);
  nor (_18087_, _17997_, _03774_);
  or (_18088_, _18087_, _18085_);
  and (_18089_, _18088_, _03375_);
  nor (_18090_, _18018_, _03375_);
  or (_18091_, _18090_, _18089_);
  and (_18092_, _18091_, _04060_);
  and (_18093_, _12642_, _05465_);
  nor (_18094_, _18093_, _17989_);
  nor (_18095_, _18094_, _04060_);
  or (_18096_, _18095_, _18092_);
  or (_18098_, _18096_, _43156_);
  or (_18099_, _43152_, \oc8051_golden_model_1.SCON [2]);
  and (_18100_, _18099_, _41894_);
  and (_43403_, _18100_, _18098_);
  not (_18101_, \oc8051_golden_model_1.SCON [3]);
  nor (_18102_, _05465_, _18101_);
  and (_18103_, _05465_, \oc8051_golden_model_1.ACC [3]);
  nor (_18104_, _18103_, _18102_);
  nor (_18105_, _18104_, _04708_);
  nor (_18106_, _04707_, _18101_);
  or (_18108_, _18106_, _18105_);
  and (_18109_, _18108_, _04722_);
  nor (_18110_, _12681_, _09001_);
  nor (_18111_, _18110_, _18102_);
  nor (_18112_, _18111_, _04722_);
  or (_18113_, _18112_, _18109_);
  and (_18114_, _18113_, _03764_);
  nor (_18115_, _06101_, _18101_);
  and (_18116_, _12674_, _06101_);
  nor (_18117_, _18116_, _18115_);
  nor (_18119_, _18117_, _03764_);
  or (_18120_, _18119_, _03848_);
  or (_18121_, _18120_, _18114_);
  and (_18122_, _05465_, _05119_);
  nor (_18123_, _18122_, _18102_);
  nand (_18124_, _18123_, _03848_);
  and (_18125_, _18124_, _18121_);
  and (_18126_, _18125_, _03855_);
  nor (_18127_, _18104_, _03855_);
  or (_18128_, _18127_, _18126_);
  and (_18130_, _18128_, _03760_);
  and (_18131_, _12667_, _06101_);
  nor (_18132_, _18131_, _18115_);
  nor (_18133_, _18132_, _03760_);
  or (_18134_, _18133_, _18130_);
  and (_18135_, _18134_, _03753_);
  nor (_18136_, _18115_, _12673_);
  nor (_18137_, _18136_, _18117_);
  and (_18138_, _18137_, _03752_);
  or (_18139_, _18138_, _18135_);
  and (_18141_, _18139_, _03747_);
  nor (_18142_, _12668_, _08987_);
  nor (_18143_, _18142_, _18115_);
  nor (_18144_, _18143_, _03747_);
  or (_18145_, _18144_, _07927_);
  or (_18146_, _18145_, _18141_);
  and (_18147_, _06964_, _05465_);
  nor (_18148_, _18102_, _03738_);
  not (_18149_, _18148_);
  nor (_18150_, _18149_, _18147_);
  and (_18152_, _18123_, _08474_);
  or (_18153_, _18152_, _03455_);
  nor (_18154_, _18153_, _18150_);
  and (_18155_, _18154_, _18146_);
  nor (_18156_, _12775_, _09001_);
  nor (_18157_, _18156_, _18102_);
  nor (_18158_, _18157_, _03820_);
  or (_18159_, _18158_, _18155_);
  and (_18160_, _18159_, _04778_);
  and (_18161_, _05465_, _06345_);
  nor (_18163_, _18161_, _18102_);
  nor (_18164_, _18163_, _04778_);
  or (_18165_, _18164_, _18160_);
  and (_18166_, _18165_, _04790_);
  and (_18167_, _12789_, _05465_);
  nor (_18168_, _18167_, _18102_);
  nor (_18169_, _18168_, _04790_);
  or (_18170_, _18169_, _18166_);
  and (_18171_, _18170_, _04792_);
  and (_18172_, _10491_, _05465_);
  nor (_18174_, _18172_, _18102_);
  nor (_18175_, _18174_, _04792_);
  nor (_18176_, _18175_, _18171_);
  nor (_18177_, _18176_, _03908_);
  nor (_18178_, _18102_, _05622_);
  not (_18179_, _18178_);
  nor (_18180_, _18163_, _03909_);
  and (_18181_, _18180_, _18179_);
  nor (_18182_, _18181_, _18177_);
  nor (_18183_, _18182_, _04027_);
  nor (_18185_, _18104_, _04785_);
  and (_18186_, _18185_, _18179_);
  or (_18187_, _18186_, _18183_);
  and (_18188_, _18187_, _06567_);
  nor (_18189_, _12788_, _09001_);
  nor (_18190_, _18189_, _18102_);
  nor (_18191_, _18190_, _06567_);
  or (_18192_, _18191_, _18188_);
  and (_18193_, _18192_, _06572_);
  nor (_18194_, _08742_, _09001_);
  nor (_18196_, _18194_, _18102_);
  nor (_18197_, _18196_, _06572_);
  or (_18198_, _18197_, _18193_);
  and (_18199_, _18198_, _03774_);
  nor (_18200_, _18111_, _03774_);
  or (_18201_, _18200_, _18199_);
  and (_18202_, _18201_, _03375_);
  nor (_18203_, _18132_, _03375_);
  or (_18204_, _18203_, _18202_);
  and (_18205_, _18204_, _04060_);
  and (_18207_, _12848_, _05465_);
  nor (_18208_, _18207_, _18102_);
  nor (_18209_, _18208_, _04060_);
  or (_18210_, _18209_, _18205_);
  or (_18211_, _18210_, _43156_);
  or (_18212_, _43152_, \oc8051_golden_model_1.SCON [3]);
  and (_18213_, _18212_, _41894_);
  and (_43404_, _18213_, _18211_);
  not (_18214_, \oc8051_golden_model_1.SCON [4]);
  nor (_18215_, _05465_, _18214_);
  and (_18217_, _05465_, \oc8051_golden_model_1.ACC [4]);
  nor (_18218_, _18217_, _18215_);
  nor (_18219_, _18218_, _04708_);
  nor (_18220_, _04707_, _18214_);
  or (_18221_, _18220_, _18219_);
  and (_18222_, _18221_, _04722_);
  nor (_18223_, _12891_, _09001_);
  nor (_18224_, _18223_, _18215_);
  nor (_18225_, _18224_, _04722_);
  or (_18226_, _18225_, _18222_);
  and (_18228_, _18226_, _03764_);
  nor (_18229_, _06101_, _18214_);
  and (_18230_, _12875_, _06101_);
  nor (_18231_, _18230_, _18229_);
  nor (_18232_, _18231_, _03764_);
  or (_18233_, _18232_, _03848_);
  or (_18234_, _18233_, _18228_);
  and (_18235_, _05950_, _05465_);
  nor (_18236_, _18235_, _18215_);
  nand (_18237_, _18236_, _03848_);
  and (_18239_, _18237_, _18234_);
  and (_18240_, _18239_, _03855_);
  nor (_18241_, _18218_, _03855_);
  or (_18242_, _18241_, _18240_);
  and (_18243_, _18242_, _03760_);
  and (_18244_, _12870_, _06101_);
  nor (_18245_, _18244_, _18229_);
  nor (_18246_, _18245_, _03760_);
  or (_18247_, _18246_, _03752_);
  or (_18248_, _18247_, _18243_);
  nor (_18250_, _18229_, _12874_);
  nor (_18251_, _18250_, _18231_);
  or (_18252_, _18251_, _03753_);
  and (_18253_, _18252_, _03747_);
  and (_18254_, _18253_, _18248_);
  nor (_18255_, _12872_, _08987_);
  nor (_18256_, _18255_, _18229_);
  nor (_18257_, _18256_, _03747_);
  or (_18258_, _18257_, _07927_);
  or (_18259_, _18258_, _18254_);
  and (_18261_, _06969_, _05465_);
  nor (_18262_, _18215_, _03738_);
  not (_18263_, _18262_);
  nor (_18264_, _18263_, _18261_);
  and (_18265_, _18236_, _08474_);
  or (_18266_, _18265_, _03455_);
  nor (_18267_, _18266_, _18264_);
  and (_18268_, _18267_, _18259_);
  nor (_18269_, _12982_, _09001_);
  nor (_18270_, _18269_, _18215_);
  nor (_18272_, _18270_, _03820_);
  or (_18273_, _18272_, _18268_);
  and (_18274_, _18273_, _04778_);
  and (_18275_, _06456_, _05465_);
  nor (_18276_, _18275_, _18215_);
  nor (_18277_, _18276_, _04778_);
  or (_18278_, _18277_, _18274_);
  nor (_18279_, _18278_, _03897_);
  and (_18280_, _12997_, _05465_);
  or (_18281_, _18215_, _04790_);
  nor (_18283_, _18281_, _18280_);
  or (_18284_, _18283_, _04018_);
  nor (_18285_, _18284_, _18279_);
  and (_18286_, _08741_, _05465_);
  nor (_18287_, _18286_, _18215_);
  nor (_18288_, _18287_, _04792_);
  nor (_18289_, _18288_, _18285_);
  nor (_18290_, _18289_, _03908_);
  nor (_18291_, _18215_, _08336_);
  not (_18292_, _18291_);
  nor (_18294_, _18276_, _03909_);
  and (_18295_, _18294_, _18292_);
  nor (_18296_, _18295_, _18290_);
  nor (_18297_, _18296_, _04027_);
  nor (_18298_, _18218_, _04785_);
  and (_18299_, _18298_, _18292_);
  nor (_18300_, _18299_, _03914_);
  not (_18301_, _18300_);
  nor (_18302_, _18301_, _18297_);
  nor (_18303_, _12996_, _09001_);
  or (_18305_, _18215_, _06567_);
  nor (_18306_, _18305_, _18303_);
  or (_18307_, _18306_, _04011_);
  nor (_18308_, _18307_, _18302_);
  nor (_18309_, _08740_, _09001_);
  nor (_18310_, _18309_, _18215_);
  nor (_18311_, _18310_, _06572_);
  or (_18312_, _18311_, _18308_);
  and (_18313_, _18312_, _03774_);
  nor (_18314_, _18224_, _03774_);
  or (_18316_, _18314_, _18313_);
  and (_18317_, _18316_, _03375_);
  nor (_18318_, _18245_, _03375_);
  or (_18319_, _18318_, _18317_);
  and (_18320_, _18319_, _04060_);
  and (_18321_, _13056_, _05465_);
  nor (_18322_, _18321_, _18215_);
  nor (_18323_, _18322_, _04060_);
  or (_18324_, _18323_, _18320_);
  or (_18325_, _18324_, _43156_);
  or (_18327_, _43152_, \oc8051_golden_model_1.SCON [4]);
  and (_18328_, _18327_, _41894_);
  and (_43405_, _18328_, _18325_);
  not (_18329_, \oc8051_golden_model_1.SCON [5]);
  nor (_18330_, _05465_, _18329_);
  and (_18331_, _05465_, \oc8051_golden_model_1.ACC [5]);
  nor (_18332_, _18331_, _18330_);
  nor (_18333_, _18332_, _04708_);
  nor (_18334_, _04707_, _18329_);
  or (_18335_, _18334_, _18333_);
  and (_18337_, _18335_, _04722_);
  nor (_18338_, _13090_, _09001_);
  nor (_18339_, _18338_, _18330_);
  nor (_18340_, _18339_, _04722_);
  or (_18341_, _18340_, _18337_);
  and (_18342_, _18341_, _03764_);
  nor (_18343_, _06101_, _18329_);
  and (_18344_, _13094_, _06101_);
  nor (_18345_, _18344_, _18343_);
  nor (_18346_, _18345_, _03764_);
  or (_18348_, _18346_, _03848_);
  or (_18349_, _18348_, _18342_);
  and (_18350_, _05857_, _05465_);
  nor (_18351_, _18350_, _18330_);
  nand (_18352_, _18351_, _03848_);
  and (_18353_, _18352_, _18349_);
  and (_18354_, _18353_, _03855_);
  nor (_18355_, _18332_, _03855_);
  or (_18356_, _18355_, _18354_);
  and (_18357_, _18356_, _03760_);
  and (_18359_, _13071_, _06101_);
  nor (_18360_, _18359_, _18343_);
  nor (_18361_, _18360_, _03760_);
  or (_18362_, _18361_, _18357_);
  and (_18363_, _18362_, _03753_);
  nor (_18364_, _18343_, _13109_);
  nor (_18365_, _18364_, _18345_);
  and (_18366_, _18365_, _03752_);
  or (_18367_, _18366_, _18363_);
  and (_18368_, _18367_, _03747_);
  nor (_18370_, _13073_, _08987_);
  nor (_18371_, _18370_, _18343_);
  nor (_18372_, _18371_, _03747_);
  or (_18373_, _18372_, _07927_);
  or (_18374_, _18373_, _18368_);
  and (_18375_, _06968_, _05465_);
  nor (_18376_, _18330_, _03738_);
  not (_18377_, _18376_);
  nor (_18378_, _18377_, _18375_);
  and (_18379_, _18351_, _08474_);
  or (_18381_, _18379_, _03455_);
  nor (_18382_, _18381_, _18378_);
  and (_18383_, _18382_, _18374_);
  nor (_18384_, _13182_, _09001_);
  nor (_18385_, _18384_, _18330_);
  nor (_18386_, _18385_, _03820_);
  or (_18387_, _18386_, _18383_);
  and (_18388_, _18387_, _04778_);
  and (_18389_, _06447_, _05465_);
  nor (_18390_, _18389_, _18330_);
  nor (_18392_, _18390_, _04778_);
  or (_18393_, _18392_, _18388_);
  nor (_18394_, _18393_, _03897_);
  and (_18395_, _13196_, _05465_);
  or (_18396_, _18330_, _04790_);
  nor (_18397_, _18396_, _18395_);
  or (_18398_, _18397_, _04018_);
  nor (_18399_, _18398_, _18394_);
  and (_18400_, _10493_, _05465_);
  nor (_18401_, _18400_, _18330_);
  nor (_18403_, _18401_, _04792_);
  nor (_18404_, _18403_, _18399_);
  nor (_18405_, _18404_, _03908_);
  nor (_18406_, _18330_, _08335_);
  not (_18407_, _18406_);
  nor (_18408_, _18390_, _03909_);
  and (_18409_, _18408_, _18407_);
  nor (_18410_, _18409_, _18405_);
  nor (_18411_, _18410_, _04027_);
  nor (_18412_, _18332_, _04785_);
  and (_18414_, _18412_, _18407_);
  nor (_18415_, _18414_, _03914_);
  not (_18416_, _18415_);
  nor (_18417_, _18416_, _18411_);
  nor (_18418_, _13195_, _09001_);
  or (_18419_, _18330_, _06567_);
  nor (_18420_, _18419_, _18418_);
  or (_18421_, _18420_, _04011_);
  nor (_18422_, _18421_, _18417_);
  nor (_18423_, _08738_, _09001_);
  nor (_18425_, _18423_, _18330_);
  nor (_18426_, _18425_, _06572_);
  or (_18427_, _18426_, _18422_);
  and (_18428_, _18427_, _03774_);
  nor (_18429_, _18339_, _03774_);
  or (_18430_, _18429_, _18428_);
  and (_18431_, _18430_, _03375_);
  nor (_18432_, _18360_, _03375_);
  or (_18433_, _18432_, _18431_);
  and (_18434_, _18433_, _04060_);
  and (_18436_, _13255_, _05465_);
  nor (_18437_, _18436_, _18330_);
  nor (_18438_, _18437_, _04060_);
  or (_18439_, _18438_, _18434_);
  or (_18440_, _18439_, _43156_);
  or (_18441_, _43152_, \oc8051_golden_model_1.SCON [5]);
  and (_18442_, _18441_, _41894_);
  and (_43406_, _18442_, _18440_);
  not (_18443_, \oc8051_golden_model_1.SCON [6]);
  nor (_18444_, _05465_, _18443_);
  and (_18446_, _05465_, \oc8051_golden_model_1.ACC [6]);
  nor (_18447_, _18446_, _18444_);
  nor (_18448_, _18447_, _04708_);
  nor (_18449_, _04707_, _18443_);
  or (_18450_, _18449_, _18448_);
  and (_18451_, _18450_, _04722_);
  nor (_18452_, _13293_, _09001_);
  nor (_18453_, _18452_, _18444_);
  nor (_18454_, _18453_, _04722_);
  or (_18455_, _18454_, _18451_);
  and (_18457_, _18455_, _03764_);
  nor (_18458_, _06101_, _18443_);
  and (_18459_, _13297_, _06101_);
  nor (_18460_, _18459_, _18458_);
  nor (_18461_, _18460_, _03764_);
  or (_18462_, _18461_, _03848_);
  or (_18463_, _18462_, _18457_);
  and (_18464_, _06065_, _05465_);
  nor (_18465_, _18464_, _18444_);
  nand (_18466_, _18465_, _03848_);
  and (_18468_, _18466_, _18463_);
  and (_18469_, _18468_, _03855_);
  nor (_18470_, _18447_, _03855_);
  or (_18471_, _18470_, _18469_);
  and (_18472_, _18471_, _03760_);
  and (_18473_, _13277_, _06101_);
  nor (_18474_, _18473_, _18458_);
  nor (_18475_, _18474_, _03760_);
  or (_18476_, _18475_, _03752_);
  or (_18477_, _18476_, _18472_);
  nor (_18479_, _18458_, _13312_);
  nor (_18480_, _18479_, _18460_);
  or (_18481_, _18480_, _03753_);
  and (_18482_, _18481_, _03747_);
  and (_18483_, _18482_, _18477_);
  nor (_18484_, _13279_, _08987_);
  nor (_18485_, _18484_, _18458_);
  nor (_18486_, _18485_, _03747_);
  or (_18487_, _18486_, _07927_);
  or (_18488_, _18487_, _18483_);
  and (_18490_, _06641_, _05465_);
  nor (_18491_, _18444_, _03738_);
  not (_18492_, _18491_);
  nor (_18493_, _18492_, _18490_);
  and (_18494_, _18465_, _08474_);
  or (_18495_, _18494_, _03455_);
  nor (_18496_, _18495_, _18493_);
  and (_18497_, _18496_, _18488_);
  nor (_18498_, _13387_, _09001_);
  nor (_18499_, _18498_, _18444_);
  nor (_18501_, _18499_, _03820_);
  or (_18502_, _18501_, _18497_);
  and (_18503_, _18502_, _04778_);
  and (_18504_, _13394_, _05465_);
  nor (_18505_, _18504_, _18444_);
  nor (_18506_, _18505_, _04778_);
  or (_18507_, _18506_, _18503_);
  nor (_18508_, _18507_, _03897_);
  and (_18509_, _13402_, _05465_);
  or (_18510_, _18444_, _04790_);
  nor (_18512_, _18510_, _18509_);
  or (_18513_, _18512_, _04018_);
  nor (_18514_, _18513_, _18508_);
  and (_18515_, _08736_, _05465_);
  nor (_18516_, _18515_, _18444_);
  nor (_18517_, _18516_, _04792_);
  nor (_18518_, _18517_, _18514_);
  nor (_18519_, _18518_, _03908_);
  nor (_18520_, _18444_, _08322_);
  not (_18521_, _18520_);
  nor (_18523_, _18505_, _03909_);
  and (_18524_, _18523_, _18521_);
  nor (_18525_, _18524_, _18519_);
  nor (_18526_, _18525_, _04027_);
  nor (_18527_, _18447_, _04785_);
  and (_18528_, _18527_, _18521_);
  or (_18529_, _18528_, _18526_);
  and (_18530_, _18529_, _06567_);
  nor (_18531_, _13401_, _09001_);
  nor (_18532_, _18531_, _18444_);
  nor (_18534_, _18532_, _06567_);
  or (_18535_, _18534_, _18530_);
  and (_18536_, _18535_, _06572_);
  nor (_18537_, _08735_, _09001_);
  nor (_18538_, _18537_, _18444_);
  nor (_18539_, _18538_, _06572_);
  or (_18540_, _18539_, _18536_);
  and (_18541_, _18540_, _03774_);
  nor (_18542_, _18453_, _03774_);
  or (_18543_, _18542_, _18541_);
  and (_18545_, _18543_, _03375_);
  nor (_18546_, _18474_, _03375_);
  or (_18547_, _18546_, _18545_);
  and (_18548_, _18547_, _04060_);
  nor (_18549_, _13460_, _09001_);
  nor (_18550_, _18549_, _18444_);
  nor (_18551_, _18550_, _04060_);
  or (_18552_, _18551_, _18548_);
  or (_18553_, _18552_, _43156_);
  or (_18554_, _43152_, \oc8051_golden_model_1.SCON [6]);
  and (_18556_, _18554_, _41894_);
  and (_43407_, _18556_, _18553_);
  not (_18557_, \oc8051_golden_model_1.PCON [0]);
  nor (_18558_, _05488_, _18557_);
  and (_18559_, _05716_, _05488_);
  nor (_18560_, _18559_, _18558_);
  and (_18561_, _18560_, _17157_);
  and (_18562_, _06962_, _05488_);
  nor (_18563_, _18558_, _03738_);
  not (_18564_, _18563_);
  nor (_18566_, _18564_, _18562_);
  and (_18567_, _05488_, _04700_);
  nor (_18568_, _18567_, _18558_);
  and (_18569_, _18568_, _08474_);
  and (_18570_, _05488_, \oc8051_golden_model_1.ACC [0]);
  nor (_18571_, _18570_, _18558_);
  nor (_18572_, _18571_, _04708_);
  nor (_18573_, _04707_, _18557_);
  or (_18574_, _18573_, _18572_);
  and (_18575_, _18574_, _04722_);
  nor (_18577_, _18560_, _04722_);
  or (_18578_, _18577_, _18575_);
  and (_18579_, _18578_, _04733_);
  nor (_18580_, _18568_, _04733_);
  nor (_18581_, _18580_, _18579_);
  nor (_18582_, _18581_, _03854_);
  nor (_18583_, _18571_, _03855_);
  or (_18584_, _18583_, _07927_);
  nor (_18585_, _18584_, _18582_);
  nor (_18586_, _18585_, _18569_);
  not (_18588_, _18586_);
  nor (_18589_, _18588_, _18566_);
  and (_18590_, _18589_, _03820_);
  nor (_18591_, _12164_, _09087_);
  nor (_18592_, _18591_, _18558_);
  nor (_18593_, _18592_, _03820_);
  or (_18594_, _18593_, _18590_);
  and (_18595_, _18594_, _04778_);
  and (_18596_, _05488_, _06479_);
  nor (_18597_, _18596_, _18558_);
  nor (_18599_, _18597_, _04778_);
  or (_18600_, _18599_, _18595_);
  and (_18601_, _18600_, _04790_);
  and (_18602_, _12178_, _05488_);
  nor (_18603_, _18602_, _18558_);
  nor (_18604_, _18603_, _04790_);
  or (_18605_, _18604_, _18601_);
  and (_18606_, _18605_, _04792_);
  nor (_18607_, _10488_, _09087_);
  nor (_18608_, _18607_, _18558_);
  not (_18610_, _18608_);
  and (_18611_, _08753_, _05488_);
  nor (_18612_, _18611_, _04792_);
  and (_18613_, _18612_, _18610_);
  nor (_18614_, _18613_, _18606_);
  nor (_18615_, _18614_, _03908_);
  and (_18616_, _12058_, _05488_);
  or (_18617_, _18616_, _18558_);
  and (_18618_, _18617_, _03908_);
  or (_18619_, _18618_, _18615_);
  and (_18621_, _18619_, _04785_);
  nor (_18622_, _18611_, _18558_);
  nor (_18623_, _18622_, _04785_);
  or (_18624_, _18623_, _18621_);
  and (_18625_, _18624_, _06567_);
  nor (_18626_, _12177_, _09087_);
  nor (_18627_, _18626_, _18558_);
  nor (_18628_, _18627_, _06567_);
  or (_18629_, _18628_, _18625_);
  and (_18630_, _18629_, _06572_);
  nor (_18632_, _18608_, _06572_);
  nor (_18633_, _18632_, _17157_);
  not (_18634_, _18633_);
  nor (_18635_, _18634_, _18630_);
  nor (_18636_, _18635_, _18561_);
  or (_18637_, _18636_, _43156_);
  or (_18638_, _43152_, \oc8051_golden_model_1.PCON [0]);
  and (_18639_, _18638_, _41894_);
  and (_43410_, _18639_, _18637_);
  and (_18640_, _05488_, _04595_);
  not (_18642_, _18640_);
  nor (_18643_, _05488_, \oc8051_golden_model_1.PCON [1]);
  nor (_18644_, _18643_, _04778_);
  and (_18645_, _18644_, _18642_);
  and (_18646_, _06961_, _05488_);
  not (_18647_, \oc8051_golden_model_1.PCON [1]);
  nor (_18648_, _05488_, _18647_);
  nor (_18649_, _18648_, _03738_);
  not (_18650_, _18649_);
  nor (_18651_, _18650_, _18646_);
  not (_18653_, _18651_);
  and (_18654_, _05488_, \oc8051_golden_model_1.ACC [1]);
  nor (_18655_, _18654_, _18648_);
  nor (_18656_, _18655_, _04708_);
  nor (_18657_, _04707_, _18647_);
  or (_18658_, _18657_, _18656_);
  and (_18659_, _18658_, _04722_);
  and (_18660_, _12262_, _05488_);
  nor (_18661_, _18660_, _18643_);
  and (_18662_, _18661_, _03850_);
  or (_18664_, _18662_, _18659_);
  and (_18665_, _18664_, _04733_);
  and (_18666_, _05488_, _04900_);
  nor (_18667_, _18666_, _18648_);
  nor (_18668_, _18667_, _04733_);
  nor (_18669_, _18668_, _18665_);
  nor (_18670_, _18669_, _03854_);
  nor (_18671_, _18655_, _03855_);
  or (_18672_, _18671_, _07927_);
  or (_18673_, _18672_, _18670_);
  and (_18675_, _18667_, _08474_);
  nor (_18676_, _18675_, _03455_);
  and (_18677_, _18676_, _18673_);
  and (_18678_, _18677_, _18653_);
  not (_18679_, _18643_);
  and (_18680_, _12352_, _05488_);
  nor (_18681_, _18680_, _03820_);
  and (_18682_, _18681_, _18679_);
  nor (_18683_, _18682_, _18678_);
  nor (_18684_, _18683_, _03903_);
  nor (_18686_, _18684_, _18645_);
  nor (_18687_, _18686_, _03897_);
  nor (_18688_, _12366_, _09087_);
  nor (_18689_, _18688_, _04790_);
  and (_18690_, _18689_, _18679_);
  nor (_18691_, _18690_, _18687_);
  nor (_18692_, _18691_, _04018_);
  nor (_18693_, _08751_, _09087_);
  nor (_18694_, _18693_, _18648_);
  and (_18695_, _08750_, _05488_);
  nor (_18697_, _18695_, _18694_);
  and (_18698_, _18697_, _04018_);
  or (_18699_, _18698_, _18692_);
  and (_18700_, _18699_, _03909_);
  and (_18701_, _12244_, _05488_);
  or (_18702_, _18701_, _18648_);
  and (_18703_, _18702_, _03908_);
  or (_18704_, _18703_, _18700_);
  and (_18705_, _18704_, _04785_);
  nor (_18706_, _18695_, _18648_);
  nor (_18708_, _18706_, _04785_);
  or (_18709_, _18708_, _18705_);
  and (_18710_, _18709_, _06567_);
  and (_18711_, _18640_, _05669_);
  nor (_18712_, _18711_, _06567_);
  and (_18713_, _18712_, _18679_);
  or (_18714_, _18713_, _18710_);
  and (_18715_, _18714_, _06572_);
  nor (_18716_, _18694_, _06572_);
  or (_18717_, _18716_, _18715_);
  nor (_18719_, _18717_, _03773_);
  nor (_18720_, _18661_, _03774_);
  or (_18721_, _18720_, _03772_);
  nor (_18722_, _18721_, _18719_);
  nor (_18723_, _18660_, _18648_);
  nor (_18724_, _18723_, _04060_);
  or (_18725_, _18724_, _18722_);
  or (_18726_, _18725_, _43156_);
  or (_18727_, _43152_, \oc8051_golden_model_1.PCON [1]);
  and (_18728_, _18727_, _41894_);
  and (_43411_, _18728_, _18726_);
  and (_18730_, _06965_, _05488_);
  not (_18731_, \oc8051_golden_model_1.PCON [2]);
  nor (_18732_, _05488_, _18731_);
  nor (_18733_, _18732_, _03738_);
  not (_18734_, _18733_);
  nor (_18735_, _18734_, _18730_);
  and (_18736_, _05488_, \oc8051_golden_model_1.ACC [2]);
  nor (_18737_, _18736_, _18732_);
  nor (_18738_, _18737_, _04708_);
  nor (_18740_, _04707_, _18731_);
  or (_18741_, _18740_, _18738_);
  and (_18742_, _18741_, _04722_);
  nor (_18743_, _12471_, _09087_);
  nor (_18744_, _18743_, _18732_);
  nor (_18745_, _18744_, _04722_);
  or (_18746_, _18745_, _18742_);
  and (_18747_, _18746_, _04733_);
  and (_18748_, _05488_, _05307_);
  nor (_18749_, _18748_, _18732_);
  nor (_18751_, _18749_, _04733_);
  nor (_18752_, _18751_, _18747_);
  nor (_18753_, _18752_, _03854_);
  nor (_18754_, _18737_, _03855_);
  or (_18755_, _18754_, _07927_);
  nor (_18756_, _18755_, _18753_);
  and (_18757_, _18749_, _08474_);
  or (_18758_, _18757_, _03455_);
  or (_18759_, _18758_, _18756_);
  nor (_18760_, _18759_, _18735_);
  nor (_18762_, _12572_, _09087_);
  nor (_18763_, _18762_, _18732_);
  nor (_18764_, _18763_, _03820_);
  or (_18765_, _18764_, _18760_);
  and (_18766_, _18765_, _04778_);
  and (_18767_, _05488_, _06495_);
  nor (_18768_, _18767_, _18732_);
  nor (_18769_, _18768_, _04778_);
  or (_18770_, _18769_, _18766_);
  and (_18771_, _18770_, _04790_);
  and (_18773_, _12586_, _05488_);
  nor (_18774_, _18773_, _18732_);
  nor (_18775_, _18774_, _04790_);
  or (_18776_, _18775_, _18771_);
  and (_18777_, _18776_, _04792_);
  and (_18778_, _08748_, _05488_);
  nor (_18779_, _18778_, _18732_);
  nor (_18780_, _18779_, _04792_);
  nor (_18781_, _18780_, _18777_);
  nor (_18782_, _18781_, _03908_);
  nor (_18784_, _18732_, _05765_);
  not (_18785_, _18784_);
  nor (_18786_, _18768_, _03909_);
  and (_18787_, _18786_, _18785_);
  nor (_18788_, _18787_, _18782_);
  nor (_18789_, _18788_, _04027_);
  nor (_18790_, _18737_, _04785_);
  and (_18791_, _18790_, _18785_);
  or (_18792_, _18791_, _18789_);
  and (_18793_, _18792_, _06567_);
  nor (_18795_, _12585_, _09087_);
  nor (_18796_, _18795_, _18732_);
  nor (_18797_, _18796_, _06567_);
  or (_18798_, _18797_, _18793_);
  and (_18799_, _18798_, _06572_);
  nor (_18800_, _08747_, _09087_);
  nor (_18801_, _18800_, _18732_);
  nor (_18802_, _18801_, _06572_);
  or (_18803_, _18802_, _03773_);
  nor (_18804_, _18803_, _18799_);
  and (_18806_, _18744_, _03773_);
  or (_18807_, _18806_, _03772_);
  nor (_18808_, _18807_, _18804_);
  and (_18809_, _12642_, _05488_);
  nor (_18810_, _18809_, _18732_);
  nor (_18811_, _18810_, _04060_);
  or (_18812_, _18811_, _18808_);
  or (_18813_, _18812_, _43156_);
  or (_18814_, _43152_, \oc8051_golden_model_1.PCON [2]);
  and (_18815_, _18814_, _41894_);
  and (_43412_, _18815_, _18813_);
  not (_18817_, \oc8051_golden_model_1.PCON [3]);
  nor (_18818_, _05488_, _18817_);
  and (_18819_, _05488_, \oc8051_golden_model_1.ACC [3]);
  nor (_18820_, _18819_, _18818_);
  nor (_18821_, _18820_, _04708_);
  nor (_18822_, _04707_, _18817_);
  or (_18823_, _18822_, _18821_);
  and (_18824_, _18823_, _04722_);
  nor (_18825_, _12681_, _09087_);
  nor (_18827_, _18825_, _18818_);
  nor (_18828_, _18827_, _04722_);
  or (_18829_, _18828_, _18824_);
  and (_18830_, _18829_, _04733_);
  and (_18831_, _05488_, _05119_);
  nor (_18832_, _18831_, _18818_);
  nor (_18833_, _18832_, _04733_);
  nor (_18834_, _18833_, _18830_);
  nor (_18835_, _18834_, _03854_);
  nor (_18836_, _18820_, _03855_);
  or (_18838_, _18836_, _07927_);
  or (_18839_, _18838_, _18835_);
  and (_18840_, _06964_, _05488_);
  nor (_18841_, _18818_, _03738_);
  not (_18842_, _18841_);
  nor (_18843_, _18842_, _18840_);
  and (_18844_, _18832_, _08474_);
  or (_18845_, _18844_, _03455_);
  nor (_18846_, _18845_, _18843_);
  and (_18847_, _18846_, _18839_);
  nor (_18849_, _12775_, _09087_);
  nor (_18850_, _18849_, _18818_);
  nor (_18851_, _18850_, _03820_);
  or (_18852_, _18851_, _18847_);
  and (_18853_, _18852_, _04778_);
  and (_18854_, _05488_, _06345_);
  nor (_18855_, _18854_, _18818_);
  nor (_18856_, _18855_, _04778_);
  or (_18857_, _18856_, _18853_);
  nor (_18858_, _18857_, _03897_);
  and (_18860_, _12789_, _05488_);
  or (_18861_, _18818_, _04790_);
  nor (_18862_, _18861_, _18860_);
  or (_18863_, _18862_, _04018_);
  nor (_18864_, _18863_, _18858_);
  and (_18865_, _10491_, _05488_);
  nor (_18866_, _18865_, _18818_);
  nor (_18867_, _18866_, _04792_);
  nor (_18868_, _18867_, _18864_);
  nor (_18869_, _18868_, _03908_);
  nor (_18871_, _18818_, _05622_);
  not (_18872_, _18871_);
  nor (_18873_, _18855_, _03909_);
  and (_18874_, _18873_, _18872_);
  nor (_18875_, _18874_, _18869_);
  nor (_18876_, _18875_, _04027_);
  nor (_18877_, _18820_, _04785_);
  and (_18878_, _18877_, _18872_);
  or (_18879_, _18878_, _18876_);
  and (_18880_, _18879_, _06567_);
  nor (_18882_, _12788_, _09087_);
  nor (_18883_, _18882_, _18818_);
  nor (_18884_, _18883_, _06567_);
  or (_18885_, _18884_, _18880_);
  and (_18886_, _18885_, _06572_);
  nor (_18887_, _08742_, _09087_);
  nor (_18888_, _18887_, _18818_);
  nor (_18889_, _18888_, _06572_);
  or (_18890_, _18889_, _03773_);
  nor (_18891_, _18890_, _18886_);
  and (_18893_, _18827_, _03773_);
  or (_18894_, _18893_, _03772_);
  nor (_18895_, _18894_, _18891_);
  and (_18896_, _12848_, _05488_);
  nor (_18897_, _18896_, _18818_);
  nor (_18898_, _18897_, _04060_);
  or (_18899_, _18898_, _18895_);
  or (_18900_, _18899_, _43156_);
  or (_18901_, _43152_, \oc8051_golden_model_1.PCON [3]);
  and (_18902_, _18901_, _41894_);
  and (_43415_, _18902_, _18900_);
  not (_18904_, \oc8051_golden_model_1.PCON [4]);
  nor (_18905_, _05488_, _18904_);
  and (_18906_, _05488_, \oc8051_golden_model_1.ACC [4]);
  nor (_18907_, _18906_, _18905_);
  nor (_18908_, _18907_, _04708_);
  nor (_18909_, _04707_, _18904_);
  or (_18910_, _18909_, _18908_);
  and (_18911_, _18910_, _04722_);
  nor (_18912_, _12891_, _09087_);
  nor (_18914_, _18912_, _18905_);
  nor (_18915_, _18914_, _04722_);
  or (_18916_, _18915_, _18911_);
  and (_18917_, _18916_, _04733_);
  and (_18918_, _05950_, _05488_);
  nor (_18919_, _18918_, _18905_);
  nor (_18920_, _18919_, _04733_);
  nor (_18921_, _18920_, _18917_);
  nor (_18922_, _18921_, _03854_);
  nor (_18923_, _18907_, _03855_);
  or (_18925_, _18923_, _07927_);
  or (_18926_, _18925_, _18922_);
  and (_18927_, _06969_, _05488_);
  nor (_18928_, _18905_, _03738_);
  not (_18929_, _18928_);
  nor (_18930_, _18929_, _18927_);
  and (_18931_, _18919_, _08474_);
  or (_18932_, _18931_, _03455_);
  nor (_18933_, _18932_, _18930_);
  and (_18934_, _18933_, _18926_);
  nor (_18936_, _12982_, _09087_);
  nor (_18937_, _18936_, _18905_);
  nor (_18938_, _18937_, _03820_);
  or (_18939_, _18938_, _18934_);
  and (_18940_, _18939_, _04778_);
  and (_18941_, _06456_, _05488_);
  nor (_18942_, _18941_, _18905_);
  nor (_18943_, _18942_, _04778_);
  or (_18944_, _18943_, _18940_);
  nor (_18945_, _18944_, _03897_);
  and (_18947_, _12997_, _05488_);
  or (_18948_, _18905_, _04790_);
  nor (_18949_, _18948_, _18947_);
  or (_18950_, _18949_, _04018_);
  nor (_18951_, _18950_, _18945_);
  and (_18952_, _08741_, _05488_);
  nor (_18953_, _18952_, _18905_);
  nor (_18954_, _18953_, _04792_);
  nor (_18955_, _18954_, _18951_);
  nor (_18956_, _18955_, _03908_);
  nor (_18958_, _18905_, _08336_);
  not (_18959_, _18958_);
  nor (_18960_, _18942_, _03909_);
  and (_18961_, _18960_, _18959_);
  nor (_18962_, _18961_, _18956_);
  nor (_18963_, _18962_, _04027_);
  nor (_18964_, _18907_, _04785_);
  and (_18965_, _18964_, _18959_);
  or (_18966_, _18965_, _18963_);
  and (_18967_, _18966_, _06567_);
  nor (_18969_, _12996_, _09087_);
  nor (_18970_, _18969_, _18905_);
  nor (_18971_, _18970_, _06567_);
  or (_18972_, _18971_, _18967_);
  and (_18973_, _18972_, _06572_);
  nor (_18974_, _08740_, _09087_);
  nor (_18975_, _18974_, _18905_);
  nor (_18976_, _18975_, _06572_);
  or (_18977_, _18976_, _03773_);
  nor (_18978_, _18977_, _18973_);
  and (_18980_, _18914_, _03773_);
  or (_18981_, _18980_, _03772_);
  nor (_18982_, _18981_, _18978_);
  and (_18983_, _13056_, _05488_);
  nor (_18984_, _18983_, _18905_);
  nor (_18985_, _18984_, _04060_);
  or (_18986_, _18985_, _18982_);
  or (_18987_, _18986_, _43156_);
  or (_18988_, _43152_, \oc8051_golden_model_1.PCON [4]);
  and (_18989_, _18988_, _41894_);
  and (_43416_, _18989_, _18987_);
  not (_18991_, \oc8051_golden_model_1.PCON [5]);
  nor (_18992_, _05488_, _18991_);
  and (_18993_, _05488_, \oc8051_golden_model_1.ACC [5]);
  nor (_18994_, _18993_, _18992_);
  nor (_18995_, _18994_, _04708_);
  nor (_18996_, _04707_, _18991_);
  or (_18997_, _18996_, _18995_);
  and (_18998_, _18997_, _04722_);
  nor (_18999_, _13090_, _09087_);
  nor (_19001_, _18999_, _18992_);
  nor (_19002_, _19001_, _04722_);
  or (_19003_, _19002_, _18998_);
  and (_19004_, _19003_, _04733_);
  and (_19005_, _05857_, _05488_);
  nor (_19006_, _19005_, _18992_);
  nor (_19007_, _19006_, _04733_);
  nor (_19008_, _19007_, _19004_);
  nor (_19009_, _19008_, _03854_);
  nor (_19010_, _18994_, _03855_);
  or (_19012_, _19010_, _07927_);
  or (_19013_, _19012_, _19009_);
  and (_19014_, _06968_, _05488_);
  nor (_19015_, _18992_, _03738_);
  not (_19016_, _19015_);
  nor (_19017_, _19016_, _19014_);
  and (_19018_, _19006_, _08474_);
  or (_19019_, _19018_, _03455_);
  nor (_19020_, _19019_, _19017_);
  and (_19021_, _19020_, _19013_);
  nor (_19023_, _13182_, _09087_);
  nor (_19024_, _19023_, _18992_);
  nor (_19025_, _19024_, _03820_);
  or (_19026_, _19025_, _19021_);
  and (_19027_, _19026_, _04778_);
  and (_19028_, _06447_, _05488_);
  nor (_19029_, _19028_, _18992_);
  nor (_19030_, _19029_, _04778_);
  or (_19031_, _19030_, _19027_);
  nor (_19032_, _19031_, _03897_);
  and (_19034_, _13196_, _05488_);
  or (_19035_, _18992_, _04790_);
  nor (_19036_, _19035_, _19034_);
  or (_19037_, _19036_, _04018_);
  nor (_19038_, _19037_, _19032_);
  and (_19039_, _10493_, _05488_);
  nor (_19040_, _19039_, _18992_);
  nor (_19041_, _19040_, _04792_);
  nor (_19042_, _19041_, _19038_);
  nor (_19043_, _19042_, _03908_);
  nor (_19045_, _18992_, _08335_);
  not (_19046_, _19045_);
  nor (_19047_, _19029_, _03909_);
  and (_19048_, _19047_, _19046_);
  nor (_19049_, _19048_, _19043_);
  nor (_19050_, _19049_, _04027_);
  nor (_19051_, _18994_, _04785_);
  and (_19052_, _19051_, _19046_);
  or (_19053_, _19052_, _19050_);
  and (_19054_, _19053_, _06567_);
  nor (_19056_, _13195_, _09087_);
  nor (_19057_, _19056_, _18992_);
  nor (_19058_, _19057_, _06567_);
  or (_19059_, _19058_, _19054_);
  and (_19060_, _19059_, _06572_);
  nor (_19061_, _08738_, _09087_);
  nor (_19062_, _19061_, _18992_);
  nor (_19063_, _19062_, _06572_);
  nor (_19064_, _19063_, _19060_);
  nor (_19065_, _19064_, _03773_);
  nor (_19067_, _19001_, _03774_);
  or (_19068_, _19067_, _03772_);
  nor (_19069_, _19068_, _19065_);
  and (_19070_, _13255_, _05488_);
  nor (_19071_, _19070_, _18992_);
  and (_19072_, _19071_, _03772_);
  nor (_19073_, _19072_, _19069_);
  or (_19074_, _19073_, _43156_);
  or (_19075_, _43152_, \oc8051_golden_model_1.PCON [5]);
  and (_19076_, _19075_, _41894_);
  and (_43417_, _19076_, _19074_);
  not (_19078_, \oc8051_golden_model_1.PCON [6]);
  nor (_19079_, _05488_, _19078_);
  and (_19080_, _05488_, \oc8051_golden_model_1.ACC [6]);
  nor (_19081_, _19080_, _19079_);
  nor (_19082_, _19081_, _04708_);
  nor (_19083_, _04707_, _19078_);
  or (_19084_, _19083_, _19082_);
  and (_19085_, _19084_, _04722_);
  nor (_19086_, _13293_, _09087_);
  nor (_19088_, _19086_, _19079_);
  nor (_19089_, _19088_, _04722_);
  or (_19090_, _19089_, _19085_);
  and (_19091_, _19090_, _04733_);
  and (_19092_, _06065_, _05488_);
  nor (_19093_, _19092_, _19079_);
  nor (_19094_, _19093_, _04733_);
  nor (_19095_, _19094_, _19091_);
  nor (_19096_, _19095_, _03854_);
  nor (_19097_, _19081_, _03855_);
  or (_19099_, _19097_, _07927_);
  or (_19100_, _19099_, _19096_);
  and (_19101_, _06641_, _05488_);
  nor (_19102_, _19079_, _03738_);
  not (_19103_, _19102_);
  nor (_19104_, _19103_, _19101_);
  and (_19105_, _19093_, _08474_);
  or (_19106_, _19105_, _03455_);
  nor (_19107_, _19106_, _19104_);
  and (_19108_, _19107_, _19100_);
  nor (_19110_, _13387_, _09087_);
  nor (_19111_, _19110_, _19079_);
  nor (_19112_, _19111_, _03820_);
  or (_19113_, _19112_, _19108_);
  and (_19114_, _19113_, _04778_);
  and (_19115_, _13394_, _05488_);
  nor (_19116_, _19115_, _19079_);
  nor (_19117_, _19116_, _04778_);
  or (_19118_, _19117_, _19114_);
  and (_19119_, _19118_, _04790_);
  and (_19121_, _13402_, _05488_);
  nor (_19122_, _19121_, _19079_);
  nor (_19123_, _19122_, _04790_);
  or (_19124_, _19123_, _19119_);
  and (_19125_, _19124_, _04792_);
  and (_19126_, _08736_, _05488_);
  nor (_19127_, _19126_, _19079_);
  nor (_19128_, _19127_, _04792_);
  nor (_19129_, _19128_, _19125_);
  nor (_19130_, _19129_, _03908_);
  nor (_19132_, _19079_, _08322_);
  not (_19133_, _19132_);
  nor (_19134_, _19116_, _03909_);
  and (_19135_, _19134_, _19133_);
  nor (_19136_, _19135_, _19130_);
  nor (_19137_, _19136_, _04027_);
  nor (_19138_, _19081_, _04785_);
  and (_19139_, _19138_, _19133_);
  nor (_19140_, _19139_, _03914_);
  not (_19141_, _19140_);
  nor (_19143_, _19141_, _19137_);
  nor (_19144_, _13401_, _09087_);
  or (_19145_, _19079_, _06567_);
  nor (_19146_, _19145_, _19144_);
  or (_19147_, _19146_, _04011_);
  nor (_19148_, _19147_, _19143_);
  nor (_19149_, _08735_, _09087_);
  nor (_19150_, _19149_, _19079_);
  nor (_19151_, _19150_, _06572_);
  or (_19152_, _19151_, _03773_);
  nor (_19154_, _19152_, _19148_);
  and (_19155_, _19088_, _03773_);
  or (_19156_, _19155_, _03772_);
  nor (_19157_, _19156_, _19154_);
  nor (_19158_, _13460_, _09087_);
  nor (_19159_, _19158_, _19079_);
  nor (_19160_, _19159_, _04060_);
  or (_19161_, _19160_, _19157_);
  or (_19162_, _19161_, _43156_);
  or (_19163_, _43152_, \oc8051_golden_model_1.PCON [6]);
  and (_19165_, _19163_, _41894_);
  and (_43418_, _19165_, _19162_);
  not (_19166_, \oc8051_golden_model_1.TCON [0]);
  nor (_19167_, _05447_, _19166_);
  and (_19168_, _05716_, _05447_);
  nor (_19169_, _19168_, _19167_);
  nor (_19170_, _19169_, _04060_);
  and (_19171_, _06962_, _05447_);
  nor (_19172_, _19167_, _03738_);
  not (_19173_, _19172_);
  nor (_19175_, _19173_, _19171_);
  nor (_19176_, _19169_, _04722_);
  nor (_19177_, _04707_, _19166_);
  and (_19178_, _05447_, \oc8051_golden_model_1.ACC [0]);
  nor (_19179_, _19178_, _19167_);
  nor (_19180_, _19179_, _04708_);
  nor (_19181_, _19180_, _19177_);
  nor (_19182_, _19181_, _03850_);
  or (_19183_, _19182_, _03763_);
  nor (_19184_, _19183_, _19176_);
  and (_19186_, _12064_, _06085_);
  nor (_19187_, _06085_, _19166_);
  or (_19188_, _19187_, _03764_);
  nor (_19189_, _19188_, _19186_);
  or (_19190_, _19189_, _03848_);
  nor (_19191_, _19190_, _19184_);
  and (_19192_, _05447_, _04700_);
  nor (_19193_, _19192_, _19167_);
  nor (_19194_, _19193_, _04733_);
  or (_19195_, _19194_, _19191_);
  and (_19197_, _19195_, _03855_);
  nor (_19198_, _19179_, _03855_);
  or (_19199_, _19198_, _19197_);
  and (_19200_, _19199_, _03760_);
  and (_19201_, _19167_, _03759_);
  or (_19202_, _19201_, _19200_);
  and (_19203_, _19202_, _03753_);
  nor (_19204_, _19169_, _03753_);
  or (_19205_, _19204_, _19203_);
  and (_19206_, _19205_, _03747_);
  and (_19208_, _19186_, _14237_);
  nor (_19209_, _19208_, _19187_);
  nor (_19210_, _19209_, _03747_);
  or (_19211_, _19210_, _07927_);
  nor (_19212_, _19211_, _19206_);
  and (_19213_, _19193_, _08474_);
  or (_19214_, _19213_, _03455_);
  or (_19215_, _19214_, _19212_);
  nor (_19216_, _19215_, _19175_);
  nor (_19217_, _12164_, _09186_);
  nor (_19219_, _19217_, _19167_);
  nor (_19220_, _19219_, _03820_);
  or (_19221_, _19220_, _19216_);
  and (_19222_, _19221_, _04778_);
  and (_19223_, _05447_, _06479_);
  nor (_19224_, _19223_, _19167_);
  nor (_19225_, _19224_, _04778_);
  or (_19226_, _19225_, _19222_);
  and (_19227_, _19226_, _04790_);
  and (_19228_, _12178_, _05447_);
  nor (_19230_, _19228_, _19167_);
  nor (_19231_, _19230_, _04790_);
  or (_19232_, _19231_, _19227_);
  and (_19233_, _19232_, _04792_);
  nor (_19234_, _10488_, _09186_);
  nor (_19235_, _19234_, _19167_);
  nand (_19236_, _08753_, _05447_);
  nand (_19237_, _19236_, _04018_);
  nor (_19238_, _19237_, _19235_);
  nor (_19239_, _19238_, _19233_);
  nor (_19241_, _19239_, _03908_);
  nor (_19242_, _19224_, _03909_);
  not (_19243_, _19242_);
  nor (_19244_, _19243_, _19168_);
  nor (_19245_, _19244_, _04027_);
  not (_19246_, _19245_);
  nor (_19247_, _19246_, _19241_);
  nor (_19248_, _19167_, _04785_);
  and (_19249_, _19248_, _19236_);
  nor (_19250_, _19249_, _19247_);
  and (_19252_, _19250_, _06567_);
  nor (_19253_, _12177_, _09186_);
  nor (_19254_, _19253_, _19167_);
  nor (_19255_, _19254_, _06567_);
  or (_19256_, _19255_, _19252_);
  and (_19257_, _19256_, _06572_);
  nor (_19258_, _19235_, _06572_);
  or (_19259_, _19258_, _03773_);
  or (_19260_, _19259_, _19257_);
  nand (_19261_, _19169_, _03773_);
  and (_19263_, _19261_, _19260_);
  nor (_19264_, _19263_, _03374_);
  nor (_19265_, _19167_, _03375_);
  nor (_19266_, _19265_, _19264_);
  and (_19267_, _19266_, _04060_);
  nor (_19268_, _19267_, _19170_);
  nand (_19269_, _19268_, _43152_);
  or (_19270_, _43152_, \oc8051_golden_model_1.TCON [0]);
  and (_19271_, _19270_, _41894_);
  and (_43419_, _19271_, _19269_);
  not (_19273_, \oc8051_golden_model_1.TCON [1]);
  nor (_19274_, _05447_, _19273_);
  nor (_19275_, _08751_, _09186_);
  or (_19276_, _19275_, _19274_);
  or (_19277_, _19276_, _06572_);
  nand (_19278_, _05447_, _04595_);
  or (_19279_, _05447_, \oc8051_golden_model_1.TCON [1]);
  and (_19280_, _19279_, _03903_);
  and (_19281_, _19280_, _19278_);
  and (_19282_, _05447_, _04900_);
  or (_19284_, _19282_, _19274_);
  or (_19285_, _19284_, _04733_);
  and (_19286_, _12262_, _05447_);
  not (_19287_, _19286_);
  and (_19288_, _19287_, _19279_);
  or (_19289_, _19288_, _04722_);
  and (_19290_, _05447_, \oc8051_golden_model_1.ACC [1]);
  or (_19291_, _19290_, _19274_);
  and (_19292_, _19291_, _04707_);
  nor (_19293_, _04707_, _19273_);
  or (_19295_, _19293_, _03850_);
  or (_19296_, _19295_, _19292_);
  and (_19297_, _19296_, _03764_);
  and (_19298_, _19297_, _19289_);
  nor (_19299_, _06085_, _19273_);
  and (_19300_, _12249_, _06085_);
  or (_19301_, _19300_, _19299_);
  and (_19302_, _19301_, _03763_);
  or (_19303_, _19302_, _03848_);
  or (_19304_, _19303_, _19298_);
  and (_19306_, _19304_, _19285_);
  or (_19307_, _19306_, _03854_);
  or (_19308_, _19291_, _03855_);
  and (_19309_, _19308_, _03760_);
  and (_19310_, _19309_, _19307_);
  and (_19311_, _12252_, _06085_);
  or (_19312_, _19311_, _19299_);
  and (_19313_, _19312_, _03759_);
  or (_19314_, _19313_, _03752_);
  or (_19315_, _19314_, _19310_);
  and (_19317_, _19300_, _12248_);
  or (_19318_, _19299_, _03753_);
  or (_19319_, _19318_, _19317_);
  and (_19320_, _19319_, _03747_);
  and (_19321_, _19320_, _19315_);
  nor (_19322_, _12293_, _09172_);
  or (_19323_, _19322_, _19299_);
  and (_19324_, _19323_, _03746_);
  or (_19325_, _19324_, _07927_);
  or (_19326_, _19325_, _19321_);
  and (_19328_, _06961_, _05447_);
  or (_19329_, _19274_, _03738_);
  or (_19330_, _19329_, _19328_);
  or (_19331_, _19284_, _07925_);
  and (_19332_, _19331_, _03820_);
  and (_19333_, _19332_, _19330_);
  and (_19334_, _19333_, _19326_);
  nor (_19335_, _12352_, _09186_);
  or (_19336_, _19335_, _19274_);
  and (_19337_, _19336_, _03455_);
  or (_19339_, _19337_, _19334_);
  and (_19340_, _19339_, _04778_);
  or (_19341_, _19340_, _19281_);
  and (_19342_, _19341_, _04790_);
  or (_19343_, _12366_, _09186_);
  and (_19344_, _19279_, _03897_);
  and (_19345_, _19344_, _19343_);
  or (_19346_, _19345_, _04018_);
  or (_19347_, _19346_, _19342_);
  and (_19348_, _08752_, _05447_);
  or (_19350_, _19348_, _19274_);
  or (_19351_, _19350_, _04792_);
  and (_19352_, _19351_, _03909_);
  and (_19353_, _19352_, _19347_);
  or (_19354_, _12244_, _09186_);
  and (_19355_, _19279_, _03908_);
  and (_19356_, _19355_, _19354_);
  or (_19357_, _19356_, _04027_);
  or (_19358_, _19357_, _19353_);
  and (_19359_, _08750_, _05447_);
  or (_19361_, _19274_, _04785_);
  or (_19362_, _19361_, _19359_);
  and (_19363_, _19362_, _06567_);
  and (_19364_, _19363_, _19358_);
  or (_19365_, _19278_, _08366_);
  and (_19366_, _19279_, _03914_);
  and (_19367_, _19366_, _19365_);
  or (_19368_, _19367_, _04011_);
  or (_19369_, _19368_, _19364_);
  and (_19370_, _19369_, _19277_);
  or (_19372_, _19370_, _03773_);
  or (_19373_, _19288_, _03774_);
  and (_19374_, _19373_, _03375_);
  and (_19375_, _19374_, _19372_);
  and (_19376_, _19312_, _03374_);
  or (_19377_, _19376_, _03772_);
  or (_19378_, _19377_, _19375_);
  or (_19379_, _19286_, _19274_);
  or (_19380_, _19379_, _04060_);
  and (_19381_, _19380_, _19378_);
  and (_19383_, _19381_, _43152_);
  nor (_19384_, \oc8051_golden_model_1.TCON [1], rst);
  nor (_19385_, _19384_, _00000_);
  or (_43420_, _19385_, _19383_);
  not (_19386_, \oc8051_golden_model_1.TCON [2]);
  nor (_19387_, _05447_, _19386_);
  and (_19388_, _05447_, \oc8051_golden_model_1.ACC [2]);
  nor (_19389_, _19388_, _19387_);
  nor (_19390_, _19389_, _04708_);
  nor (_19391_, _04707_, _19386_);
  or (_19393_, _19391_, _19390_);
  and (_19394_, _19393_, _04722_);
  nor (_19395_, _12471_, _09186_);
  nor (_19396_, _19395_, _19387_);
  nor (_19397_, _19396_, _04722_);
  or (_19398_, _19397_, _19394_);
  and (_19399_, _19398_, _03764_);
  nor (_19400_, _06085_, _19386_);
  and (_19401_, _12464_, _06085_);
  nor (_19402_, _19401_, _19400_);
  nor (_19404_, _19402_, _03764_);
  or (_19405_, _19404_, _19399_);
  and (_19406_, _19405_, _04733_);
  and (_19407_, _05447_, _05307_);
  nor (_19408_, _19407_, _19387_);
  nor (_19409_, _19408_, _04733_);
  or (_19410_, _19409_, _19406_);
  and (_19411_, _19410_, _03855_);
  nor (_19412_, _19389_, _03855_);
  or (_19413_, _19412_, _19411_);
  and (_19415_, _19413_, _03760_);
  and (_19416_, _12467_, _06085_);
  nor (_19417_, _19416_, _19400_);
  nor (_19418_, _19417_, _03760_);
  or (_19419_, _19418_, _19415_);
  and (_19420_, _19419_, _03753_);
  and (_19421_, _19401_, _12463_);
  or (_19422_, _19421_, _19400_);
  and (_19423_, _19422_, _03752_);
  or (_19424_, _19423_, _19420_);
  and (_19426_, _19424_, _03747_);
  nor (_19427_, _12514_, _09172_);
  nor (_19428_, _19427_, _19400_);
  nor (_19429_, _19428_, _03747_);
  or (_19430_, _19429_, _07927_);
  or (_19431_, _19430_, _19426_);
  and (_19432_, _06965_, _05447_);
  nor (_19433_, _19387_, _03738_);
  not (_19434_, _19433_);
  nor (_19435_, _19434_, _19432_);
  and (_19437_, _19408_, _08474_);
  or (_19438_, _19437_, _03455_);
  nor (_19439_, _19438_, _19435_);
  and (_19440_, _19439_, _19431_);
  nor (_19441_, _12572_, _09186_);
  nor (_19442_, _19441_, _19387_);
  nor (_19443_, _19442_, _03820_);
  or (_19444_, _19443_, _19440_);
  and (_19445_, _19444_, _04778_);
  and (_19446_, _05447_, _06495_);
  nor (_19448_, _19446_, _19387_);
  nor (_19449_, _19448_, _04778_);
  or (_19450_, _19449_, _19445_);
  nor (_19451_, _19450_, _03897_);
  and (_19452_, _12586_, _05447_);
  or (_19453_, _19387_, _04790_);
  nor (_19454_, _19453_, _19452_);
  or (_19455_, _19454_, _04018_);
  nor (_19456_, _19455_, _19451_);
  and (_19457_, _08748_, _05447_);
  nor (_19459_, _19457_, _19387_);
  nor (_19460_, _19459_, _04792_);
  nor (_19461_, _19460_, _19456_);
  nor (_19462_, _19461_, _03908_);
  nor (_19463_, _19387_, _05765_);
  not (_19464_, _19463_);
  nor (_19465_, _19448_, _03909_);
  and (_19466_, _19465_, _19464_);
  nor (_19467_, _19466_, _19462_);
  nor (_19468_, _19467_, _04027_);
  nor (_19470_, _19389_, _04785_);
  and (_19471_, _19470_, _19464_);
  or (_19472_, _19471_, _19468_);
  and (_19473_, _19472_, _06567_);
  nor (_19474_, _12585_, _09186_);
  nor (_19475_, _19474_, _19387_);
  nor (_19476_, _19475_, _06567_);
  or (_19477_, _19476_, _19473_);
  and (_19478_, _19477_, _06572_);
  nor (_19479_, _08747_, _09186_);
  nor (_19481_, _19479_, _19387_);
  nor (_19482_, _19481_, _06572_);
  or (_19483_, _19482_, _19478_);
  and (_19484_, _19483_, _03774_);
  nor (_19485_, _19396_, _03774_);
  or (_19486_, _19485_, _19484_);
  and (_19487_, _19486_, _03375_);
  nor (_19488_, _19417_, _03375_);
  or (_19489_, _19488_, _19487_);
  and (_19490_, _19489_, _04060_);
  and (_19492_, _12642_, _05447_);
  nor (_19493_, _19492_, _19387_);
  nor (_19494_, _19493_, _04060_);
  or (_19495_, _19494_, _19490_);
  or (_19496_, _19495_, _43156_);
  or (_19497_, _43152_, \oc8051_golden_model_1.TCON [2]);
  and (_19498_, _19497_, _41894_);
  and (_43421_, _19498_, _19496_);
  not (_19499_, \oc8051_golden_model_1.TCON [3]);
  nor (_19500_, _05447_, _19499_);
  and (_19502_, _05447_, \oc8051_golden_model_1.ACC [3]);
  nor (_19503_, _19502_, _19500_);
  nor (_19504_, _19503_, _04708_);
  nor (_19505_, _04707_, _19499_);
  or (_19506_, _19505_, _19504_);
  and (_19507_, _19506_, _04722_);
  nor (_19508_, _12681_, _09186_);
  nor (_19509_, _19508_, _19500_);
  nor (_19510_, _19509_, _04722_);
  or (_19511_, _19510_, _19507_);
  and (_19513_, _19511_, _03764_);
  nor (_19514_, _06085_, _19499_);
  and (_19515_, _12674_, _06085_);
  nor (_19516_, _19515_, _19514_);
  nor (_19517_, _19516_, _03764_);
  or (_19518_, _19517_, _03848_);
  or (_19519_, _19518_, _19513_);
  and (_19520_, _05447_, _05119_);
  nor (_19521_, _19520_, _19500_);
  nand (_19522_, _19521_, _03848_);
  and (_19524_, _19522_, _19519_);
  and (_19525_, _19524_, _03855_);
  nor (_19526_, _19503_, _03855_);
  or (_19527_, _19526_, _19525_);
  and (_19528_, _19527_, _03760_);
  and (_19529_, _12667_, _06085_);
  nor (_19530_, _19529_, _19514_);
  nor (_19531_, _19530_, _03760_);
  or (_19532_, _19531_, _03752_);
  or (_19533_, _19532_, _19528_);
  nor (_19535_, _19514_, _12673_);
  nor (_19536_, _19535_, _19516_);
  or (_19537_, _19536_, _03753_);
  and (_19538_, _19537_, _03747_);
  and (_19539_, _19538_, _19533_);
  nor (_19540_, _12668_, _09172_);
  nor (_19541_, _19540_, _19514_);
  nor (_19542_, _19541_, _03747_);
  or (_19543_, _19542_, _07927_);
  or (_19544_, _19543_, _19539_);
  and (_19546_, _06964_, _05447_);
  nor (_19547_, _19500_, _03738_);
  not (_19548_, _19547_);
  nor (_19549_, _19548_, _19546_);
  and (_19550_, _19521_, _08474_);
  or (_19551_, _19550_, _03455_);
  nor (_19552_, _19551_, _19549_);
  and (_19553_, _19552_, _19544_);
  nor (_19554_, _12775_, _09186_);
  nor (_19555_, _19554_, _19500_);
  nor (_19557_, _19555_, _03820_);
  or (_19558_, _19557_, _19553_);
  and (_19559_, _19558_, _04778_);
  and (_19560_, _05447_, _06345_);
  nor (_19561_, _19560_, _19500_);
  nor (_19562_, _19561_, _04778_);
  or (_19563_, _19562_, _19559_);
  and (_19564_, _19563_, _04790_);
  and (_19565_, _12789_, _05447_);
  nor (_19566_, _19565_, _19500_);
  nor (_19568_, _19566_, _04790_);
  or (_19569_, _19568_, _19564_);
  and (_19570_, _19569_, _04792_);
  and (_19571_, _10491_, _05447_);
  nor (_19572_, _19571_, _19500_);
  nor (_19573_, _19572_, _04792_);
  nor (_19574_, _19573_, _19570_);
  nor (_19575_, _19574_, _03908_);
  nor (_19576_, _19500_, _05622_);
  not (_19577_, _19576_);
  nor (_19579_, _19561_, _03909_);
  and (_19580_, _19579_, _19577_);
  nor (_19581_, _19580_, _19575_);
  nor (_19582_, _19581_, _04027_);
  nor (_19583_, _19503_, _04785_);
  and (_19584_, _19583_, _19577_);
  or (_19585_, _19584_, _19582_);
  and (_19586_, _19585_, _06567_);
  nor (_19587_, _12788_, _09186_);
  nor (_19588_, _19587_, _19500_);
  nor (_19590_, _19588_, _06567_);
  or (_19591_, _19590_, _19586_);
  and (_19592_, _19591_, _06572_);
  nor (_19593_, _08742_, _09186_);
  nor (_19594_, _19593_, _19500_);
  nor (_19595_, _19594_, _06572_);
  or (_19596_, _19595_, _19592_);
  and (_19597_, _19596_, _03774_);
  nor (_19598_, _19509_, _03774_);
  or (_19599_, _19598_, _19597_);
  and (_19601_, _19599_, _03375_);
  nor (_19602_, _19530_, _03375_);
  or (_19603_, _19602_, _19601_);
  and (_19604_, _19603_, _04060_);
  and (_19605_, _12848_, _05447_);
  nor (_19606_, _19605_, _19500_);
  nor (_19607_, _19606_, _04060_);
  or (_19608_, _19607_, _19604_);
  or (_19609_, _19608_, _43156_);
  or (_19610_, _43152_, \oc8051_golden_model_1.TCON [3]);
  and (_19612_, _19610_, _41894_);
  and (_43422_, _19612_, _19609_);
  not (_19613_, \oc8051_golden_model_1.TCON [4]);
  nor (_19614_, _05447_, _19613_);
  and (_19615_, _05447_, \oc8051_golden_model_1.ACC [4]);
  nor (_19616_, _19615_, _19614_);
  nor (_19617_, _19616_, _04708_);
  nor (_19618_, _04707_, _19613_);
  or (_19619_, _19618_, _19617_);
  and (_19620_, _19619_, _04722_);
  nor (_19622_, _12891_, _09186_);
  nor (_19623_, _19622_, _19614_);
  nor (_19624_, _19623_, _04722_);
  or (_19625_, _19624_, _19620_);
  and (_19626_, _19625_, _03764_);
  nor (_19627_, _06085_, _19613_);
  and (_19628_, _12875_, _06085_);
  nor (_19629_, _19628_, _19627_);
  nor (_19630_, _19629_, _03764_);
  or (_19631_, _19630_, _03848_);
  or (_19633_, _19631_, _19626_);
  and (_19634_, _05950_, _05447_);
  nor (_19635_, _19634_, _19614_);
  nand (_19636_, _19635_, _03848_);
  and (_19637_, _19636_, _19633_);
  and (_19638_, _19637_, _03855_);
  nor (_19639_, _19616_, _03855_);
  or (_19640_, _19639_, _19638_);
  and (_19641_, _19640_, _03760_);
  and (_19642_, _12870_, _06085_);
  nor (_19644_, _19642_, _19627_);
  nor (_19645_, _19644_, _03760_);
  or (_19646_, _19645_, _19641_);
  and (_19647_, _19646_, _03753_);
  nor (_19648_, _19627_, _12874_);
  nor (_19649_, _19648_, _19629_);
  and (_19650_, _19649_, _03752_);
  or (_19651_, _19650_, _19647_);
  and (_19652_, _19651_, _03747_);
  nor (_19653_, _12872_, _09172_);
  nor (_19655_, _19653_, _19627_);
  nor (_19656_, _19655_, _03747_);
  or (_19657_, _19656_, _07927_);
  or (_19658_, _19657_, _19652_);
  and (_19659_, _06969_, _05447_);
  nor (_19660_, _19614_, _03738_);
  not (_19661_, _19660_);
  nor (_19662_, _19661_, _19659_);
  and (_19663_, _19635_, _08474_);
  or (_19664_, _19663_, _03455_);
  nor (_19666_, _19664_, _19662_);
  and (_19667_, _19666_, _19658_);
  nor (_19668_, _12982_, _09186_);
  nor (_19669_, _19668_, _19614_);
  nor (_19670_, _19669_, _03820_);
  or (_19671_, _19670_, _19667_);
  and (_19672_, _19671_, _04778_);
  and (_19673_, _06456_, _05447_);
  nor (_19674_, _19673_, _19614_);
  nor (_19675_, _19674_, _04778_);
  or (_19677_, _19675_, _19672_);
  and (_19678_, _19677_, _04790_);
  and (_19679_, _12997_, _05447_);
  nor (_19680_, _19679_, _19614_);
  nor (_19681_, _19680_, _04790_);
  or (_19682_, _19681_, _19678_);
  and (_19683_, _19682_, _04792_);
  and (_19684_, _08741_, _05447_);
  nor (_19685_, _19684_, _19614_);
  nor (_19686_, _19685_, _04792_);
  nor (_19688_, _19686_, _19683_);
  nor (_19689_, _19688_, _03908_);
  nor (_19690_, _19614_, _08336_);
  not (_19691_, _19690_);
  nor (_19692_, _19674_, _03909_);
  and (_19693_, _19692_, _19691_);
  nor (_19694_, _19693_, _19689_);
  nor (_19695_, _19694_, _04027_);
  nor (_19696_, _19616_, _04785_);
  and (_19697_, _19696_, _19691_);
  or (_19699_, _19697_, _19695_);
  and (_19700_, _19699_, _06567_);
  nor (_19701_, _12996_, _09186_);
  nor (_19702_, _19701_, _19614_);
  nor (_19703_, _19702_, _06567_);
  or (_19704_, _19703_, _19700_);
  and (_19705_, _19704_, _06572_);
  nor (_19706_, _08740_, _09186_);
  nor (_19707_, _19706_, _19614_);
  nor (_19708_, _19707_, _06572_);
  or (_19710_, _19708_, _19705_);
  and (_19711_, _19710_, _03774_);
  nor (_19712_, _19623_, _03774_);
  or (_19713_, _19712_, _19711_);
  and (_19714_, _19713_, _03375_);
  nor (_19715_, _19644_, _03375_);
  or (_19716_, _19715_, _19714_);
  and (_19717_, _19716_, _04060_);
  and (_19718_, _13056_, _05447_);
  nor (_19719_, _19718_, _19614_);
  nor (_19721_, _19719_, _04060_);
  or (_19722_, _19721_, _19717_);
  or (_19723_, _19722_, _43156_);
  or (_19724_, _43152_, \oc8051_golden_model_1.TCON [4]);
  and (_19725_, _19724_, _41894_);
  and (_43423_, _19725_, _19723_);
  not (_19726_, \oc8051_golden_model_1.TCON [5]);
  nor (_19727_, _05447_, _19726_);
  and (_19728_, _05447_, \oc8051_golden_model_1.ACC [5]);
  nor (_19729_, _19728_, _19727_);
  nor (_19731_, _19729_, _04708_);
  nor (_19732_, _04707_, _19726_);
  or (_19733_, _19732_, _19731_);
  and (_19734_, _19733_, _04722_);
  nor (_19735_, _13090_, _09186_);
  nor (_19736_, _19735_, _19727_);
  nor (_19737_, _19736_, _04722_);
  or (_19738_, _19737_, _19734_);
  and (_19739_, _19738_, _03764_);
  nor (_19740_, _06085_, _19726_);
  and (_19742_, _13094_, _06085_);
  nor (_19743_, _19742_, _19740_);
  nor (_19744_, _19743_, _03764_);
  or (_19745_, _19744_, _03848_);
  or (_19746_, _19745_, _19739_);
  and (_19747_, _05857_, _05447_);
  nor (_19748_, _19747_, _19727_);
  nand (_19749_, _19748_, _03848_);
  and (_19750_, _19749_, _19746_);
  and (_19751_, _19750_, _03855_);
  nor (_19753_, _19729_, _03855_);
  or (_19754_, _19753_, _19751_);
  and (_19755_, _19754_, _03760_);
  and (_19756_, _13071_, _06085_);
  nor (_19757_, _19756_, _19740_);
  nor (_19758_, _19757_, _03760_);
  or (_19759_, _19758_, _03752_);
  or (_19760_, _19759_, _19755_);
  nor (_19761_, _19740_, _13109_);
  nor (_19762_, _19761_, _19743_);
  or (_19764_, _19762_, _03753_);
  and (_19765_, _19764_, _03747_);
  and (_19766_, _19765_, _19760_);
  nor (_19767_, _13073_, _09172_);
  nor (_19768_, _19767_, _19740_);
  nor (_19769_, _19768_, _03747_);
  or (_19770_, _19769_, _07927_);
  or (_19771_, _19770_, _19766_);
  and (_19772_, _06968_, _05447_);
  nor (_19773_, _19727_, _03738_);
  not (_19775_, _19773_);
  nor (_19776_, _19775_, _19772_);
  and (_19777_, _19748_, _08474_);
  or (_19778_, _19777_, _03455_);
  nor (_19779_, _19778_, _19776_);
  and (_19780_, _19779_, _19771_);
  nor (_19781_, _13182_, _09186_);
  nor (_19782_, _19781_, _19727_);
  nor (_19783_, _19782_, _03820_);
  or (_19784_, _19783_, _19780_);
  and (_19786_, _19784_, _04778_);
  and (_19787_, _06447_, _05447_);
  nor (_19788_, _19787_, _19727_);
  nor (_19789_, _19788_, _04778_);
  or (_19790_, _19789_, _19786_);
  nor (_19791_, _19790_, _03897_);
  and (_19792_, _13196_, _05447_);
  or (_19793_, _19727_, _04790_);
  nor (_19794_, _19793_, _19792_);
  or (_19795_, _19794_, _04018_);
  nor (_19797_, _19795_, _19791_);
  and (_19798_, _10493_, _05447_);
  nor (_19799_, _19798_, _19727_);
  nor (_19800_, _19799_, _04792_);
  nor (_19801_, _19800_, _19797_);
  nor (_19802_, _19801_, _03908_);
  nor (_19803_, _19727_, _08335_);
  not (_19804_, _19803_);
  nor (_19805_, _19788_, _03909_);
  and (_19806_, _19805_, _19804_);
  nor (_19808_, _19806_, _19802_);
  nor (_19809_, _19808_, _04027_);
  nor (_19810_, _19729_, _04785_);
  and (_19811_, _19810_, _19804_);
  or (_19812_, _19811_, _19809_);
  and (_19813_, _19812_, _06567_);
  nor (_19814_, _13195_, _09186_);
  nor (_19815_, _19814_, _19727_);
  nor (_19816_, _19815_, _06567_);
  or (_19817_, _19816_, _19813_);
  and (_19819_, _19817_, _06572_);
  nor (_19820_, _08738_, _09186_);
  nor (_19821_, _19820_, _19727_);
  nor (_19822_, _19821_, _06572_);
  or (_19823_, _19822_, _19819_);
  and (_19824_, _19823_, _03774_);
  nor (_19825_, _19736_, _03774_);
  or (_19826_, _19825_, _19824_);
  and (_19827_, _19826_, _03375_);
  nor (_19828_, _19757_, _03375_);
  or (_19830_, _19828_, _19827_);
  and (_19831_, _19830_, _04060_);
  and (_19832_, _13255_, _05447_);
  nor (_19833_, _19832_, _19727_);
  nor (_19834_, _19833_, _04060_);
  or (_19835_, _19834_, _19831_);
  or (_19836_, _19835_, _43156_);
  or (_19837_, _43152_, \oc8051_golden_model_1.TCON [5]);
  and (_19838_, _19837_, _41894_);
  and (_43424_, _19838_, _19836_);
  not (_19840_, \oc8051_golden_model_1.TCON [6]);
  nor (_19841_, _05447_, _19840_);
  and (_19842_, _05447_, \oc8051_golden_model_1.ACC [6]);
  nor (_19843_, _19842_, _19841_);
  nor (_19844_, _19843_, _04708_);
  nor (_19845_, _04707_, _19840_);
  or (_19846_, _19845_, _19844_);
  and (_19847_, _19846_, _04722_);
  nor (_19848_, _13293_, _09186_);
  nor (_19849_, _19848_, _19841_);
  nor (_19851_, _19849_, _04722_);
  or (_19852_, _19851_, _19847_);
  and (_19853_, _19852_, _03764_);
  nor (_19854_, _06085_, _19840_);
  and (_19855_, _13297_, _06085_);
  nor (_19856_, _19855_, _19854_);
  nor (_19857_, _19856_, _03764_);
  or (_19858_, _19857_, _03848_);
  or (_19859_, _19858_, _19853_);
  and (_19860_, _06065_, _05447_);
  nor (_19862_, _19860_, _19841_);
  nand (_19863_, _19862_, _03848_);
  and (_19864_, _19863_, _19859_);
  and (_19865_, _19864_, _03855_);
  nor (_19866_, _19843_, _03855_);
  or (_19867_, _19866_, _19865_);
  and (_19868_, _19867_, _03760_);
  and (_19869_, _13277_, _06085_);
  nor (_19870_, _19869_, _19854_);
  nor (_19871_, _19870_, _03760_);
  or (_19873_, _19871_, _03752_);
  or (_19874_, _19873_, _19868_);
  nor (_19875_, _19854_, _13312_);
  nor (_19876_, _19875_, _19856_);
  or (_19877_, _19876_, _03753_);
  and (_19878_, _19877_, _03747_);
  and (_19879_, _19878_, _19874_);
  nor (_19880_, _13279_, _09172_);
  nor (_19881_, _19880_, _19854_);
  nor (_19882_, _19881_, _03747_);
  or (_19884_, _19882_, _07927_);
  or (_19885_, _19884_, _19879_);
  and (_19886_, _06641_, _05447_);
  nor (_19887_, _19841_, _03738_);
  not (_19888_, _19887_);
  nor (_19889_, _19888_, _19886_);
  and (_19890_, _19862_, _08474_);
  or (_19891_, _19890_, _03455_);
  nor (_19892_, _19891_, _19889_);
  and (_19893_, _19892_, _19885_);
  nor (_19895_, _13387_, _09186_);
  nor (_19896_, _19895_, _19841_);
  nor (_19897_, _19896_, _03820_);
  or (_19898_, _19897_, _19893_);
  and (_19899_, _19898_, _04778_);
  and (_19900_, _13394_, _05447_);
  nor (_19901_, _19900_, _19841_);
  nor (_19902_, _19901_, _04778_);
  or (_19903_, _19902_, _19899_);
  and (_19904_, _19903_, _04790_);
  and (_19906_, _13402_, _05447_);
  nor (_19907_, _19906_, _19841_);
  nor (_19908_, _19907_, _04790_);
  or (_19909_, _19908_, _19904_);
  and (_19910_, _19909_, _04792_);
  and (_19911_, _08736_, _05447_);
  nor (_19912_, _19911_, _19841_);
  nor (_19913_, _19912_, _04792_);
  nor (_19914_, _19913_, _19910_);
  nor (_19915_, _19914_, _03908_);
  nor (_19917_, _19841_, _08322_);
  not (_19918_, _19917_);
  nor (_19919_, _19901_, _03909_);
  and (_19920_, _19919_, _19918_);
  nor (_19921_, _19920_, _19915_);
  nor (_19922_, _19921_, _04027_);
  nor (_19923_, _19843_, _04785_);
  and (_19924_, _19923_, _19918_);
  nor (_19925_, _19924_, _03914_);
  not (_19926_, _19925_);
  nor (_19928_, _19926_, _19922_);
  nor (_19929_, _13401_, _09186_);
  or (_19930_, _19841_, _06567_);
  nor (_19931_, _19930_, _19929_);
  or (_19932_, _19931_, _04011_);
  nor (_19933_, _19932_, _19928_);
  nor (_19934_, _08735_, _09186_);
  nor (_19935_, _19934_, _19841_);
  nor (_19936_, _19935_, _06572_);
  or (_19937_, _19936_, _19933_);
  and (_19939_, _19937_, _03774_);
  nor (_19940_, _19849_, _03774_);
  or (_19941_, _19940_, _19939_);
  and (_19942_, _19941_, _03375_);
  nor (_19943_, _19870_, _03375_);
  or (_19944_, _19943_, _19942_);
  and (_19945_, _19944_, _04060_);
  nor (_19946_, _13460_, _09186_);
  nor (_19947_, _19946_, _19841_);
  nor (_19948_, _19947_, _04060_);
  or (_19950_, _19948_, _19945_);
  or (_19951_, _19950_, _43156_);
  or (_19952_, _43152_, \oc8051_golden_model_1.TCON [6]);
  and (_19953_, _19952_, _41894_);
  and (_43425_, _19953_, _19951_);
  not (_19954_, \oc8051_golden_model_1.TL0 [0]);
  nor (_19955_, _05589_, _19954_);
  and (_19956_, _05716_, _05589_);
  nor (_19957_, _19956_, _19955_);
  and (_19958_, _19957_, _17157_);
  nand (_19960_, _08753_, _05589_);
  nor (_19961_, _19955_, _04785_);
  and (_19962_, _19961_, _19960_);
  nor (_19963_, _19955_, _03738_);
  or (_19964_, _06733_, _09271_);
  and (_19965_, _19964_, _19963_);
  and (_19966_, _05589_, _04700_);
  nor (_19967_, _19966_, _19955_);
  and (_19968_, _19967_, _08474_);
  and (_19969_, _05589_, \oc8051_golden_model_1.ACC [0]);
  nor (_19971_, _19969_, _19955_);
  nor (_19972_, _19971_, _04708_);
  nor (_19973_, _04707_, _19954_);
  or (_19974_, _19973_, _19972_);
  and (_19975_, _19974_, _04722_);
  nor (_19976_, _19957_, _04722_);
  or (_19977_, _19976_, _19975_);
  and (_19978_, _19977_, _04733_);
  nor (_19979_, _19967_, _04733_);
  nor (_19980_, _19979_, _19978_);
  nor (_19982_, _19980_, _03854_);
  nor (_19983_, _19971_, _03855_);
  or (_19984_, _19983_, _07927_);
  nor (_19985_, _19984_, _19982_);
  nor (_19986_, _19985_, _19968_);
  not (_19987_, _19986_);
  nor (_19988_, _19987_, _19965_);
  and (_19989_, _19988_, _03820_);
  not (_19990_, _05480_);
  nor (_19991_, _12164_, _19990_);
  nor (_19993_, _19991_, _19955_);
  nor (_19994_, _19993_, _03820_);
  or (_19995_, _19994_, _19989_);
  and (_19996_, _19995_, _04778_);
  and (_19997_, _05589_, _06479_);
  nor (_19998_, _19997_, _19955_);
  nor (_19999_, _19998_, _04778_);
  or (_20000_, _19999_, _19996_);
  and (_20001_, _20000_, _04790_);
  and (_20002_, _12178_, _05480_);
  nor (_20004_, _20002_, _19955_);
  nor (_20005_, _20004_, _04790_);
  or (_20006_, _20005_, _20001_);
  and (_20007_, _20006_, _04792_);
  nor (_20008_, _10488_, _09271_);
  nor (_20009_, _20008_, _19955_);
  nand (_20010_, _19960_, _04018_);
  nor (_20011_, _20010_, _20009_);
  nor (_20012_, _20011_, _20007_);
  nor (_20013_, _20012_, _03908_);
  nor (_20015_, _19998_, _03909_);
  not (_20016_, _20015_);
  nor (_20017_, _20016_, _19956_);
  nor (_20018_, _20017_, _04027_);
  not (_20019_, _20018_);
  nor (_20020_, _20019_, _20013_);
  nor (_20021_, _20020_, _19962_);
  and (_20022_, _20021_, _06567_);
  nor (_20023_, _12177_, _19990_);
  nor (_20024_, _20023_, _19955_);
  nor (_20026_, _20024_, _06567_);
  or (_20027_, _20026_, _20022_);
  and (_20028_, _20027_, _06572_);
  nor (_20029_, _20009_, _06572_);
  nor (_20030_, _20029_, _17157_);
  not (_20031_, _20030_);
  nor (_20032_, _20031_, _20028_);
  nor (_20033_, _20032_, _19958_);
  or (_20034_, _20033_, _43156_);
  or (_20035_, _43152_, \oc8051_golden_model_1.TL0 [0]);
  and (_20037_, _20035_, _41894_);
  and (_43428_, _20037_, _20034_);
  nor (_20038_, _05589_, \oc8051_golden_model_1.TL0 [1]);
  nor (_20039_, _20038_, _04778_);
  and (_20040_, _05589_, _04595_);
  not (_20041_, _20040_);
  and (_20042_, _20041_, _20039_);
  not (_20043_, \oc8051_golden_model_1.TL0 [1]);
  nor (_20044_, _05589_, _20043_);
  nor (_20045_, _20044_, _03738_);
  or (_20047_, _06688_, _09271_);
  and (_20048_, _20047_, _20045_);
  not (_20049_, _20048_);
  and (_20050_, _05480_, \oc8051_golden_model_1.ACC [1]);
  nor (_20051_, _20050_, _20044_);
  nor (_20052_, _20051_, _04708_);
  nor (_20053_, _04707_, _20043_);
  or (_20054_, _20053_, _20052_);
  and (_20055_, _20054_, _04722_);
  and (_20056_, _12262_, _05480_);
  nor (_20058_, _20056_, _20038_);
  and (_20059_, _20058_, _03850_);
  or (_20060_, _20059_, _20055_);
  and (_20061_, _20060_, _04733_);
  and (_20062_, _05589_, _04900_);
  nor (_20063_, _20062_, _20044_);
  nor (_20064_, _20063_, _04733_);
  nor (_20065_, _20064_, _20061_);
  nor (_20066_, _20065_, _03854_);
  nor (_20067_, _20051_, _03855_);
  or (_20069_, _20067_, _07927_);
  or (_20070_, _20069_, _20066_);
  and (_20071_, _20063_, _08474_);
  nor (_20072_, _20071_, _03455_);
  and (_20073_, _20072_, _20070_);
  and (_20074_, _20073_, _20049_);
  nor (_20075_, _12352_, _19990_);
  nor (_20076_, _20075_, _20044_);
  nor (_20077_, _20076_, _03820_);
  nor (_20078_, _20077_, _20074_);
  nor (_20080_, _20078_, _03903_);
  nor (_20081_, _20080_, _20042_);
  nor (_20082_, _20081_, _03897_);
  and (_20083_, _12366_, _05480_);
  or (_20084_, _20083_, _20044_);
  and (_20085_, _20084_, _03897_);
  nor (_20086_, _20085_, _20082_);
  nor (_20087_, _20086_, _04018_);
  nor (_20088_, _08751_, _09271_);
  nor (_20089_, _20088_, _20044_);
  and (_20091_, _20050_, _08366_);
  nor (_20092_, _20091_, _20089_);
  and (_20093_, _20092_, _04018_);
  or (_20094_, _20093_, _20087_);
  and (_20095_, _20094_, _03909_);
  and (_20096_, _12244_, _05480_);
  or (_20097_, _20096_, _20044_);
  and (_20098_, _20097_, _03908_);
  or (_20099_, _20098_, _20095_);
  and (_20100_, _20099_, _04785_);
  nor (_20102_, _20091_, _20044_);
  nor (_20103_, _20102_, _04785_);
  or (_20104_, _20103_, _20100_);
  and (_20105_, _20104_, _06567_);
  nor (_20106_, _12365_, _19990_);
  or (_20107_, _20106_, _20044_);
  and (_20108_, _20107_, _03914_);
  or (_20109_, _20108_, _20105_);
  and (_20110_, _20109_, _06572_);
  nor (_20111_, _20089_, _06572_);
  or (_20113_, _20111_, _20110_);
  nor (_20114_, _20113_, _03773_);
  nor (_20115_, _20058_, _03774_);
  or (_20116_, _20115_, _03772_);
  nor (_20117_, _20116_, _20114_);
  nor (_20118_, _20056_, _20044_);
  nor (_20119_, _20118_, _04060_);
  or (_20120_, _20119_, _20117_);
  or (_20121_, _20120_, _43156_);
  or (_20122_, _43152_, \oc8051_golden_model_1.TL0 [1]);
  and (_20124_, _20122_, _41894_);
  and (_43429_, _20124_, _20121_);
  not (_20125_, \oc8051_golden_model_1.TL0 [2]);
  nor (_20126_, _05589_, _20125_);
  nor (_20127_, _20126_, _03738_);
  or (_20128_, _06824_, _09271_);
  and (_20129_, _20128_, _20127_);
  not (_20130_, _20129_);
  and (_20131_, _05589_, _05307_);
  nor (_20132_, _20131_, _20126_);
  and (_20134_, _20132_, _08474_);
  and (_20135_, _05589_, \oc8051_golden_model_1.ACC [2]);
  nor (_20136_, _20135_, _20126_);
  nor (_20137_, _20136_, _04708_);
  nor (_20138_, _04707_, _20125_);
  or (_20139_, _20138_, _20137_);
  and (_20140_, _20139_, _04722_);
  nor (_20141_, _12471_, _09271_);
  nor (_20142_, _20141_, _20126_);
  nor (_20143_, _20142_, _04722_);
  or (_20145_, _20143_, _20140_);
  and (_20146_, _20145_, _04733_);
  nor (_20147_, _20132_, _04733_);
  nor (_20148_, _20147_, _20146_);
  nor (_20149_, _20148_, _03854_);
  nor (_20150_, _20136_, _03855_);
  or (_20151_, _20150_, _07927_);
  nor (_20152_, _20151_, _20149_);
  nor (_20153_, _20152_, _20134_);
  and (_20154_, _20153_, _20130_);
  and (_20156_, _20154_, _03820_);
  nor (_20157_, _12572_, _19990_);
  nor (_20158_, _20157_, _20126_);
  nor (_20159_, _20158_, _03820_);
  or (_20160_, _20159_, _20156_);
  and (_20161_, _20160_, _04778_);
  and (_20162_, _05589_, _06495_);
  nor (_20163_, _20162_, _20126_);
  nor (_20164_, _20163_, _04778_);
  or (_20165_, _20164_, _20161_);
  and (_20167_, _20165_, _04790_);
  and (_20168_, _12586_, _05480_);
  nor (_20169_, _20168_, _20126_);
  nor (_20170_, _20169_, _04790_);
  or (_20171_, _20170_, _20167_);
  and (_20172_, _20171_, _04792_);
  and (_20173_, _08748_, _05480_);
  nor (_20174_, _20173_, _20126_);
  nor (_20175_, _20174_, _04792_);
  nor (_20176_, _20175_, _20172_);
  nor (_20178_, _20176_, _03908_);
  nor (_20179_, _20126_, _05765_);
  not (_20180_, _20179_);
  nor (_20181_, _20163_, _03909_);
  and (_20182_, _20181_, _20180_);
  nor (_20183_, _20182_, _20178_);
  nor (_20184_, _20183_, _04027_);
  nor (_20185_, _20136_, _04785_);
  and (_20186_, _20185_, _20180_);
  nor (_20187_, _20186_, _03914_);
  not (_20189_, _20187_);
  nor (_20190_, _20189_, _20184_);
  or (_20191_, _12585_, _09271_);
  nor (_20192_, _20126_, _06567_);
  and (_20193_, _20192_, _20191_);
  or (_20194_, _20193_, _04011_);
  nor (_20195_, _20194_, _20190_);
  nor (_20196_, _08747_, _09271_);
  nor (_20197_, _20196_, _20126_);
  nor (_20198_, _20197_, _06572_);
  or (_20200_, _20198_, _03773_);
  nor (_20201_, _20200_, _20195_);
  and (_20202_, _20142_, _03773_);
  or (_20203_, _20202_, _03772_);
  nor (_20204_, _20203_, _20201_);
  and (_20205_, _12642_, _05480_);
  nor (_20206_, _20205_, _20126_);
  nor (_20207_, _20206_, _04060_);
  or (_20208_, _20207_, _20204_);
  or (_20209_, _20208_, _43156_);
  or (_20211_, _43152_, \oc8051_golden_model_1.TL0 [2]);
  and (_20212_, _20211_, _41894_);
  and (_43430_, _20212_, _20209_);
  not (_20213_, \oc8051_golden_model_1.TL0 [3]);
  nor (_20214_, _05589_, _20213_);
  and (_20215_, _05589_, \oc8051_golden_model_1.ACC [3]);
  nor (_20216_, _20215_, _20214_);
  nor (_20217_, _20216_, _04708_);
  nor (_20218_, _04707_, _20213_);
  or (_20219_, _20218_, _20217_);
  and (_20221_, _20219_, _04722_);
  nor (_20222_, _12681_, _09271_);
  nor (_20223_, _20222_, _20214_);
  nor (_20224_, _20223_, _04722_);
  or (_20225_, _20224_, _20221_);
  and (_20226_, _20225_, _04733_);
  and (_20227_, _05589_, _05119_);
  nor (_20228_, _20227_, _20214_);
  nor (_20229_, _20228_, _04733_);
  nor (_20230_, _20229_, _20226_);
  nor (_20232_, _20230_, _03854_);
  nor (_20233_, _20216_, _03855_);
  or (_20234_, _20233_, _07927_);
  or (_20235_, _20234_, _20232_);
  nor (_20236_, _20214_, _03738_);
  or (_20237_, _06779_, _09271_);
  and (_20238_, _20237_, _20236_);
  and (_20239_, _20228_, _08474_);
  or (_20240_, _20239_, _03455_);
  nor (_20241_, _20240_, _20238_);
  and (_20243_, _20241_, _20235_);
  nor (_20244_, _12775_, _09271_);
  nor (_20245_, _20244_, _20214_);
  nor (_20246_, _20245_, _03820_);
  or (_20247_, _20246_, _20243_);
  and (_20248_, _20247_, _04778_);
  and (_20249_, _05589_, _06345_);
  nor (_20250_, _20249_, _20214_);
  nor (_20251_, _20250_, _04778_);
  or (_20252_, _20251_, _20248_);
  nor (_20254_, _20252_, _03897_);
  nand (_20255_, _12789_, _05589_);
  nor (_20256_, _20214_, _04790_);
  and (_20257_, _20256_, _20255_);
  or (_20258_, _20257_, _04018_);
  nor (_20259_, _20258_, _20254_);
  and (_20260_, _10491_, _05480_);
  nor (_20261_, _20260_, _20214_);
  nor (_20262_, _20261_, _04792_);
  nor (_20263_, _20262_, _20259_);
  nor (_20265_, _20263_, _03908_);
  nor (_20266_, _20214_, _05622_);
  not (_20267_, _20266_);
  nor (_20268_, _20250_, _03909_);
  and (_20269_, _20268_, _20267_);
  nor (_20270_, _20269_, _20265_);
  nor (_20271_, _20270_, _04027_);
  nor (_20272_, _20216_, _04785_);
  and (_20273_, _20272_, _20267_);
  or (_20274_, _20273_, _20271_);
  and (_20276_, _20274_, _06567_);
  nor (_20277_, _12788_, _19990_);
  nor (_20278_, _20277_, _20214_);
  nor (_20279_, _20278_, _06567_);
  or (_20280_, _20279_, _20276_);
  and (_20281_, _20280_, _06572_);
  nor (_20282_, _08742_, _09271_);
  nor (_20283_, _20282_, _20214_);
  nor (_20284_, _20283_, _06572_);
  or (_20285_, _20284_, _03773_);
  nor (_20287_, _20285_, _20281_);
  and (_20288_, _20223_, _03773_);
  or (_20289_, _20288_, _03772_);
  nor (_20290_, _20289_, _20287_);
  and (_20291_, _12848_, _05480_);
  nor (_20292_, _20291_, _20214_);
  nor (_20293_, _20292_, _04060_);
  or (_20294_, _20293_, _20290_);
  or (_20295_, _20294_, _43156_);
  or (_20296_, _43152_, \oc8051_golden_model_1.TL0 [3]);
  and (_20298_, _20296_, _41894_);
  and (_43431_, _20298_, _20295_);
  not (_20299_, \oc8051_golden_model_1.TL0 [4]);
  nor (_20300_, _05589_, _20299_);
  and (_20301_, _05589_, \oc8051_golden_model_1.ACC [4]);
  nor (_20302_, _20301_, _20300_);
  nor (_20303_, _20302_, _04708_);
  nor (_20304_, _04707_, _20299_);
  or (_20305_, _20304_, _20303_);
  and (_20306_, _20305_, _04722_);
  nor (_20308_, _12891_, _09271_);
  nor (_20309_, _20308_, _20300_);
  nor (_20310_, _20309_, _04722_);
  or (_20311_, _20310_, _20306_);
  and (_20312_, _20311_, _04733_);
  and (_20313_, _05950_, _05589_);
  nor (_20314_, _20313_, _20300_);
  nor (_20315_, _20314_, _04733_);
  nor (_20316_, _20315_, _20312_);
  nor (_20317_, _20316_, _03854_);
  nor (_20319_, _20302_, _03855_);
  or (_20320_, _20319_, _07927_);
  nor (_20321_, _20320_, _20317_);
  nor (_20322_, _20300_, _03738_);
  or (_20323_, _06918_, _09271_);
  and (_20324_, _20323_, _20322_);
  and (_20325_, _20314_, _08474_);
  or (_20326_, _20325_, _03455_);
  or (_20327_, _20326_, _20324_);
  nor (_20328_, _20327_, _20321_);
  nor (_20330_, _12982_, _09271_);
  nor (_20331_, _20330_, _20300_);
  nor (_20332_, _20331_, _03820_);
  or (_20333_, _20332_, _20328_);
  and (_20334_, _20333_, _04778_);
  and (_20335_, _06456_, _05589_);
  nor (_20336_, _20335_, _20300_);
  nor (_20337_, _20336_, _04778_);
  or (_20338_, _20337_, _20334_);
  and (_20339_, _20338_, _04790_);
  and (_20341_, _12997_, _05480_);
  nor (_20342_, _20341_, _20300_);
  nor (_20343_, _20342_, _04790_);
  or (_20344_, _20343_, _20339_);
  and (_20345_, _20344_, _04792_);
  and (_20346_, _08741_, _05480_);
  nor (_20347_, _20346_, _20300_);
  nor (_20348_, _20347_, _04792_);
  nor (_20349_, _20348_, _20345_);
  nor (_20350_, _20349_, _03908_);
  nor (_20352_, _20300_, _08336_);
  not (_20353_, _20352_);
  nor (_20354_, _20336_, _03909_);
  and (_20355_, _20354_, _20353_);
  nor (_20356_, _20355_, _20350_);
  nor (_20357_, _20356_, _04027_);
  nor (_20358_, _20302_, _04785_);
  and (_20359_, _20358_, _20353_);
  nor (_20360_, _20359_, _03914_);
  not (_20361_, _20360_);
  nor (_20363_, _20361_, _20357_);
  or (_20364_, _12996_, _09271_);
  nor (_20365_, _20300_, _06567_);
  and (_20366_, _20365_, _20364_);
  or (_20367_, _20366_, _04011_);
  nor (_20368_, _20367_, _20363_);
  nor (_20369_, _08740_, _09271_);
  nor (_20370_, _20369_, _20300_);
  nor (_20371_, _20370_, _06572_);
  or (_20372_, _20371_, _03773_);
  nor (_20374_, _20372_, _20368_);
  and (_20375_, _20309_, _03773_);
  or (_20376_, _20375_, _03772_);
  nor (_20377_, _20376_, _20374_);
  and (_20378_, _13056_, _05480_);
  nor (_20379_, _20378_, _20300_);
  nor (_20380_, _20379_, _04060_);
  or (_20381_, _20380_, _20377_);
  or (_20382_, _20381_, _43156_);
  or (_20383_, _43152_, \oc8051_golden_model_1.TL0 [4]);
  and (_20385_, _20383_, _41894_);
  and (_43432_, _20385_, _20382_);
  not (_20386_, \oc8051_golden_model_1.TL0 [5]);
  nor (_20387_, _05589_, _20386_);
  and (_20388_, _05589_, \oc8051_golden_model_1.ACC [5]);
  nor (_20389_, _20388_, _20387_);
  nor (_20390_, _20389_, _04708_);
  nor (_20391_, _04707_, _20386_);
  or (_20392_, _20391_, _20390_);
  and (_20393_, _20392_, _04722_);
  nor (_20395_, _13090_, _09271_);
  nor (_20396_, _20395_, _20387_);
  nor (_20397_, _20396_, _04722_);
  or (_20398_, _20397_, _20393_);
  and (_20399_, _20398_, _04733_);
  and (_20400_, _05857_, _05589_);
  nor (_20401_, _20400_, _20387_);
  nor (_20402_, _20401_, _04733_);
  nor (_20403_, _20402_, _20399_);
  nor (_20404_, _20403_, _03854_);
  nor (_20406_, _20389_, _03855_);
  or (_20407_, _20406_, _07927_);
  or (_20408_, _20407_, _20404_);
  nor (_20409_, _20387_, _03738_);
  or (_20410_, _06873_, _09271_);
  and (_20411_, _20410_, _20409_);
  and (_20412_, _20401_, _08474_);
  or (_20413_, _20412_, _03455_);
  nor (_20414_, _20413_, _20411_);
  and (_20415_, _20414_, _20408_);
  nor (_20417_, _13182_, _09271_);
  nor (_20418_, _20417_, _20387_);
  nor (_20419_, _20418_, _03820_);
  or (_20420_, _20419_, _20415_);
  and (_20421_, _20420_, _04778_);
  and (_20422_, _06447_, _05589_);
  nor (_20423_, _20422_, _20387_);
  nor (_20424_, _20423_, _04778_);
  or (_20425_, _20424_, _20421_);
  nor (_20426_, _20425_, _03897_);
  nand (_20428_, _13196_, _05589_);
  nor (_20429_, _20387_, _04790_);
  and (_20430_, _20429_, _20428_);
  or (_20431_, _20430_, _04018_);
  nor (_20432_, _20431_, _20426_);
  and (_20433_, _10493_, _05480_);
  nor (_20434_, _20433_, _20387_);
  nor (_20435_, _20434_, _04792_);
  nor (_20436_, _20435_, _20432_);
  nor (_20437_, _20436_, _03908_);
  nor (_20439_, _20387_, _08335_);
  not (_20440_, _20439_);
  nor (_20441_, _20423_, _03909_);
  and (_20442_, _20441_, _20440_);
  nor (_20443_, _20442_, _20437_);
  nor (_20444_, _20443_, _04027_);
  nor (_20445_, _20389_, _04785_);
  and (_20446_, _20445_, _20440_);
  or (_20447_, _20446_, _20444_);
  and (_20448_, _20447_, _06567_);
  nor (_20450_, _13195_, _19990_);
  nor (_20451_, _20450_, _20387_);
  nor (_20452_, _20451_, _06567_);
  or (_20453_, _20452_, _20448_);
  and (_20454_, _20453_, _06572_);
  nor (_20455_, _08738_, _09271_);
  nor (_20456_, _20455_, _20387_);
  nor (_20457_, _20456_, _06572_);
  nor (_20458_, _20457_, _20454_);
  nor (_20459_, _20458_, _03773_);
  nor (_20461_, _20396_, _03774_);
  or (_20462_, _20461_, _03772_);
  nor (_20463_, _20462_, _20459_);
  and (_20464_, _13255_, _05480_);
  nor (_20465_, _20464_, _20387_);
  and (_20466_, _20465_, _03772_);
  nor (_20467_, _20466_, _20463_);
  or (_20468_, _20467_, _43156_);
  or (_20469_, _43152_, \oc8051_golden_model_1.TL0 [5]);
  and (_20470_, _20469_, _41894_);
  and (_43435_, _20470_, _20468_);
  not (_20472_, \oc8051_golden_model_1.TL0 [6]);
  nor (_20473_, _05589_, _20472_);
  and (_20474_, _05589_, \oc8051_golden_model_1.ACC [6]);
  nor (_20475_, _20474_, _20473_);
  nor (_20476_, _20475_, _04708_);
  nor (_20477_, _04707_, _20472_);
  or (_20478_, _20477_, _20476_);
  and (_20479_, _20478_, _04722_);
  nor (_20480_, _13293_, _09271_);
  nor (_20482_, _20480_, _20473_);
  nor (_20483_, _20482_, _04722_);
  or (_20484_, _20483_, _20479_);
  and (_20485_, _20484_, _04733_);
  and (_20486_, _06065_, _05589_);
  nor (_20487_, _20486_, _20473_);
  nor (_20488_, _20487_, _04733_);
  nor (_20489_, _20488_, _20485_);
  nor (_20490_, _20489_, _03854_);
  nor (_20491_, _20475_, _03855_);
  or (_20493_, _20491_, _07927_);
  nor (_20494_, _20493_, _20490_);
  nor (_20495_, _20473_, _03738_);
  nand (_20496_, _06641_, _05589_);
  and (_20497_, _20496_, _20495_);
  and (_20498_, _20487_, _08474_);
  or (_20499_, _20498_, _03455_);
  or (_20500_, _20499_, _20497_);
  nor (_20501_, _20500_, _20494_);
  nor (_20502_, _13387_, _09271_);
  nor (_20504_, _20502_, _20473_);
  nor (_20505_, _20504_, _03820_);
  or (_20506_, _20505_, _20501_);
  and (_20507_, _20506_, _04778_);
  and (_20508_, _13394_, _05589_);
  nor (_20509_, _20508_, _20473_);
  nor (_20510_, _20509_, _04778_);
  or (_20511_, _20510_, _20507_);
  and (_20512_, _20511_, _04790_);
  and (_20513_, _13402_, _05480_);
  nor (_20515_, _20513_, _20473_);
  nor (_20516_, _20515_, _04790_);
  or (_20517_, _20516_, _20512_);
  and (_20518_, _20517_, _04792_);
  and (_20519_, _08736_, _05480_);
  nor (_20520_, _20519_, _20473_);
  nor (_20521_, _20520_, _04792_);
  nor (_20522_, _20521_, _20518_);
  nor (_20523_, _20522_, _03908_);
  nor (_20524_, _20473_, _08322_);
  not (_20526_, _20524_);
  nor (_20527_, _20509_, _03909_);
  and (_20528_, _20527_, _20526_);
  nor (_20529_, _20528_, _20523_);
  nor (_20530_, _20529_, _04027_);
  nor (_20531_, _20475_, _04785_);
  and (_20532_, _20531_, _20526_);
  nor (_20533_, _20532_, _03914_);
  not (_20534_, _20533_);
  nor (_20535_, _20534_, _20530_);
  or (_20537_, _13401_, _09271_);
  nor (_20538_, _20473_, _06567_);
  and (_20539_, _20538_, _20537_);
  or (_20540_, _20539_, _04011_);
  nor (_20541_, _20540_, _20535_);
  nor (_20542_, _08735_, _09271_);
  nor (_20543_, _20542_, _20473_);
  nor (_20544_, _20543_, _06572_);
  or (_20545_, _20544_, _03773_);
  nor (_20546_, _20545_, _20541_);
  and (_20548_, _20482_, _03773_);
  or (_20549_, _20548_, _03772_);
  nor (_20550_, _20549_, _20546_);
  nor (_20551_, _13460_, _19990_);
  nor (_20552_, _20551_, _20473_);
  nor (_20553_, _20552_, _04060_);
  or (_20554_, _20553_, _20550_);
  or (_20555_, _20554_, _43156_);
  or (_20556_, _43152_, \oc8051_golden_model_1.TL0 [6]);
  and (_20557_, _20556_, _41894_);
  and (_43436_, _20557_, _20555_);
  not (_20559_, \oc8051_golden_model_1.TL1 [0]);
  nor (_20560_, _05587_, _20559_);
  and (_20561_, _05716_, _05587_);
  nor (_20562_, _20561_, _20560_);
  and (_20563_, _20562_, _17157_);
  and (_20564_, _05587_, _04700_);
  nor (_20565_, _20564_, _20560_);
  and (_20566_, _20565_, _08474_);
  nor (_20567_, _20562_, _04722_);
  nor (_20569_, _04707_, _20559_);
  and (_20570_, _05461_, \oc8051_golden_model_1.ACC [0]);
  nor (_20571_, _20570_, _20560_);
  nor (_20572_, _20571_, _04708_);
  nor (_20573_, _20572_, _20569_);
  nor (_20574_, _20573_, _03850_);
  or (_20575_, _20574_, _20567_);
  and (_20576_, _20575_, _04733_);
  nor (_20577_, _20565_, _04733_);
  or (_20578_, _20577_, _20576_);
  and (_20580_, _20578_, _03855_);
  nor (_20581_, _20571_, _03855_);
  or (_20582_, _20581_, _07927_);
  nor (_20583_, _20582_, _20580_);
  nor (_20584_, _20583_, _20566_);
  nor (_20585_, _20560_, _03738_);
  or (_20586_, _06733_, _09351_);
  nand (_20587_, _20586_, _20585_);
  and (_20588_, _20587_, _20584_);
  and (_20589_, _20588_, _03820_);
  not (_20591_, _05461_);
  nor (_20592_, _12164_, _20591_);
  nor (_20593_, _20592_, _20560_);
  nor (_20594_, _20593_, _03820_);
  or (_20595_, _20594_, _20589_);
  and (_20596_, _20595_, _04778_);
  and (_20597_, _05461_, _06479_);
  nor (_20598_, _20597_, _20560_);
  nor (_20599_, _20598_, _04778_);
  or (_20600_, _20599_, _20596_);
  and (_20602_, _20600_, _04790_);
  and (_20603_, _12178_, _05461_);
  nor (_20604_, _20603_, _20560_);
  nor (_20605_, _20604_, _04790_);
  or (_20606_, _20605_, _20602_);
  and (_20607_, _20606_, _04792_);
  nor (_20608_, _10488_, _09351_);
  nor (_20609_, _20608_, _20560_);
  and (_20610_, _20570_, _10262_);
  or (_20611_, _20610_, _04792_);
  nor (_20613_, _20611_, _20609_);
  nor (_20614_, _20613_, _20607_);
  nor (_20615_, _20614_, _03908_);
  and (_20616_, _12058_, _05461_);
  or (_20617_, _20616_, _20560_);
  and (_20618_, _20617_, _03908_);
  or (_20619_, _20618_, _20615_);
  and (_20620_, _20619_, _04785_);
  nor (_20621_, _20610_, _20560_);
  nor (_20622_, _20621_, _04785_);
  or (_20624_, _20622_, _20620_);
  and (_20625_, _20624_, _06567_);
  nor (_20626_, _12177_, _20591_);
  nor (_20627_, _20626_, _20560_);
  nor (_20628_, _20627_, _06567_);
  or (_20629_, _20628_, _20625_);
  and (_20630_, _20629_, _06572_);
  nor (_20631_, _20609_, _06572_);
  nor (_20632_, _20631_, _17157_);
  not (_20633_, _20632_);
  nor (_20635_, _20633_, _20630_);
  nor (_20636_, _20635_, _20563_);
  or (_20637_, _20636_, _43156_);
  or (_20638_, _43152_, \oc8051_golden_model_1.TL1 [0]);
  and (_20639_, _20638_, _41894_);
  and (_43437_, _20639_, _20637_);
  nor (_20640_, _05587_, \oc8051_golden_model_1.TL1 [1]);
  nor (_20641_, _20640_, _04778_);
  and (_20642_, _05587_, _04595_);
  not (_20643_, _20642_);
  and (_20645_, _20643_, _20641_);
  not (_20646_, \oc8051_golden_model_1.TL1 [1]);
  nor (_20647_, _05587_, _20646_);
  nor (_20648_, _20647_, _03738_);
  or (_20649_, _06688_, _09351_);
  and (_20650_, _20649_, _20648_);
  not (_20651_, _20650_);
  and (_20652_, _05461_, \oc8051_golden_model_1.ACC [1]);
  nor (_20653_, _20652_, _20647_);
  nor (_20654_, _20653_, _04708_);
  nor (_20656_, _04707_, _20646_);
  or (_20657_, _20656_, _20654_);
  and (_20658_, _20657_, _04722_);
  and (_20659_, _12262_, _05461_);
  nor (_20660_, _20659_, _20640_);
  and (_20661_, _20660_, _03850_);
  or (_20662_, _20661_, _20658_);
  and (_20663_, _20662_, _04733_);
  and (_20664_, _05587_, _04900_);
  nor (_20665_, _20664_, _20647_);
  nor (_20667_, _20665_, _04733_);
  nor (_20668_, _20667_, _20663_);
  nor (_20669_, _20668_, _03854_);
  nor (_20670_, _20653_, _03855_);
  or (_20671_, _20670_, _07927_);
  or (_20672_, _20671_, _20669_);
  and (_20673_, _20665_, _08474_);
  nor (_20674_, _20673_, _03455_);
  and (_20675_, _20674_, _20672_);
  and (_20676_, _20675_, _20651_);
  nor (_20678_, _12352_, _20591_);
  nor (_20679_, _20678_, _20647_);
  nor (_20680_, _20679_, _03820_);
  nor (_20681_, _20680_, _20676_);
  nor (_20682_, _20681_, _03903_);
  nor (_20683_, _20682_, _20645_);
  nor (_20684_, _20683_, _03897_);
  and (_20685_, _12366_, _05461_);
  or (_20686_, _20685_, _20647_);
  and (_20687_, _20686_, _03897_);
  nor (_20689_, _20687_, _20684_);
  nor (_20690_, _20689_, _04018_);
  nor (_20691_, _08751_, _09351_);
  nor (_20692_, _20691_, _20647_);
  and (_20693_, _20652_, _08366_);
  nor (_20694_, _20693_, _20692_);
  and (_20695_, _20694_, _04018_);
  or (_20696_, _20695_, _20690_);
  and (_20697_, _20696_, _03909_);
  and (_20698_, _12244_, _05461_);
  or (_20700_, _20698_, _20647_);
  and (_20701_, _20700_, _03908_);
  or (_20702_, _20701_, _20697_);
  and (_20703_, _20702_, _04785_);
  nor (_20704_, _20693_, _20647_);
  nor (_20705_, _20704_, _04785_);
  or (_20706_, _20705_, _20703_);
  and (_20707_, _20706_, _06567_);
  nor (_20708_, _12365_, _20591_);
  or (_20709_, _20708_, _20647_);
  and (_20711_, _20709_, _03914_);
  or (_20712_, _20711_, _20707_);
  and (_20713_, _20712_, _06572_);
  nor (_20714_, _20692_, _06572_);
  or (_20715_, _20714_, _20713_);
  nor (_20716_, _20715_, _03773_);
  nor (_20717_, _20660_, _03774_);
  or (_20718_, _20717_, _03772_);
  nor (_20719_, _20718_, _20716_);
  nor (_20720_, _20659_, _20647_);
  nor (_20722_, _20720_, _04060_);
  or (_20723_, _20722_, _20719_);
  or (_20724_, _20723_, _43156_);
  or (_20725_, _43152_, \oc8051_golden_model_1.TL1 [1]);
  and (_20726_, _20725_, _41894_);
  and (_43439_, _20726_, _20724_);
  not (_20727_, \oc8051_golden_model_1.TL1 [2]);
  nor (_20728_, _05587_, _20727_);
  nor (_20729_, _20728_, _03738_);
  or (_20730_, _06824_, _09351_);
  and (_20732_, _20730_, _20729_);
  and (_20733_, _05461_, \oc8051_golden_model_1.ACC [2]);
  nor (_20734_, _20733_, _20728_);
  nor (_20735_, _20734_, _04708_);
  nor (_20736_, _04707_, _20727_);
  or (_20737_, _20736_, _20735_);
  and (_20738_, _20737_, _04722_);
  nor (_20739_, _12471_, _09351_);
  nor (_20740_, _20739_, _20728_);
  nor (_20741_, _20740_, _04722_);
  or (_20743_, _20741_, _20738_);
  and (_20744_, _20743_, _04733_);
  and (_20745_, _05587_, _05307_);
  nor (_20746_, _20745_, _20728_);
  nor (_20747_, _20746_, _04733_);
  nor (_20748_, _20747_, _20744_);
  nor (_20749_, _20748_, _03854_);
  nor (_20750_, _20734_, _03855_);
  or (_20751_, _20750_, _07927_);
  nor (_20752_, _20751_, _20749_);
  and (_20754_, _20746_, _08474_);
  or (_20755_, _20754_, _03455_);
  or (_20756_, _20755_, _20752_);
  nor (_20757_, _20756_, _20732_);
  nor (_20758_, _12572_, _09351_);
  nor (_20759_, _20758_, _20728_);
  nor (_20760_, _20759_, _03820_);
  or (_20761_, _20760_, _20757_);
  and (_20762_, _20761_, _04778_);
  and (_20763_, _05461_, _06495_);
  nor (_20765_, _20763_, _20728_);
  nor (_20766_, _20765_, _04778_);
  or (_20767_, _20766_, _20762_);
  nor (_20768_, _20767_, _03897_);
  nand (_20769_, _12586_, _05587_);
  nor (_20770_, _20728_, _04790_);
  and (_20771_, _20770_, _20769_);
  or (_20772_, _20771_, _04018_);
  nor (_20773_, _20772_, _20768_);
  and (_20774_, _08748_, _05461_);
  nor (_20776_, _20774_, _20728_);
  nor (_20777_, _20776_, _04792_);
  nor (_20778_, _20777_, _20773_);
  nor (_20779_, _20778_, _03908_);
  nor (_20780_, _20728_, _05765_);
  not (_20781_, _20780_);
  nor (_20782_, _20765_, _03909_);
  and (_20783_, _20782_, _20781_);
  nor (_20784_, _20783_, _20779_);
  nor (_20785_, _20784_, _04027_);
  nor (_20787_, _20734_, _04785_);
  and (_20788_, _20787_, _20781_);
  or (_20789_, _20788_, _20785_);
  and (_20790_, _20789_, _06567_);
  nor (_20791_, _12585_, _20591_);
  nor (_20792_, _20791_, _20728_);
  nor (_20793_, _20792_, _06567_);
  or (_20794_, _20793_, _20790_);
  and (_20795_, _20794_, _06572_);
  nor (_20796_, _08747_, _09351_);
  nor (_20798_, _20796_, _20728_);
  nor (_20799_, _20798_, _06572_);
  or (_20800_, _20799_, _03773_);
  nor (_20801_, _20800_, _20795_);
  and (_20802_, _20740_, _03773_);
  or (_20803_, _20802_, _03772_);
  nor (_20804_, _20803_, _20801_);
  and (_20805_, _12642_, _05461_);
  nor (_20806_, _20805_, _20728_);
  nor (_20807_, _20806_, _04060_);
  or (_20809_, _20807_, _20804_);
  or (_20810_, _20809_, _43156_);
  or (_20811_, _43152_, \oc8051_golden_model_1.TL1 [2]);
  and (_20812_, _20811_, _41894_);
  and (_43440_, _20812_, _20810_);
  not (_20813_, \oc8051_golden_model_1.TL1 [3]);
  nor (_20814_, _05587_, _20813_);
  and (_20815_, _05461_, \oc8051_golden_model_1.ACC [3]);
  nor (_20816_, _20815_, _20814_);
  nor (_20817_, _20816_, _04708_);
  nor (_20819_, _04707_, _20813_);
  or (_20820_, _20819_, _20817_);
  and (_20821_, _20820_, _04722_);
  nor (_20822_, _12681_, _09351_);
  nor (_20823_, _20822_, _20814_);
  nor (_20824_, _20823_, _04722_);
  or (_20825_, _20824_, _20821_);
  and (_20826_, _20825_, _04733_);
  and (_20827_, _05587_, _05119_);
  nor (_20828_, _20827_, _20814_);
  nor (_20830_, _20828_, _04733_);
  nor (_20831_, _20830_, _20826_);
  nor (_20832_, _20831_, _03854_);
  nor (_20833_, _20816_, _03855_);
  or (_20834_, _20833_, _07927_);
  nor (_20835_, _20834_, _20832_);
  nor (_20836_, _20814_, _03738_);
  or (_20837_, _06779_, _09351_);
  and (_20838_, _20837_, _20836_);
  and (_20839_, _20828_, _08474_);
  or (_20841_, _20839_, _03455_);
  or (_20842_, _20841_, _20838_);
  nor (_20843_, _20842_, _20835_);
  nor (_20844_, _12775_, _09351_);
  nor (_20845_, _20844_, _20814_);
  nor (_20846_, _20845_, _03820_);
  or (_20847_, _20846_, _20843_);
  and (_20848_, _20847_, _04778_);
  and (_20849_, _05461_, _06345_);
  nor (_20850_, _20849_, _20814_);
  nor (_20852_, _20850_, _04778_);
  or (_20853_, _20852_, _20848_);
  nor (_20854_, _20853_, _03897_);
  nand (_20855_, _12789_, _05587_);
  nor (_20856_, _20814_, _04790_);
  and (_20857_, _20856_, _20855_);
  or (_20858_, _20857_, _04018_);
  nor (_20859_, _20858_, _20854_);
  and (_20860_, _10491_, _05461_);
  nor (_20861_, _20860_, _20814_);
  nor (_20863_, _20861_, _04792_);
  nor (_20864_, _20863_, _20859_);
  nor (_20865_, _20864_, _03908_);
  nor (_20866_, _20814_, _05622_);
  not (_20867_, _20866_);
  nor (_20868_, _20850_, _03909_);
  and (_20869_, _20868_, _20867_);
  nor (_20870_, _20869_, _20865_);
  nor (_20871_, _20870_, _04027_);
  nor (_20872_, _20816_, _04785_);
  and (_20874_, _20872_, _20867_);
  or (_20875_, _20874_, _20871_);
  and (_20876_, _20875_, _06567_);
  nor (_20877_, _12788_, _20591_);
  nor (_20878_, _20877_, _20814_);
  nor (_20879_, _20878_, _06567_);
  or (_20880_, _20879_, _20876_);
  and (_20881_, _20880_, _06572_);
  nor (_20882_, _08742_, _09351_);
  nor (_20883_, _20882_, _20814_);
  nor (_20885_, _20883_, _06572_);
  or (_20886_, _20885_, _03773_);
  nor (_20887_, _20886_, _20881_);
  and (_20888_, _20823_, _03773_);
  or (_20889_, _20888_, _03772_);
  nor (_20890_, _20889_, _20887_);
  and (_20891_, _12848_, _05461_);
  nor (_20892_, _20891_, _20814_);
  nor (_20893_, _20892_, _04060_);
  or (_20894_, _20893_, _20890_);
  or (_20896_, _20894_, _43156_);
  or (_20897_, _43152_, \oc8051_golden_model_1.TL1 [3]);
  and (_20898_, _20897_, _41894_);
  and (_43441_, _20898_, _20896_);
  not (_20899_, \oc8051_golden_model_1.TL1 [4]);
  nor (_20900_, _05587_, _20899_);
  and (_20901_, _05461_, \oc8051_golden_model_1.ACC [4]);
  nor (_20902_, _20901_, _20900_);
  nor (_20903_, _20902_, _04708_);
  nor (_20904_, _04707_, _20899_);
  or (_20906_, _20904_, _20903_);
  and (_20907_, _20906_, _04722_);
  nor (_20908_, _12891_, _09351_);
  nor (_20909_, _20908_, _20900_);
  nor (_20910_, _20909_, _04722_);
  or (_20911_, _20910_, _20907_);
  and (_20912_, _20911_, _04733_);
  and (_20913_, _05950_, _05587_);
  nor (_20914_, _20913_, _20900_);
  nor (_20915_, _20914_, _04733_);
  nor (_20916_, _20915_, _20912_);
  nor (_20917_, _20916_, _03854_);
  nor (_20918_, _20902_, _03855_);
  or (_20919_, _20918_, _07927_);
  or (_20920_, _20919_, _20917_);
  nor (_20921_, _20900_, _03738_);
  or (_20922_, _06918_, _09351_);
  and (_20923_, _20922_, _20921_);
  and (_20924_, _20914_, _08474_);
  or (_20925_, _20924_, _03455_);
  nor (_20927_, _20925_, _20923_);
  and (_20928_, _20927_, _20920_);
  nor (_20929_, _12982_, _09351_);
  nor (_20930_, _20929_, _20900_);
  nor (_20931_, _20930_, _03820_);
  or (_20932_, _20931_, _20928_);
  and (_20933_, _20932_, _04778_);
  and (_20934_, _06456_, _05461_);
  nor (_20935_, _20934_, _20900_);
  nor (_20936_, _20935_, _04778_);
  or (_20938_, _20936_, _20933_);
  nor (_20939_, _20938_, _03897_);
  nand (_20940_, _12997_, _05587_);
  nor (_20941_, _20900_, _04790_);
  and (_20942_, _20941_, _20940_);
  or (_20943_, _20942_, _04018_);
  nor (_20944_, _20943_, _20939_);
  and (_20945_, _08741_, _05461_);
  nor (_20946_, _20945_, _20900_);
  nor (_20947_, _20946_, _04792_);
  nor (_20949_, _20947_, _20944_);
  nor (_20950_, _20949_, _03908_);
  nor (_20951_, _20900_, _08336_);
  not (_20952_, _20951_);
  nor (_20953_, _20935_, _03909_);
  and (_20954_, _20953_, _20952_);
  nor (_20955_, _20954_, _20950_);
  nor (_20956_, _20955_, _04027_);
  nor (_20957_, _20902_, _04785_);
  and (_20958_, _20957_, _20952_);
  or (_20959_, _20958_, _20956_);
  and (_20960_, _20959_, _06567_);
  nor (_20961_, _12996_, _20591_);
  nor (_20962_, _20961_, _20900_);
  nor (_20963_, _20962_, _06567_);
  or (_20964_, _20963_, _20960_);
  and (_20965_, _20964_, _06572_);
  nor (_20966_, _08740_, _09351_);
  nor (_20967_, _20966_, _20900_);
  nor (_20968_, _20967_, _06572_);
  or (_20970_, _20968_, _03773_);
  nor (_20971_, _20970_, _20965_);
  and (_20972_, _20909_, _03773_);
  or (_20973_, _20972_, _03772_);
  nor (_20974_, _20973_, _20971_);
  and (_20975_, _13056_, _05461_);
  nor (_20976_, _20975_, _20900_);
  nor (_20977_, _20976_, _04060_);
  or (_20978_, _20977_, _20974_);
  or (_20979_, _20978_, _43156_);
  or (_20981_, _43152_, \oc8051_golden_model_1.TL1 [4]);
  and (_20982_, _20981_, _41894_);
  and (_43442_, _20982_, _20979_);
  not (_20983_, \oc8051_golden_model_1.TL1 [5]);
  nor (_20984_, _05587_, _20983_);
  nor (_20985_, _13090_, _09351_);
  nor (_20986_, _20985_, _20984_);
  nor (_20987_, _20986_, _04722_);
  nor (_20988_, _04707_, _20983_);
  and (_20989_, _05461_, \oc8051_golden_model_1.ACC [5]);
  nor (_20990_, _20989_, _20984_);
  nor (_20991_, _20990_, _04708_);
  nor (_20992_, _20991_, _20988_);
  nor (_20993_, _20992_, _03850_);
  or (_20994_, _20993_, _20987_);
  and (_20995_, _20994_, _04733_);
  and (_20996_, _05857_, _05587_);
  nor (_20997_, _20996_, _20984_);
  nor (_20998_, _20997_, _04733_);
  or (_20999_, _20998_, _20995_);
  and (_21001_, _20999_, _03855_);
  nor (_21002_, _20990_, _03855_);
  or (_21003_, _21002_, _07927_);
  or (_21004_, _21003_, _21001_);
  nor (_21005_, _20984_, _03738_);
  or (_21006_, _06873_, _09351_);
  and (_21007_, _21006_, _21005_);
  and (_21008_, _20997_, _08474_);
  or (_21009_, _21008_, _03455_);
  nor (_21010_, _21009_, _21007_);
  and (_21012_, _21010_, _21004_);
  nor (_21013_, _13182_, _09351_);
  nor (_21014_, _21013_, _20984_);
  nor (_21015_, _21014_, _03820_);
  or (_21016_, _21015_, _21012_);
  and (_21017_, _21016_, _04778_);
  and (_21018_, _06447_, _05461_);
  nor (_21019_, _21018_, _20984_);
  nor (_21020_, _21019_, _04778_);
  or (_21021_, _21020_, _21017_);
  nor (_21022_, _21021_, _03897_);
  nand (_21023_, _13196_, _05587_);
  nor (_21024_, _20984_, _04790_);
  and (_21025_, _21024_, _21023_);
  or (_21026_, _21025_, _04018_);
  nor (_21027_, _21026_, _21022_);
  and (_21028_, _10493_, _05461_);
  nor (_21029_, _21028_, _20984_);
  nor (_21030_, _21029_, _04792_);
  nor (_21031_, _21030_, _21027_);
  nor (_21033_, _21031_, _03908_);
  nor (_21034_, _20984_, _08335_);
  not (_21035_, _21034_);
  nor (_21036_, _21019_, _03909_);
  and (_21037_, _21036_, _21035_);
  nor (_21038_, _21037_, _21033_);
  nor (_21039_, _21038_, _04027_);
  nor (_21040_, _20990_, _04785_);
  and (_21041_, _21040_, _21035_);
  or (_21042_, _21041_, _21039_);
  and (_21044_, _21042_, _06567_);
  nor (_21045_, _13195_, _20591_);
  nor (_21046_, _21045_, _20984_);
  nor (_21047_, _21046_, _06567_);
  or (_21048_, _21047_, _21044_);
  and (_21049_, _21048_, _06572_);
  nor (_21050_, _08738_, _09351_);
  nor (_21051_, _21050_, _20984_);
  nor (_21052_, _21051_, _06572_);
  nor (_21053_, _21052_, _21049_);
  nor (_21054_, _21053_, _03773_);
  nor (_21055_, _20986_, _03774_);
  or (_21056_, _21055_, _03772_);
  nor (_21057_, _21056_, _21054_);
  and (_21058_, _13255_, _05461_);
  nor (_21059_, _21058_, _20984_);
  and (_21060_, _21059_, _03772_);
  nor (_21061_, _21060_, _21057_);
  or (_21062_, _21061_, _43156_);
  or (_21063_, _43152_, \oc8051_golden_model_1.TL1 [5]);
  and (_21065_, _21063_, _41894_);
  and (_43443_, _21065_, _21062_);
  not (_21066_, \oc8051_golden_model_1.TL1 [6]);
  nor (_21067_, _05587_, _21066_);
  and (_21068_, _05461_, \oc8051_golden_model_1.ACC [6]);
  nor (_21069_, _21068_, _21067_);
  nor (_21070_, _21069_, _04708_);
  nor (_21071_, _04707_, _21066_);
  or (_21072_, _21071_, _21070_);
  and (_21073_, _21072_, _04722_);
  nor (_21075_, _13293_, _09351_);
  nor (_21076_, _21075_, _21067_);
  nor (_21077_, _21076_, _04722_);
  or (_21078_, _21077_, _21073_);
  and (_21079_, _21078_, _04733_);
  and (_21080_, _06065_, _05587_);
  nor (_21081_, _21080_, _21067_);
  nor (_21082_, _21081_, _04733_);
  nor (_21083_, _21082_, _21079_);
  nor (_21084_, _21083_, _03854_);
  nor (_21085_, _21069_, _03855_);
  or (_21086_, _21085_, _07927_);
  or (_21087_, _21086_, _21084_);
  nor (_21088_, _21067_, _03738_);
  nand (_21089_, _06641_, _05587_);
  and (_21090_, _21089_, _21088_);
  and (_21091_, _21081_, _08474_);
  or (_21092_, _21091_, _03455_);
  nor (_21093_, _21092_, _21090_);
  and (_21094_, _21093_, _21087_);
  nor (_21096_, _13387_, _09351_);
  nor (_21097_, _21096_, _21067_);
  nor (_21098_, _21097_, _03820_);
  or (_21099_, _21098_, _21094_);
  and (_21100_, _21099_, _04778_);
  and (_21101_, _13394_, _05461_);
  nor (_21102_, _21101_, _21067_);
  nor (_21103_, _21102_, _04778_);
  or (_21104_, _21103_, _21100_);
  nor (_21105_, _21104_, _03897_);
  nand (_21107_, _13402_, _05587_);
  nor (_21108_, _21067_, _04790_);
  and (_21109_, _21108_, _21107_);
  or (_21110_, _21109_, _04018_);
  nor (_21111_, _21110_, _21105_);
  and (_21112_, _08736_, _05461_);
  nor (_21113_, _21112_, _21067_);
  nor (_21114_, _21113_, _04792_);
  nor (_21115_, _21114_, _21111_);
  nor (_21116_, _21115_, _03908_);
  nor (_21117_, _21067_, _08322_);
  not (_21118_, _21117_);
  nor (_21119_, _21102_, _03909_);
  and (_21120_, _21119_, _21118_);
  nor (_21121_, _21120_, _21116_);
  nor (_21122_, _21121_, _04027_);
  nor (_21123_, _21069_, _04785_);
  and (_21124_, _21123_, _21118_);
  nor (_21125_, _21124_, _03914_);
  not (_21126_, _21125_);
  nor (_21128_, _21126_, _21122_);
  or (_21129_, _13401_, _09351_);
  nor (_21130_, _21067_, _06567_);
  and (_21131_, _21130_, _21129_);
  or (_21132_, _21131_, _04011_);
  nor (_21133_, _21132_, _21128_);
  nor (_21134_, _08735_, _09351_);
  nor (_21135_, _21134_, _21067_);
  nor (_21136_, _21135_, _06572_);
  or (_21137_, _21136_, _03773_);
  nor (_21139_, _21137_, _21133_);
  and (_21140_, _21076_, _03773_);
  or (_21141_, _21140_, _03772_);
  nor (_21142_, _21141_, _21139_);
  nor (_21143_, _13460_, _20591_);
  nor (_21144_, _21143_, _21067_);
  nor (_21145_, _21144_, _04060_);
  or (_21146_, _21145_, _21142_);
  or (_21147_, _21146_, _43156_);
  or (_21148_, _43152_, \oc8051_golden_model_1.TL1 [6]);
  and (_21149_, _21148_, _41894_);
  and (_43444_, _21149_, _21147_);
  not (_21150_, \oc8051_golden_model_1.TH0 [0]);
  nor (_21151_, _05451_, _21150_);
  and (_21152_, _05716_, _05451_);
  nor (_21153_, _21152_, _21151_);
  and (_21154_, _21153_, _17157_);
  and (_21155_, _06962_, _05451_);
  nor (_21156_, _21151_, _03738_);
  not (_21157_, _21156_);
  nor (_21159_, _21157_, _21155_);
  and (_21160_, _05451_, _04700_);
  nor (_21161_, _21160_, _21151_);
  and (_21162_, _21161_, _08474_);
  nor (_21163_, _21153_, _04722_);
  nor (_21164_, _04707_, _21150_);
  and (_21165_, _05451_, \oc8051_golden_model_1.ACC [0]);
  nor (_21166_, _21165_, _21151_);
  nor (_21167_, _21166_, _04708_);
  nor (_21168_, _21167_, _21164_);
  nor (_21170_, _21168_, _03850_);
  or (_21171_, _21170_, _21163_);
  and (_21172_, _21171_, _04733_);
  nor (_21173_, _21161_, _04733_);
  or (_21174_, _21173_, _21172_);
  and (_21175_, _21174_, _03855_);
  nor (_21176_, _21166_, _03855_);
  or (_21177_, _21176_, _07927_);
  nor (_21178_, _21177_, _21175_);
  nor (_21179_, _21178_, _21162_);
  not (_21180_, _21179_);
  nor (_21181_, _21180_, _21159_);
  and (_21182_, _21181_, _03820_);
  nor (_21183_, _12164_, _09432_);
  nor (_21184_, _21183_, _21151_);
  nor (_21185_, _21184_, _03820_);
  or (_21186_, _21185_, _21182_);
  and (_21187_, _21186_, _04778_);
  and (_21188_, _05451_, _06479_);
  nor (_21189_, _21188_, _21151_);
  nor (_21191_, _21189_, _04778_);
  or (_21192_, _21191_, _21187_);
  and (_21193_, _21192_, _04790_);
  and (_21194_, _12178_, _05451_);
  nor (_21195_, _21194_, _21151_);
  nor (_21196_, _21195_, _04790_);
  or (_21197_, _21196_, _21193_);
  and (_21198_, _21197_, _04792_);
  nor (_21199_, _10488_, _09432_);
  nor (_21200_, _21199_, _21151_);
  not (_21202_, _21200_);
  and (_21203_, _08753_, _05451_);
  nor (_21204_, _21203_, _04792_);
  and (_21205_, _21204_, _21202_);
  nor (_21206_, _21205_, _21198_);
  nor (_21207_, _21206_, _03908_);
  and (_21208_, _12058_, _05451_);
  or (_21209_, _21208_, _21151_);
  and (_21210_, _21209_, _03908_);
  or (_21211_, _21210_, _21207_);
  and (_21212_, _21211_, _04785_);
  nor (_21213_, _21203_, _21151_);
  nor (_21214_, _21213_, _04785_);
  or (_21215_, _21214_, _21212_);
  and (_21216_, _21215_, _06567_);
  nor (_21217_, _12177_, _09432_);
  nor (_21218_, _21217_, _21151_);
  nor (_21219_, _21218_, _06567_);
  or (_21220_, _21219_, _21216_);
  and (_21221_, _21220_, _06572_);
  nor (_21223_, _21200_, _06572_);
  nor (_21224_, _21223_, _17157_);
  not (_21225_, _21224_);
  nor (_21226_, _21225_, _21221_);
  nor (_21227_, _21226_, _21154_);
  or (_21228_, _21227_, _43156_);
  or (_21229_, _43152_, \oc8051_golden_model_1.TH0 [0]);
  and (_21230_, _21229_, _41894_);
  and (_43447_, _21230_, _21228_);
  and (_21231_, _06961_, _05451_);
  not (_21233_, \oc8051_golden_model_1.TH0 [1]);
  nor (_21234_, _05451_, _21233_);
  nor (_21235_, _21234_, _03738_);
  not (_21236_, _21235_);
  nor (_21237_, _21236_, _21231_);
  not (_21238_, _21237_);
  and (_21239_, _05451_, \oc8051_golden_model_1.ACC [1]);
  nor (_21240_, _21239_, _21234_);
  nor (_21241_, _21240_, _04708_);
  nor (_21242_, _04707_, _21233_);
  or (_21243_, _21242_, _21241_);
  and (_21244_, _21243_, _04722_);
  nor (_21245_, _05451_, \oc8051_golden_model_1.TH0 [1]);
  and (_21246_, _12262_, _05451_);
  nor (_21247_, _21246_, _21245_);
  and (_21248_, _21247_, _03850_);
  or (_21249_, _21248_, _21244_);
  and (_21250_, _21249_, _04733_);
  and (_21251_, _05451_, _04900_);
  nor (_21252_, _21251_, _21234_);
  nor (_21254_, _21252_, _04733_);
  nor (_21255_, _21254_, _21250_);
  nor (_21256_, _21255_, _03854_);
  nor (_21257_, _21240_, _03855_);
  or (_21258_, _21257_, _07927_);
  or (_21259_, _21258_, _21256_);
  and (_21260_, _21252_, _08474_);
  nor (_21261_, _21260_, _03455_);
  and (_21262_, _21261_, _21259_);
  and (_21263_, _21262_, _21238_);
  and (_21265_, _12352_, _05451_);
  or (_21266_, _21265_, _03820_);
  nor (_21267_, _21266_, _21245_);
  nor (_21268_, _21267_, _21263_);
  nor (_21269_, _21268_, _03903_);
  and (_21270_, _05451_, _04595_);
  not (_21271_, _21270_);
  nor (_21272_, _21245_, _04778_);
  and (_21273_, _21272_, _21271_);
  nor (_21274_, _21273_, _21269_);
  nor (_21275_, _21274_, _03897_);
  and (_21276_, _12366_, _05451_);
  or (_21277_, _21276_, _21234_);
  and (_21278_, _21277_, _03897_);
  nor (_21279_, _21278_, _21275_);
  nor (_21280_, _21279_, _04018_);
  nor (_21281_, _08751_, _09432_);
  nor (_21282_, _21281_, _21234_);
  and (_21283_, _08750_, _05451_);
  nor (_21284_, _21283_, _21282_);
  and (_21286_, _21284_, _04018_);
  or (_21287_, _21286_, _21280_);
  and (_21288_, _21287_, _03909_);
  and (_21289_, _12244_, _05451_);
  or (_21290_, _21289_, _21234_);
  and (_21291_, _21290_, _03908_);
  or (_21292_, _21291_, _21288_);
  and (_21293_, _21292_, _04785_);
  nor (_21294_, _21283_, _21234_);
  nor (_21295_, _21294_, _04785_);
  or (_21297_, _21295_, _21293_);
  and (_21298_, _21297_, _06567_);
  nor (_21299_, _12365_, _09432_);
  or (_21300_, _21299_, _21234_);
  and (_21301_, _21300_, _03914_);
  or (_21302_, _21301_, _21298_);
  and (_21303_, _21302_, _06572_);
  nor (_21304_, _21282_, _06572_);
  or (_21305_, _21304_, _21303_);
  nor (_21306_, _21305_, _03773_);
  nor (_21307_, _21247_, _03774_);
  or (_21308_, _21307_, _03772_);
  nor (_21309_, _21308_, _21306_);
  nor (_21310_, _21246_, _21234_);
  nor (_21311_, _21310_, _04060_);
  or (_21312_, _21311_, _21309_);
  or (_21313_, _21312_, _43156_);
  or (_21314_, _43152_, \oc8051_golden_model_1.TH0 [1]);
  and (_21315_, _21314_, _41894_);
  and (_43448_, _21315_, _21313_);
  and (_21317_, _06965_, _05451_);
  not (_21318_, \oc8051_golden_model_1.TH0 [2]);
  nor (_21319_, _05451_, _21318_);
  nor (_21320_, _21319_, _03738_);
  not (_21321_, _21320_);
  nor (_21322_, _21321_, _21317_);
  not (_21323_, _21322_);
  and (_21324_, _05451_, _05307_);
  nor (_21325_, _21324_, _21319_);
  and (_21326_, _21325_, _08474_);
  and (_21328_, _05451_, \oc8051_golden_model_1.ACC [2]);
  nor (_21329_, _21328_, _21319_);
  nor (_21330_, _21329_, _04708_);
  nor (_21331_, _04707_, _21318_);
  or (_21332_, _21331_, _21330_);
  and (_21333_, _21332_, _04722_);
  nor (_21334_, _12471_, _09432_);
  nor (_21335_, _21334_, _21319_);
  nor (_21336_, _21335_, _04722_);
  or (_21337_, _21336_, _21333_);
  and (_21339_, _21337_, _04733_);
  nor (_21340_, _21325_, _04733_);
  nor (_21341_, _21340_, _21339_);
  nor (_21342_, _21341_, _03854_);
  nor (_21343_, _21329_, _03855_);
  or (_21344_, _21343_, _07927_);
  nor (_21345_, _21344_, _21342_);
  nor (_21346_, _21345_, _21326_);
  and (_21347_, _21346_, _21323_);
  and (_21348_, _21347_, _03820_);
  nor (_21349_, _12572_, _09432_);
  nor (_21350_, _21349_, _21319_);
  nor (_21351_, _21350_, _03820_);
  or (_21352_, _21351_, _21348_);
  and (_21353_, _21352_, _04778_);
  and (_21354_, _05451_, _06495_);
  nor (_21355_, _21354_, _21319_);
  nor (_21356_, _21355_, _04778_);
  or (_21357_, _21356_, _21353_);
  and (_21358_, _21357_, _04790_);
  and (_21360_, _12586_, _05451_);
  nor (_21361_, _21360_, _21319_);
  nor (_21362_, _21361_, _04790_);
  or (_21363_, _21362_, _21358_);
  and (_21364_, _21363_, _04792_);
  and (_21365_, _08748_, _05451_);
  nor (_21366_, _21365_, _21319_);
  nor (_21367_, _21366_, _04792_);
  nor (_21368_, _21367_, _21364_);
  nor (_21369_, _21368_, _03908_);
  nor (_21371_, _21319_, _05765_);
  not (_21372_, _21371_);
  nor (_21373_, _21355_, _03909_);
  and (_21374_, _21373_, _21372_);
  nor (_21375_, _21374_, _21369_);
  nor (_21376_, _21375_, _04027_);
  nor (_21377_, _21329_, _04785_);
  and (_21378_, _21377_, _21372_);
  or (_21379_, _21378_, _21376_);
  and (_21380_, _21379_, _06567_);
  nor (_21382_, _12585_, _09432_);
  nor (_21383_, _21382_, _21319_);
  nor (_21384_, _21383_, _06567_);
  or (_21385_, _21384_, _21380_);
  and (_21386_, _21385_, _06572_);
  nor (_21387_, _08747_, _09432_);
  nor (_21388_, _21387_, _21319_);
  nor (_21389_, _21388_, _06572_);
  or (_21390_, _21389_, _03773_);
  nor (_21391_, _21390_, _21386_);
  and (_21393_, _21335_, _03773_);
  or (_21394_, _21393_, _03772_);
  nor (_21395_, _21394_, _21391_);
  and (_21396_, _12642_, _05451_);
  nor (_21397_, _21396_, _21319_);
  nor (_21398_, _21397_, _04060_);
  or (_21399_, _21398_, _21395_);
  or (_21400_, _21399_, _43156_);
  or (_21401_, _43152_, \oc8051_golden_model_1.TH0 [2]);
  and (_21402_, _21401_, _41894_);
  and (_43449_, _21402_, _21400_);
  not (_21405_, \oc8051_golden_model_1.TH0 [3]);
  nor (_21406_, _05451_, _21405_);
  and (_21407_, _05451_, \oc8051_golden_model_1.ACC [3]);
  nor (_21408_, _21407_, _21406_);
  nor (_21409_, _21408_, _04708_);
  nor (_21410_, _04707_, _21405_);
  or (_21411_, _21410_, _21409_);
  and (_21412_, _21411_, _04722_);
  nor (_21413_, _12681_, _09432_);
  nor (_21416_, _21413_, _21406_);
  nor (_21417_, _21416_, _04722_);
  or (_21418_, _21417_, _21412_);
  and (_21419_, _21418_, _04733_);
  and (_21420_, _05451_, _05119_);
  nor (_21421_, _21420_, _21406_);
  nor (_21422_, _21421_, _04733_);
  nor (_21423_, _21422_, _21419_);
  nor (_21424_, _21423_, _03854_);
  nor (_21425_, _21408_, _03855_);
  or (_21428_, _21425_, _07927_);
  or (_21429_, _21428_, _21424_);
  and (_21430_, _06964_, _05451_);
  nor (_21431_, _21406_, _03738_);
  not (_21432_, _21431_);
  nor (_21433_, _21432_, _21430_);
  and (_21434_, _21421_, _08474_);
  or (_21435_, _21434_, _03455_);
  nor (_21436_, _21435_, _21433_);
  and (_21437_, _21436_, _21429_);
  nor (_21439_, _12775_, _09432_);
  nor (_21440_, _21439_, _21406_);
  nor (_21441_, _21440_, _03820_);
  or (_21442_, _21441_, _21437_);
  and (_21443_, _21442_, _04778_);
  and (_21444_, _05451_, _06345_);
  nor (_21445_, _21444_, _21406_);
  nor (_21446_, _21445_, _04778_);
  or (_21447_, _21446_, _21443_);
  nor (_21448_, _21447_, _03897_);
  and (_21451_, _12789_, _05451_);
  or (_21452_, _21406_, _04790_);
  nor (_21453_, _21452_, _21451_);
  or (_21454_, _21453_, _04018_);
  nor (_21455_, _21454_, _21448_);
  and (_21456_, _10491_, _05451_);
  nor (_21457_, _21456_, _21406_);
  nor (_21458_, _21457_, _04792_);
  nor (_21459_, _21458_, _21455_);
  nor (_21460_, _21459_, _03908_);
  nor (_21461_, _21406_, _05622_);
  not (_21462_, _21461_);
  nor (_21463_, _21445_, _03909_);
  and (_21464_, _21463_, _21462_);
  nor (_21465_, _21464_, _21460_);
  nor (_21466_, _21465_, _04027_);
  nor (_21467_, _21408_, _04785_);
  and (_21468_, _21467_, _21462_);
  nor (_21469_, _21468_, _03914_);
  not (_21470_, _21469_);
  nor (_21472_, _21470_, _21466_);
  nor (_21473_, _12788_, _09432_);
  or (_21474_, _21406_, _06567_);
  nor (_21475_, _21474_, _21473_);
  or (_21476_, _21475_, _04011_);
  nor (_21477_, _21476_, _21472_);
  nor (_21478_, _08742_, _09432_);
  nor (_21479_, _21478_, _21406_);
  nor (_21480_, _21479_, _06572_);
  or (_21481_, _21480_, _03773_);
  nor (_21483_, _21481_, _21477_);
  and (_21484_, _21416_, _03773_);
  or (_21485_, _21484_, _03772_);
  nor (_21486_, _21485_, _21483_);
  and (_21487_, _12848_, _05451_);
  nor (_21488_, _21487_, _21406_);
  nor (_21489_, _21488_, _04060_);
  or (_21490_, _21489_, _21486_);
  or (_21491_, _21490_, _43156_);
  or (_21492_, _43152_, \oc8051_golden_model_1.TH0 [3]);
  and (_21494_, _21492_, _41894_);
  and (_43450_, _21494_, _21491_);
  not (_21495_, \oc8051_golden_model_1.TH0 [4]);
  nor (_21496_, _05451_, _21495_);
  and (_21497_, _05451_, \oc8051_golden_model_1.ACC [4]);
  nor (_21498_, _21497_, _21496_);
  nor (_21499_, _21498_, _04708_);
  nor (_21500_, _04707_, _21495_);
  or (_21501_, _21500_, _21499_);
  and (_21502_, _21501_, _04722_);
  nor (_21504_, _12891_, _09432_);
  nor (_21505_, _21504_, _21496_);
  nor (_21506_, _21505_, _04722_);
  or (_21507_, _21506_, _21502_);
  and (_21508_, _21507_, _04733_);
  and (_21509_, _05950_, _05451_);
  nor (_21510_, _21509_, _21496_);
  nor (_21511_, _21510_, _04733_);
  nor (_21512_, _21511_, _21508_);
  nor (_21513_, _21512_, _03854_);
  nor (_21515_, _21498_, _03855_);
  or (_21516_, _21515_, _07927_);
  or (_21517_, _21516_, _21513_);
  and (_21518_, _06969_, _05451_);
  nor (_21519_, _21496_, _03738_);
  not (_21520_, _21519_);
  nor (_21521_, _21520_, _21518_);
  and (_21522_, _21510_, _08474_);
  or (_21523_, _21522_, _03455_);
  nor (_21524_, _21523_, _21521_);
  and (_21526_, _21524_, _21517_);
  nor (_21527_, _12982_, _09432_);
  nor (_21528_, _21527_, _21496_);
  nor (_21529_, _21528_, _03820_);
  or (_21530_, _21529_, _21526_);
  and (_21531_, _21530_, _04778_);
  and (_21532_, _06456_, _05451_);
  nor (_21533_, _21532_, _21496_);
  nor (_21534_, _21533_, _04778_);
  or (_21535_, _21534_, _21531_);
  nor (_21537_, _21535_, _03897_);
  and (_21538_, _12997_, _05451_);
  or (_21539_, _21496_, _04790_);
  nor (_21540_, _21539_, _21538_);
  or (_21541_, _21540_, _04018_);
  nor (_21542_, _21541_, _21537_);
  and (_21543_, _08741_, _05451_);
  nor (_21544_, _21543_, _21496_);
  nor (_21545_, _21544_, _04792_);
  nor (_21546_, _21545_, _21542_);
  nor (_21548_, _21546_, _03908_);
  nor (_21549_, _21496_, _08336_);
  not (_21550_, _21549_);
  nor (_21551_, _21533_, _03909_);
  and (_21552_, _21551_, _21550_);
  nor (_21553_, _21552_, _21548_);
  nor (_21554_, _21553_, _04027_);
  nor (_21555_, _21498_, _04785_);
  and (_21556_, _21555_, _21550_);
  or (_21557_, _21556_, _21554_);
  and (_21559_, _21557_, _06567_);
  nor (_21560_, _12996_, _09432_);
  nor (_21561_, _21560_, _21496_);
  nor (_21562_, _21561_, _06567_);
  or (_21563_, _21562_, _21559_);
  and (_21564_, _21563_, _06572_);
  nor (_21565_, _08740_, _09432_);
  nor (_21566_, _21565_, _21496_);
  nor (_21567_, _21566_, _06572_);
  or (_21568_, _21567_, _03773_);
  nor (_21569_, _21568_, _21564_);
  and (_21570_, _21505_, _03773_);
  or (_21571_, _21570_, _03772_);
  nor (_21572_, _21571_, _21569_);
  and (_21573_, _13056_, _05451_);
  nor (_21574_, _21573_, _21496_);
  nor (_21575_, _21574_, _04060_);
  or (_21576_, _21575_, _21572_);
  or (_21577_, _21576_, _43156_);
  or (_21578_, _43152_, \oc8051_golden_model_1.TH0 [4]);
  and (_21579_, _21578_, _41894_);
  and (_43451_, _21579_, _21577_);
  not (_21580_, \oc8051_golden_model_1.TH0 [5]);
  nor (_21581_, _05451_, _21580_);
  and (_21582_, _05451_, \oc8051_golden_model_1.ACC [5]);
  nor (_21583_, _21582_, _21581_);
  nor (_21584_, _21583_, _04708_);
  nor (_21585_, _04707_, _21580_);
  or (_21586_, _21585_, _21584_);
  and (_21587_, _21586_, _04722_);
  nor (_21589_, _13090_, _09432_);
  nor (_21590_, _21589_, _21581_);
  nor (_21591_, _21590_, _04722_);
  or (_21592_, _21591_, _21587_);
  and (_21593_, _21592_, _04733_);
  and (_21594_, _05857_, _05451_);
  nor (_21595_, _21594_, _21581_);
  nor (_21596_, _21595_, _04733_);
  nor (_21597_, _21596_, _21593_);
  nor (_21598_, _21597_, _03854_);
  nor (_21600_, _21583_, _03855_);
  or (_21601_, _21600_, _07927_);
  or (_21602_, _21601_, _21598_);
  and (_21603_, _06968_, _05451_);
  nor (_21604_, _21581_, _03738_);
  not (_21605_, _21604_);
  nor (_21606_, _21605_, _21603_);
  and (_21607_, _21595_, _08474_);
  or (_21608_, _21607_, _03455_);
  nor (_21609_, _21608_, _21606_);
  and (_21611_, _21609_, _21602_);
  nor (_21612_, _13182_, _09432_);
  nor (_21613_, _21612_, _21581_);
  nor (_21614_, _21613_, _03820_);
  or (_21615_, _21614_, _21611_);
  and (_21616_, _21615_, _04778_);
  and (_21617_, _06447_, _05451_);
  nor (_21618_, _21617_, _21581_);
  nor (_21619_, _21618_, _04778_);
  or (_21620_, _21619_, _21616_);
  and (_21622_, _21620_, _04790_);
  and (_21623_, _13196_, _05451_);
  nor (_21624_, _21623_, _21581_);
  nor (_21625_, _21624_, _04790_);
  or (_21626_, _21625_, _21622_);
  and (_21627_, _21626_, _04792_);
  and (_21628_, _10493_, _05451_);
  nor (_21629_, _21628_, _21581_);
  nor (_21630_, _21629_, _04792_);
  nor (_21631_, _21630_, _21627_);
  nor (_21633_, _21631_, _03908_);
  nor (_21634_, _21581_, _08335_);
  not (_21635_, _21634_);
  nor (_21636_, _21618_, _03909_);
  and (_21637_, _21636_, _21635_);
  nor (_21638_, _21637_, _21633_);
  nor (_21639_, _21638_, _04027_);
  nor (_21640_, _21583_, _04785_);
  and (_21641_, _21640_, _21635_);
  or (_21642_, _21641_, _21639_);
  and (_21644_, _21642_, _06567_);
  nor (_21645_, _13195_, _09432_);
  nor (_21646_, _21645_, _21581_);
  nor (_21647_, _21646_, _06567_);
  or (_21648_, _21647_, _21644_);
  and (_21649_, _21648_, _06572_);
  nor (_21650_, _08738_, _09432_);
  nor (_21651_, _21650_, _21581_);
  nor (_21652_, _21651_, _06572_);
  nor (_21653_, _21652_, _21649_);
  nor (_21655_, _21653_, _03773_);
  nor (_21656_, _21590_, _03774_);
  or (_21657_, _21656_, _03772_);
  nor (_21658_, _21657_, _21655_);
  and (_21659_, _13255_, _05451_);
  nor (_21660_, _21659_, _21581_);
  and (_21661_, _21660_, _03772_);
  nor (_21662_, _21661_, _21658_);
  or (_21663_, _21662_, _43156_);
  or (_21664_, _43152_, \oc8051_golden_model_1.TH0 [5]);
  and (_21666_, _21664_, _41894_);
  and (_43452_, _21666_, _21663_);
  not (_21667_, \oc8051_golden_model_1.TH0 [6]);
  nor (_21668_, _05451_, _21667_);
  and (_21669_, _05451_, \oc8051_golden_model_1.ACC [6]);
  nor (_21670_, _21669_, _21668_);
  nor (_21671_, _21670_, _04708_);
  nor (_21672_, _04707_, _21667_);
  or (_21673_, _21672_, _21671_);
  and (_21674_, _21673_, _04722_);
  nor (_21676_, _13293_, _09432_);
  nor (_21677_, _21676_, _21668_);
  nor (_21678_, _21677_, _04722_);
  or (_21679_, _21678_, _21674_);
  and (_21680_, _21679_, _04733_);
  and (_21681_, _06065_, _05451_);
  nor (_21682_, _21681_, _21668_);
  nor (_21683_, _21682_, _04733_);
  nor (_21684_, _21683_, _21680_);
  nor (_21685_, _21684_, _03854_);
  nor (_21687_, _21670_, _03855_);
  or (_21688_, _21687_, _07927_);
  or (_21689_, _21688_, _21685_);
  and (_21690_, _06641_, _05451_);
  nor (_21691_, _21668_, _03738_);
  not (_21692_, _21691_);
  nor (_21693_, _21692_, _21690_);
  and (_21694_, _21682_, _08474_);
  or (_21695_, _21694_, _03455_);
  nor (_21696_, _21695_, _21693_);
  and (_21698_, _21696_, _21689_);
  nor (_21699_, _13387_, _09432_);
  nor (_21700_, _21699_, _21668_);
  nor (_21701_, _21700_, _03820_);
  or (_21702_, _21701_, _21698_);
  and (_21703_, _21702_, _04778_);
  and (_21704_, _13394_, _05451_);
  nor (_21705_, _21704_, _21668_);
  nor (_21706_, _21705_, _04778_);
  or (_21707_, _21706_, _21703_);
  and (_21709_, _21707_, _04790_);
  and (_21710_, _13402_, _05451_);
  nor (_21711_, _21710_, _21668_);
  nor (_21712_, _21711_, _04790_);
  or (_21713_, _21712_, _21709_);
  and (_21714_, _21713_, _04792_);
  and (_21715_, _08736_, _05451_);
  nor (_21716_, _21715_, _21668_);
  nor (_21717_, _21716_, _04792_);
  nor (_21718_, _21717_, _21714_);
  nor (_21720_, _21718_, _03908_);
  nor (_21721_, _21668_, _08322_);
  not (_21722_, _21721_);
  nor (_21723_, _21705_, _03909_);
  and (_21724_, _21723_, _21722_);
  nor (_21725_, _21724_, _21720_);
  nor (_21726_, _21725_, _04027_);
  nor (_21727_, _21670_, _04785_);
  and (_21728_, _21727_, _21722_);
  or (_21729_, _21728_, _21726_);
  and (_21731_, _21729_, _06567_);
  nor (_21732_, _13401_, _09432_);
  nor (_21733_, _21732_, _21668_);
  nor (_21734_, _21733_, _06567_);
  or (_21735_, _21734_, _21731_);
  and (_21736_, _21735_, _06572_);
  nor (_21737_, _08735_, _09432_);
  nor (_21738_, _21737_, _21668_);
  nor (_21739_, _21738_, _06572_);
  or (_21740_, _21739_, _03773_);
  nor (_21742_, _21740_, _21736_);
  and (_21743_, _21677_, _03773_);
  or (_21744_, _21743_, _03772_);
  nor (_21745_, _21744_, _21742_);
  nor (_21746_, _13460_, _09432_);
  nor (_21747_, _21746_, _21668_);
  nor (_21748_, _21747_, _04060_);
  or (_21749_, _21748_, _21745_);
  or (_21750_, _21749_, _43156_);
  or (_21751_, _43152_, \oc8051_golden_model_1.TH0 [6]);
  and (_21753_, _21751_, _41894_);
  and (_43453_, _21753_, _21750_);
  not (_21754_, \oc8051_golden_model_1.TH1 [0]);
  nor (_21755_, _05469_, _21754_);
  and (_21756_, _05716_, _05469_);
  nor (_21757_, _21756_, _21755_);
  and (_21758_, _21757_, _17157_);
  and (_21759_, _06962_, _05469_);
  nor (_21760_, _21755_, _03738_);
  not (_21761_, _21760_);
  nor (_21763_, _21761_, _21759_);
  and (_21764_, _05469_, _04700_);
  nor (_21765_, _21764_, _21755_);
  and (_21766_, _21765_, _08474_);
  and (_21767_, _05469_, \oc8051_golden_model_1.ACC [0]);
  nor (_21768_, _21767_, _21755_);
  nor (_21769_, _21768_, _04708_);
  nor (_21770_, _04707_, _21754_);
  or (_21771_, _21770_, _21769_);
  and (_21772_, _21771_, _04722_);
  nor (_21774_, _21757_, _04722_);
  or (_21775_, _21774_, _21772_);
  and (_21776_, _21775_, _04733_);
  nor (_21777_, _21765_, _04733_);
  nor (_21778_, _21777_, _21776_);
  nor (_21779_, _21778_, _03854_);
  nor (_21780_, _21768_, _03855_);
  or (_21781_, _21780_, _07927_);
  nor (_21782_, _21781_, _21779_);
  nor (_21783_, _21782_, _21766_);
  not (_21785_, _21783_);
  nor (_21786_, _21785_, _21763_);
  and (_21787_, _21786_, _03820_);
  nor (_21788_, _12164_, _09514_);
  nor (_21789_, _21788_, _21755_);
  nor (_21790_, _21789_, _03820_);
  or (_21791_, _21790_, _21787_);
  and (_21792_, _21791_, _04778_);
  and (_21793_, _05469_, _06479_);
  nor (_21794_, _21793_, _21755_);
  nor (_21796_, _21794_, _04778_);
  or (_21797_, _21796_, _21792_);
  and (_21798_, _21797_, _04790_);
  and (_21799_, _12178_, _05469_);
  nor (_21800_, _21799_, _21755_);
  nor (_21801_, _21800_, _04790_);
  or (_21802_, _21801_, _21798_);
  and (_21803_, _21802_, _04792_);
  nor (_21804_, _10488_, _09514_);
  nor (_21805_, _21804_, _21755_);
  not (_21807_, _21805_);
  and (_21808_, _08753_, _05469_);
  nor (_21809_, _21808_, _04792_);
  and (_21810_, _21809_, _21807_);
  nor (_21811_, _21810_, _21803_);
  nor (_21812_, _21811_, _03908_);
  and (_21813_, _12058_, _05469_);
  or (_21814_, _21813_, _21755_);
  and (_21815_, _21814_, _03908_);
  or (_21816_, _21815_, _21812_);
  and (_21818_, _21816_, _04785_);
  nor (_21819_, _21808_, _21755_);
  nor (_21820_, _21819_, _04785_);
  or (_21821_, _21820_, _21818_);
  and (_21822_, _21821_, _06567_);
  nor (_21823_, _12177_, _09514_);
  nor (_21824_, _21823_, _21755_);
  nor (_21825_, _21824_, _06567_);
  or (_21826_, _21825_, _21822_);
  and (_21827_, _21826_, _06572_);
  nor (_21829_, _21805_, _06572_);
  nor (_21830_, _21829_, _17157_);
  not (_21831_, _21830_);
  nor (_21832_, _21831_, _21827_);
  nor (_21833_, _21832_, _21758_);
  or (_21834_, _21833_, _43156_);
  or (_21835_, _43152_, \oc8051_golden_model_1.TH1 [0]);
  and (_21836_, _21835_, _41894_);
  and (_43455_, _21836_, _21834_);
  and (_21837_, _05469_, _04595_);
  not (_21839_, _21837_);
  nor (_21840_, _05469_, \oc8051_golden_model_1.TH1 [1]);
  nor (_21841_, _21840_, _04778_);
  and (_21842_, _21841_, _21839_);
  and (_21843_, _06961_, _05469_);
  not (_21844_, \oc8051_golden_model_1.TH1 [1]);
  nor (_21845_, _05469_, _21844_);
  nor (_21846_, _21845_, _03738_);
  not (_21847_, _21846_);
  nor (_21848_, _21847_, _21843_);
  not (_21850_, _21848_);
  and (_21851_, _05469_, \oc8051_golden_model_1.ACC [1]);
  nor (_21852_, _21851_, _21845_);
  nor (_21853_, _21852_, _04708_);
  nor (_21854_, _04707_, _21844_);
  or (_21855_, _21854_, _21853_);
  and (_21856_, _21855_, _04722_);
  and (_21857_, _12262_, _05469_);
  nor (_21858_, _21857_, _21840_);
  and (_21859_, _21858_, _03850_);
  or (_21861_, _21859_, _21856_);
  and (_21862_, _21861_, _04733_);
  and (_21863_, _05469_, _04900_);
  nor (_21864_, _21863_, _21845_);
  nor (_21865_, _21864_, _04733_);
  nor (_21866_, _21865_, _21862_);
  nor (_21867_, _21866_, _03854_);
  nor (_21868_, _21852_, _03855_);
  or (_21869_, _21868_, _07927_);
  or (_21870_, _21869_, _21867_);
  and (_21872_, _21864_, _08474_);
  nor (_21873_, _21872_, _03455_);
  and (_21874_, _21873_, _21870_);
  and (_21875_, _21874_, _21850_);
  not (_21876_, _21840_);
  and (_21877_, _12352_, _05469_);
  nor (_21878_, _21877_, _03820_);
  and (_21879_, _21878_, _21876_);
  nor (_21880_, _21879_, _21875_);
  nor (_21881_, _21880_, _03903_);
  nor (_21883_, _21881_, _21842_);
  nor (_21884_, _21883_, _03897_);
  nor (_21885_, _12366_, _09514_);
  nor (_21886_, _21885_, _04790_);
  and (_21887_, _21886_, _21876_);
  nor (_21888_, _21887_, _21884_);
  nor (_21889_, _21888_, _04018_);
  nor (_21890_, _08751_, _09514_);
  nor (_21891_, _21890_, _21845_);
  and (_21892_, _08750_, _05469_);
  nor (_21894_, _21892_, _21891_);
  and (_21895_, _21894_, _04018_);
  or (_21896_, _21895_, _21889_);
  and (_21897_, _21896_, _03909_);
  and (_21898_, _12244_, _05469_);
  or (_21899_, _21898_, _21845_);
  and (_21900_, _21899_, _03908_);
  or (_21901_, _21900_, _21897_);
  and (_21902_, _21901_, _04785_);
  nor (_21903_, _21892_, _21845_);
  nor (_21905_, _21903_, _04785_);
  or (_21906_, _21905_, _21902_);
  and (_21907_, _21906_, _06567_);
  and (_21908_, _21837_, _05669_);
  nor (_21909_, _21908_, _06567_);
  and (_21910_, _21909_, _21876_);
  or (_21911_, _21910_, _21907_);
  and (_21912_, _21911_, _06572_);
  nor (_21913_, _21891_, _06572_);
  or (_21914_, _21913_, _21912_);
  nor (_21916_, _21914_, _03773_);
  nor (_21917_, _21858_, _03774_);
  or (_21918_, _21917_, _03772_);
  nor (_21919_, _21918_, _21916_);
  nor (_21920_, _21857_, _21845_);
  nor (_21921_, _21920_, _04060_);
  or (_21922_, _21921_, _21919_);
  or (_21923_, _21922_, _43156_);
  or (_21924_, _43152_, \oc8051_golden_model_1.TH1 [1]);
  and (_21925_, _21924_, _41894_);
  and (_43456_, _21925_, _21923_);
  and (_21927_, _06965_, _05469_);
  not (_21928_, \oc8051_golden_model_1.TH1 [2]);
  nor (_21929_, _05469_, _21928_);
  nor (_21930_, _21929_, _03738_);
  not (_21931_, _21930_);
  nor (_21932_, _21931_, _21927_);
  and (_21933_, _05469_, \oc8051_golden_model_1.ACC [2]);
  nor (_21934_, _21933_, _21929_);
  nor (_21935_, _21934_, _04708_);
  nor (_21937_, _04707_, _21928_);
  or (_21938_, _21937_, _21935_);
  and (_21939_, _21938_, _04722_);
  nor (_21940_, _12471_, _09514_);
  nor (_21941_, _21940_, _21929_);
  nor (_21942_, _21941_, _04722_);
  or (_21943_, _21942_, _21939_);
  and (_21944_, _21943_, _04733_);
  and (_21945_, _05469_, _05307_);
  nor (_21946_, _21945_, _21929_);
  nor (_21947_, _21946_, _04733_);
  nor (_21948_, _21947_, _21944_);
  nor (_21949_, _21948_, _03854_);
  nor (_21950_, _21934_, _03855_);
  or (_21951_, _21950_, _07927_);
  nor (_21952_, _21951_, _21949_);
  and (_21953_, _21946_, _08474_);
  or (_21954_, _21953_, _03455_);
  or (_21955_, _21954_, _21952_);
  nor (_21956_, _21955_, _21932_);
  nor (_21959_, _12572_, _09514_);
  nor (_21960_, _21959_, _21929_);
  nor (_21961_, _21960_, _03820_);
  or (_21962_, _21961_, _21956_);
  and (_21963_, _21962_, _04778_);
  and (_21964_, _05469_, _06495_);
  nor (_21965_, _21964_, _21929_);
  nor (_21966_, _21965_, _04778_);
  or (_21967_, _21966_, _21963_);
  nor (_21968_, _21967_, _03897_);
  and (_21970_, _12586_, _05469_);
  or (_21971_, _21929_, _04790_);
  nor (_21972_, _21971_, _21970_);
  or (_21973_, _21972_, _04018_);
  nor (_21974_, _21973_, _21968_);
  and (_21975_, _08748_, _05469_);
  nor (_21976_, _21975_, _21929_);
  nor (_21977_, _21976_, _04792_);
  nor (_21978_, _21977_, _21974_);
  nor (_21979_, _21978_, _03908_);
  nor (_21981_, _21929_, _05765_);
  not (_21982_, _21981_);
  nor (_21983_, _21965_, _03909_);
  and (_21984_, _21983_, _21982_);
  nor (_21985_, _21984_, _21979_);
  nor (_21986_, _21985_, _04027_);
  nor (_21987_, _21934_, _04785_);
  and (_21988_, _21987_, _21982_);
  nor (_21989_, _21988_, _03914_);
  not (_21990_, _21989_);
  nor (_21992_, _21990_, _21986_);
  nor (_21993_, _12585_, _09514_);
  or (_21994_, _21929_, _06567_);
  nor (_21995_, _21994_, _21993_);
  or (_21996_, _21995_, _04011_);
  nor (_21997_, _21996_, _21992_);
  nor (_21998_, _08747_, _09514_);
  nor (_21999_, _21998_, _21929_);
  nor (_22000_, _21999_, _06572_);
  or (_22001_, _22000_, _03773_);
  nor (_22003_, _22001_, _21997_);
  and (_22004_, _21941_, _03773_);
  or (_22005_, _22004_, _03772_);
  nor (_22006_, _22005_, _22003_);
  and (_22007_, _12642_, _05469_);
  nor (_22008_, _22007_, _21929_);
  nor (_22009_, _22008_, _04060_);
  or (_22010_, _22009_, _22006_);
  or (_22011_, _22010_, _43156_);
  or (_22012_, _43152_, \oc8051_golden_model_1.TH1 [2]);
  and (_22014_, _22012_, _41894_);
  and (_43457_, _22014_, _22011_);
  not (_22015_, \oc8051_golden_model_1.TH1 [3]);
  nor (_22016_, _05469_, _22015_);
  and (_22017_, _05469_, \oc8051_golden_model_1.ACC [3]);
  nor (_22018_, _22017_, _22016_);
  nor (_22019_, _22018_, _04708_);
  nor (_22020_, _04707_, _22015_);
  or (_22021_, _22020_, _22019_);
  and (_22022_, _22021_, _04722_);
  nor (_22024_, _12681_, _09514_);
  nor (_22025_, _22024_, _22016_);
  nor (_22026_, _22025_, _04722_);
  or (_22027_, _22026_, _22022_);
  and (_22028_, _22027_, _04733_);
  and (_22029_, _05469_, _05119_);
  nor (_22030_, _22029_, _22016_);
  nor (_22031_, _22030_, _04733_);
  nor (_22032_, _22031_, _22028_);
  nor (_22033_, _22032_, _03854_);
  nor (_22035_, _22018_, _03855_);
  or (_22036_, _22035_, _07927_);
  or (_22037_, _22036_, _22033_);
  and (_22038_, _06964_, _05469_);
  nor (_22039_, _22016_, _03738_);
  not (_22040_, _22039_);
  nor (_22041_, _22040_, _22038_);
  and (_22042_, _22030_, _08474_);
  or (_22043_, _22042_, _03455_);
  nor (_22044_, _22043_, _22041_);
  and (_22046_, _22044_, _22037_);
  nor (_22047_, _12775_, _09514_);
  nor (_22048_, _22047_, _22016_);
  nor (_22049_, _22048_, _03820_);
  or (_22050_, _22049_, _22046_);
  and (_22051_, _22050_, _04778_);
  and (_22052_, _05469_, _06345_);
  nor (_22053_, _22052_, _22016_);
  nor (_22054_, _22053_, _04778_);
  or (_22055_, _22054_, _22051_);
  and (_22057_, _22055_, _04790_);
  and (_22058_, _12789_, _05469_);
  nor (_22059_, _22058_, _22016_);
  nor (_22060_, _22059_, _04790_);
  or (_22061_, _22060_, _22057_);
  and (_22062_, _22061_, _04792_);
  and (_22063_, _10491_, _05469_);
  nor (_22064_, _22063_, _22016_);
  nor (_22065_, _22064_, _04792_);
  nor (_22066_, _22065_, _22062_);
  nor (_22068_, _22066_, _03908_);
  nor (_22069_, _22016_, _05622_);
  not (_22070_, _22069_);
  nor (_22071_, _22053_, _03909_);
  and (_22072_, _22071_, _22070_);
  nor (_22073_, _22072_, _22068_);
  nor (_22074_, _22073_, _04027_);
  nor (_22075_, _22018_, _04785_);
  and (_22076_, _22075_, _22070_);
  or (_22077_, _22076_, _22074_);
  and (_22079_, _22077_, _06567_);
  nor (_22080_, _12788_, _09514_);
  nor (_22081_, _22080_, _22016_);
  nor (_22082_, _22081_, _06567_);
  or (_22083_, _22082_, _22079_);
  and (_22084_, _22083_, _06572_);
  nor (_22085_, _08742_, _09514_);
  nor (_22086_, _22085_, _22016_);
  nor (_22087_, _22086_, _06572_);
  or (_22088_, _22087_, _03773_);
  nor (_22090_, _22088_, _22084_);
  and (_22091_, _22025_, _03773_);
  or (_22092_, _22091_, _03772_);
  nor (_22093_, _22092_, _22090_);
  and (_22094_, _12848_, _05469_);
  nor (_22095_, _22094_, _22016_);
  nor (_22096_, _22095_, _04060_);
  or (_22097_, _22096_, _22093_);
  or (_22098_, _22097_, _43156_);
  or (_22099_, _43152_, \oc8051_golden_model_1.TH1 [3]);
  and (_22101_, _22099_, _41894_);
  and (_43458_, _22101_, _22098_);
  not (_22102_, \oc8051_golden_model_1.TH1 [4]);
  nor (_22103_, _05469_, _22102_);
  and (_22104_, _05469_, \oc8051_golden_model_1.ACC [4]);
  nor (_22105_, _22104_, _22103_);
  nor (_22106_, _22105_, _04708_);
  nor (_22107_, _04707_, _22102_);
  or (_22108_, _22107_, _22106_);
  and (_22109_, _22108_, _04722_);
  nor (_22111_, _12891_, _09514_);
  nor (_22112_, _22111_, _22103_);
  nor (_22113_, _22112_, _04722_);
  or (_22114_, _22113_, _22109_);
  and (_22115_, _22114_, _04733_);
  and (_22116_, _05950_, _05469_);
  nor (_22117_, _22116_, _22103_);
  nor (_22118_, _22117_, _04733_);
  nor (_22119_, _22118_, _22115_);
  nor (_22120_, _22119_, _03854_);
  nor (_22122_, _22105_, _03855_);
  or (_22123_, _22122_, _07927_);
  or (_22124_, _22123_, _22120_);
  and (_22125_, _06969_, _05469_);
  nor (_22126_, _22103_, _03738_);
  not (_22127_, _22126_);
  nor (_22128_, _22127_, _22125_);
  and (_22129_, _22117_, _08474_);
  or (_22130_, _22129_, _03455_);
  nor (_22131_, _22130_, _22128_);
  and (_22133_, _22131_, _22124_);
  nor (_22134_, _12982_, _09514_);
  nor (_22135_, _22134_, _22103_);
  nor (_22136_, _22135_, _03820_);
  or (_22137_, _22136_, _22133_);
  and (_22138_, _22137_, _04778_);
  and (_22139_, _06456_, _05469_);
  nor (_22140_, _22139_, _22103_);
  nor (_22141_, _22140_, _04778_);
  or (_22142_, _22141_, _22138_);
  and (_22144_, _22142_, _04790_);
  and (_22145_, _12997_, _05469_);
  nor (_22146_, _22145_, _22103_);
  nor (_22147_, _22146_, _04790_);
  or (_22148_, _22147_, _22144_);
  and (_22149_, _22148_, _04792_);
  and (_22150_, _08741_, _05469_);
  nor (_22151_, _22150_, _22103_);
  nor (_22152_, _22151_, _04792_);
  nor (_22153_, _22152_, _22149_);
  nor (_22155_, _22153_, _03908_);
  nor (_22156_, _22103_, _08336_);
  not (_22157_, _22156_);
  nor (_22158_, _22140_, _03909_);
  and (_22159_, _22158_, _22157_);
  nor (_22160_, _22159_, _22155_);
  nor (_22161_, _22160_, _04027_);
  nor (_22162_, _22105_, _04785_);
  and (_22163_, _22162_, _22157_);
  nor (_22164_, _22163_, _03914_);
  not (_22166_, _22164_);
  nor (_22167_, _22166_, _22161_);
  nor (_22168_, _12996_, _09514_);
  or (_22169_, _22103_, _06567_);
  nor (_22170_, _22169_, _22168_);
  or (_22171_, _22170_, _04011_);
  nor (_22172_, _22171_, _22167_);
  nor (_22173_, _08740_, _09514_);
  nor (_22174_, _22173_, _22103_);
  nor (_22175_, _22174_, _06572_);
  or (_22177_, _22175_, _03773_);
  nor (_22178_, _22177_, _22172_);
  and (_22179_, _22112_, _03773_);
  or (_22180_, _22179_, _03772_);
  nor (_22181_, _22180_, _22178_);
  and (_22182_, _13056_, _05469_);
  nor (_22183_, _22182_, _22103_);
  nor (_22184_, _22183_, _04060_);
  or (_22185_, _22184_, _22181_);
  or (_22186_, _22185_, _43156_);
  or (_22188_, _43152_, \oc8051_golden_model_1.TH1 [4]);
  and (_22189_, _22188_, _41894_);
  and (_43459_, _22189_, _22186_);
  not (_22190_, \oc8051_golden_model_1.TH1 [5]);
  nor (_22191_, _05469_, _22190_);
  and (_22192_, _05469_, \oc8051_golden_model_1.ACC [5]);
  nor (_22193_, _22192_, _22191_);
  nor (_22194_, _22193_, _04708_);
  nor (_22195_, _04707_, _22190_);
  or (_22196_, _22195_, _22194_);
  and (_22198_, _22196_, _04722_);
  nor (_22199_, _13090_, _09514_);
  nor (_22200_, _22199_, _22191_);
  nor (_22201_, _22200_, _04722_);
  or (_22202_, _22201_, _22198_);
  and (_22203_, _22202_, _04733_);
  and (_22204_, _05857_, _05469_);
  nor (_22205_, _22204_, _22191_);
  nor (_22206_, _22205_, _04733_);
  nor (_22207_, _22206_, _22203_);
  nor (_22209_, _22207_, _03854_);
  nor (_22210_, _22193_, _03855_);
  or (_22211_, _22210_, _07927_);
  or (_22212_, _22211_, _22209_);
  and (_22213_, _06968_, _05469_);
  nor (_22214_, _22191_, _03738_);
  not (_22215_, _22214_);
  nor (_22216_, _22215_, _22213_);
  and (_22217_, _22205_, _08474_);
  or (_22218_, _22217_, _03455_);
  nor (_22221_, _22218_, _22216_);
  and (_22222_, _22221_, _22212_);
  nor (_22223_, _13182_, _09514_);
  nor (_22224_, _22223_, _22191_);
  nor (_22225_, _22224_, _03820_);
  or (_22226_, _22225_, _22222_);
  and (_22227_, _22226_, _04778_);
  and (_22228_, _06447_, _05469_);
  nor (_22229_, _22228_, _22191_);
  nor (_22230_, _22229_, _04778_);
  or (_22232_, _22230_, _22227_);
  and (_22233_, _22232_, _04790_);
  and (_22234_, _13196_, _05469_);
  nor (_22235_, _22234_, _22191_);
  nor (_22236_, _22235_, _04790_);
  or (_22237_, _22236_, _22233_);
  and (_22238_, _22237_, _04792_);
  and (_22239_, _10493_, _05469_);
  nor (_22240_, _22239_, _22191_);
  nor (_22241_, _22240_, _04792_);
  nor (_22243_, _22241_, _22238_);
  nor (_22244_, _22243_, _03908_);
  nor (_22245_, _22191_, _08335_);
  not (_22246_, _22245_);
  nor (_22247_, _22229_, _03909_);
  and (_22248_, _22247_, _22246_);
  nor (_22249_, _22248_, _22244_);
  nor (_22250_, _22249_, _04027_);
  nor (_22251_, _22193_, _04785_);
  and (_22252_, _22251_, _22246_);
  or (_22254_, _22252_, _22250_);
  and (_22255_, _22254_, _06567_);
  nor (_22256_, _13195_, _09514_);
  nor (_22257_, _22256_, _22191_);
  nor (_22258_, _22257_, _06567_);
  or (_22259_, _22258_, _22255_);
  and (_22260_, _22259_, _06572_);
  nor (_22261_, _08738_, _09514_);
  nor (_22262_, _22261_, _22191_);
  nor (_22263_, _22262_, _06572_);
  nor (_22265_, _22263_, _22260_);
  nor (_22266_, _22265_, _03773_);
  nor (_22267_, _22200_, _03774_);
  or (_22268_, _22267_, _03772_);
  nor (_22269_, _22268_, _22266_);
  and (_22270_, _13255_, _05469_);
  nor (_22271_, _22270_, _22191_);
  and (_22272_, _22271_, _03772_);
  nor (_22273_, _22272_, _22269_);
  or (_22274_, _22273_, _43156_);
  or (_22276_, _43152_, \oc8051_golden_model_1.TH1 [5]);
  and (_22277_, _22276_, _41894_);
  and (_43460_, _22277_, _22274_);
  not (_22278_, \oc8051_golden_model_1.TH1 [6]);
  nor (_22279_, _05469_, _22278_);
  and (_22280_, _05469_, \oc8051_golden_model_1.ACC [6]);
  nor (_22281_, _22280_, _22279_);
  nor (_22282_, _22281_, _04708_);
  nor (_22283_, _04707_, _22278_);
  or (_22284_, _22283_, _22282_);
  and (_22286_, _22284_, _04722_);
  nor (_22287_, _13293_, _09514_);
  nor (_22288_, _22287_, _22279_);
  nor (_22289_, _22288_, _04722_);
  or (_22290_, _22289_, _22286_);
  and (_22291_, _22290_, _04733_);
  and (_22292_, _06065_, _05469_);
  nor (_22293_, _22292_, _22279_);
  nor (_22294_, _22293_, _04733_);
  nor (_22295_, _22294_, _22291_);
  nor (_22297_, _22295_, _03854_);
  nor (_22298_, _22281_, _03855_);
  or (_22299_, _22298_, _07927_);
  or (_22300_, _22299_, _22297_);
  and (_22301_, _06641_, _05469_);
  nor (_22302_, _22279_, _03738_);
  not (_22303_, _22302_);
  nor (_22304_, _22303_, _22301_);
  and (_22305_, _22293_, _08474_);
  or (_22306_, _22305_, _03455_);
  nor (_22308_, _22306_, _22304_);
  and (_22309_, _22308_, _22300_);
  nor (_22310_, _13387_, _09514_);
  nor (_22311_, _22310_, _22279_);
  nor (_22312_, _22311_, _03820_);
  or (_22313_, _22312_, _22309_);
  and (_22314_, _22313_, _04778_);
  and (_22315_, _13394_, _05469_);
  nor (_22316_, _22315_, _22279_);
  nor (_22317_, _22316_, _04778_);
  or (_22319_, _22317_, _22314_);
  nor (_22320_, _22319_, _03897_);
  and (_22321_, _13402_, _05469_);
  or (_22322_, _22279_, _04790_);
  nor (_22323_, _22322_, _22321_);
  or (_22324_, _22323_, _04018_);
  nor (_22325_, _22324_, _22320_);
  and (_22326_, _08736_, _05469_);
  nor (_22327_, _22326_, _22279_);
  nor (_22328_, _22327_, _04792_);
  nor (_22331_, _22328_, _22325_);
  nor (_22332_, _22331_, _03908_);
  nor (_22333_, _22279_, _08322_);
  not (_22334_, _22333_);
  nor (_22335_, _22316_, _03909_);
  and (_22336_, _22335_, _22334_);
  nor (_22337_, _22336_, _22332_);
  nor (_22338_, _22337_, _04027_);
  nor (_22339_, _22281_, _04785_);
  and (_22340_, _22339_, _22334_);
  or (_22342_, _22340_, _22338_);
  and (_22343_, _22342_, _06567_);
  nor (_22344_, _13401_, _09514_);
  nor (_22345_, _22344_, _22279_);
  nor (_22346_, _22345_, _06567_);
  or (_22347_, _22346_, _22343_);
  and (_22348_, _22347_, _06572_);
  nor (_22349_, _08735_, _09514_);
  nor (_22350_, _22349_, _22279_);
  nor (_22351_, _22350_, _06572_);
  or (_22353_, _22351_, _03773_);
  nor (_22354_, _22353_, _22348_);
  and (_22355_, _22288_, _03773_);
  or (_22356_, _22355_, _03772_);
  nor (_22357_, _22356_, _22354_);
  nor (_22358_, _13460_, _09514_);
  nor (_22359_, _22358_, _22279_);
  nor (_22360_, _22359_, _04060_);
  or (_22361_, _22360_, _22357_);
  or (_22362_, _22361_, _43156_);
  or (_22364_, _43152_, \oc8051_golden_model_1.TH1 [6]);
  and (_22365_, _22364_, _41894_);
  and (_43461_, _22365_, _22362_);
  not (_22366_, \oc8051_golden_model_1.TMOD [0]);
  nor (_22367_, _05475_, _22366_);
  and (_22368_, _05716_, _05475_);
  nor (_22369_, _22368_, _22367_);
  and (_22370_, _22369_, _17157_);
  and (_22371_, _06962_, _05475_);
  nor (_22372_, _22367_, _03738_);
  not (_22374_, _22372_);
  nor (_22375_, _22374_, _22371_);
  and (_22376_, _05475_, _04700_);
  nor (_22377_, _22376_, _22367_);
  and (_22378_, _22377_, _08474_);
  nor (_22379_, _22369_, _04722_);
  nor (_22380_, _04707_, _22366_);
  and (_22381_, _05475_, \oc8051_golden_model_1.ACC [0]);
  nor (_22382_, _22381_, _22367_);
  nor (_22383_, _22382_, _04708_);
  nor (_22385_, _22383_, _22380_);
  nor (_22386_, _22385_, _03850_);
  or (_22387_, _22386_, _22379_);
  and (_22388_, _22387_, _04733_);
  nor (_22389_, _22377_, _04733_);
  or (_22390_, _22389_, _22388_);
  and (_22391_, _22390_, _03855_);
  nor (_22392_, _22382_, _03855_);
  or (_22393_, _22392_, _07927_);
  nor (_22394_, _22393_, _22391_);
  nor (_22396_, _22394_, _22378_);
  not (_22397_, _22396_);
  nor (_22398_, _22397_, _22375_);
  and (_22399_, _22398_, _03820_);
  nor (_22400_, _12164_, _09595_);
  nor (_22401_, _22400_, _22367_);
  nor (_22402_, _22401_, _03820_);
  or (_22403_, _22402_, _22399_);
  and (_22404_, _22403_, _04778_);
  and (_22405_, _05475_, _06479_);
  nor (_22407_, _22405_, _22367_);
  nor (_22408_, _22407_, _04778_);
  or (_22409_, _22408_, _22404_);
  and (_22410_, _22409_, _04790_);
  and (_22411_, _12178_, _05475_);
  nor (_22412_, _22411_, _22367_);
  nor (_22413_, _22412_, _04790_);
  or (_22414_, _22413_, _22410_);
  and (_22415_, _22414_, _04792_);
  nor (_22416_, _10488_, _09595_);
  nor (_22418_, _22416_, _22367_);
  not (_22419_, _22418_);
  and (_22420_, _08753_, _05475_);
  nor (_22421_, _22420_, _04792_);
  and (_22422_, _22421_, _22419_);
  nor (_22423_, _22422_, _22415_);
  nor (_22424_, _22423_, _03908_);
  and (_22425_, _12058_, _05475_);
  or (_22426_, _22425_, _22367_);
  and (_22427_, _22426_, _03908_);
  or (_22429_, _22427_, _22424_);
  and (_22430_, _22429_, _04785_);
  nor (_22431_, _22420_, _22367_);
  nor (_22432_, _22431_, _04785_);
  or (_22433_, _22432_, _22430_);
  and (_22434_, _22433_, _06567_);
  nor (_22435_, _12177_, _09595_);
  nor (_22436_, _22435_, _22367_);
  nor (_22437_, _22436_, _06567_);
  or (_22438_, _22437_, _22434_);
  and (_22440_, _22438_, _06572_);
  nor (_22441_, _22418_, _06572_);
  nor (_22442_, _22441_, _17157_);
  not (_22443_, _22442_);
  nor (_22444_, _22443_, _22440_);
  nor (_22445_, _22444_, _22370_);
  or (_22446_, _22445_, _43156_);
  or (_22447_, _43152_, \oc8051_golden_model_1.TMOD [0]);
  and (_22448_, _22447_, _41894_);
  and (_43464_, _22448_, _22446_);
  and (_22450_, _05475_, _04595_);
  not (_22451_, _22450_);
  nor (_22452_, _05475_, \oc8051_golden_model_1.TMOD [1]);
  nor (_22453_, _22452_, _04778_);
  and (_22454_, _22453_, _22451_);
  and (_22455_, _06961_, _05475_);
  not (_22456_, \oc8051_golden_model_1.TMOD [1]);
  nor (_22457_, _05475_, _22456_);
  nor (_22458_, _22457_, _03738_);
  not (_22459_, _22458_);
  nor (_22461_, _22459_, _22455_);
  not (_22462_, _22461_);
  and (_22463_, _05475_, \oc8051_golden_model_1.ACC [1]);
  nor (_22464_, _22463_, _22457_);
  nor (_22465_, _22464_, _04708_);
  nor (_22466_, _04707_, _22456_);
  or (_22467_, _22466_, _22465_);
  and (_22468_, _22467_, _04722_);
  and (_22469_, _12262_, _05475_);
  nor (_22470_, _22469_, _22452_);
  and (_22472_, _22470_, _03850_);
  or (_22473_, _22472_, _22468_);
  and (_22474_, _22473_, _04733_);
  and (_22475_, _05475_, _04900_);
  nor (_22476_, _22475_, _22457_);
  nor (_22477_, _22476_, _04733_);
  nor (_22478_, _22477_, _22474_);
  nor (_22479_, _22478_, _03854_);
  nor (_22480_, _22464_, _03855_);
  or (_22481_, _22480_, _07927_);
  or (_22483_, _22481_, _22479_);
  and (_22484_, _22476_, _08474_);
  nor (_22485_, _22484_, _03455_);
  and (_22486_, _22485_, _22483_);
  and (_22487_, _22486_, _22462_);
  and (_22488_, _12352_, _05475_);
  or (_22489_, _22488_, _03820_);
  nor (_22490_, _22489_, _22452_);
  nor (_22491_, _22490_, _22487_);
  nor (_22492_, _22491_, _03903_);
  nor (_22494_, _22492_, _22454_);
  nor (_22495_, _22494_, _03897_);
  and (_22496_, _12366_, _05475_);
  or (_22497_, _22496_, _22457_);
  and (_22498_, _22497_, _03897_);
  nor (_22499_, _22498_, _22495_);
  nor (_22500_, _22499_, _04018_);
  nor (_22501_, _08751_, _09595_);
  nor (_22502_, _22501_, _22457_);
  and (_22503_, _08750_, _05475_);
  nor (_22505_, _22503_, _22502_);
  and (_22506_, _22505_, _04018_);
  or (_22507_, _22506_, _22500_);
  and (_22508_, _22507_, _03909_);
  and (_22509_, _12244_, _05475_);
  or (_22510_, _22509_, _22457_);
  and (_22511_, _22510_, _03908_);
  or (_22512_, _22511_, _22508_);
  and (_22513_, _22512_, _04785_);
  nor (_22514_, _22503_, _22457_);
  nor (_22516_, _22514_, _04785_);
  or (_22517_, _22516_, _22513_);
  and (_22518_, _22517_, _06567_);
  nor (_22519_, _12365_, _09595_);
  or (_22520_, _22519_, _22457_);
  and (_22521_, _22520_, _03914_);
  or (_22522_, _22521_, _22518_);
  and (_22523_, _22522_, _06572_);
  nor (_22524_, _22502_, _06572_);
  or (_22525_, _22524_, _22523_);
  nor (_22527_, _22525_, _03773_);
  nor (_22528_, _22470_, _03774_);
  or (_22529_, _22528_, _03772_);
  nor (_22530_, _22529_, _22527_);
  nor (_22531_, _22469_, _22457_);
  nor (_22532_, _22531_, _04060_);
  or (_22533_, _22532_, _22530_);
  or (_22534_, _22533_, _43156_);
  or (_22535_, _43152_, \oc8051_golden_model_1.TMOD [1]);
  and (_22536_, _22535_, _41894_);
  and (_43465_, _22536_, _22534_);
  and (_22538_, _06965_, _05475_);
  not (_22539_, \oc8051_golden_model_1.TMOD [2]);
  nor (_22540_, _05475_, _22539_);
  nor (_22541_, _22540_, _03738_);
  not (_22542_, _22541_);
  nor (_22543_, _22542_, _22538_);
  and (_22544_, _05475_, \oc8051_golden_model_1.ACC [2]);
  nor (_22545_, _22544_, _22540_);
  nor (_22546_, _22545_, _04708_);
  nor (_22548_, _04707_, _22539_);
  or (_22549_, _22548_, _22546_);
  and (_22550_, _22549_, _04722_);
  nor (_22551_, _12471_, _09595_);
  nor (_22552_, _22551_, _22540_);
  nor (_22553_, _22552_, _04722_);
  or (_22554_, _22553_, _22550_);
  and (_22555_, _22554_, _04733_);
  and (_22556_, _05475_, _05307_);
  nor (_22557_, _22556_, _22540_);
  nor (_22559_, _22557_, _04733_);
  nor (_22560_, _22559_, _22555_);
  nor (_22561_, _22560_, _03854_);
  nor (_22562_, _22545_, _03855_);
  or (_22563_, _22562_, _07927_);
  nor (_22564_, _22563_, _22561_);
  and (_22565_, _22557_, _08474_);
  or (_22566_, _22565_, _03455_);
  or (_22567_, _22566_, _22564_);
  nor (_22568_, _22567_, _22543_);
  nor (_22570_, _12572_, _09595_);
  nor (_22571_, _22570_, _22540_);
  nor (_22572_, _22571_, _03820_);
  or (_22573_, _22572_, _22568_);
  and (_22574_, _22573_, _04778_);
  and (_22575_, _05475_, _06495_);
  nor (_22576_, _22575_, _22540_);
  nor (_22577_, _22576_, _04778_);
  or (_22578_, _22577_, _22574_);
  nor (_22579_, _22578_, _03897_);
  and (_22581_, _12586_, _05475_);
  or (_22582_, _22540_, _04790_);
  nor (_22583_, _22582_, _22581_);
  or (_22584_, _22583_, _04018_);
  nor (_22585_, _22584_, _22579_);
  and (_22586_, _08748_, _05475_);
  nor (_22587_, _22586_, _22540_);
  nor (_22588_, _22587_, _04792_);
  nor (_22589_, _22588_, _22585_);
  nor (_22590_, _22589_, _03908_);
  nor (_22592_, _22540_, _05765_);
  not (_22593_, _22592_);
  nor (_22594_, _22576_, _03909_);
  and (_22595_, _22594_, _22593_);
  nor (_22596_, _22595_, _22590_);
  nor (_22597_, _22596_, _04027_);
  nor (_22598_, _22545_, _04785_);
  and (_22599_, _22598_, _22593_);
  or (_22600_, _22599_, _22597_);
  and (_22601_, _22600_, _06567_);
  nor (_22603_, _12585_, _09595_);
  nor (_22604_, _22603_, _22540_);
  nor (_22605_, _22604_, _06567_);
  or (_22606_, _22605_, _22601_);
  and (_22607_, _22606_, _06572_);
  nor (_22608_, _08747_, _09595_);
  nor (_22609_, _22608_, _22540_);
  nor (_22610_, _22609_, _06572_);
  or (_22611_, _22610_, _03773_);
  nor (_22612_, _22611_, _22607_);
  and (_22614_, _22552_, _03773_);
  or (_22615_, _22614_, _03772_);
  nor (_22616_, _22615_, _22612_);
  and (_22617_, _12642_, _05475_);
  nor (_22618_, _22617_, _22540_);
  nor (_22619_, _22618_, _04060_);
  or (_22620_, _22619_, _22616_);
  or (_22621_, _22620_, _43156_);
  or (_22622_, _43152_, \oc8051_golden_model_1.TMOD [2]);
  and (_22623_, _22622_, _41894_);
  and (_43466_, _22623_, _22621_);
  not (_22625_, \oc8051_golden_model_1.TMOD [3]);
  nor (_22626_, _05475_, _22625_);
  and (_22627_, _05475_, \oc8051_golden_model_1.ACC [3]);
  nor (_22628_, _22627_, _22626_);
  nor (_22629_, _22628_, _04708_);
  nor (_22630_, _04707_, _22625_);
  or (_22631_, _22630_, _22629_);
  and (_22632_, _22631_, _04722_);
  nor (_22633_, _12681_, _09595_);
  nor (_22635_, _22633_, _22626_);
  nor (_22636_, _22635_, _04722_);
  or (_22637_, _22636_, _22632_);
  and (_22638_, _22637_, _04733_);
  and (_22639_, _05475_, _05119_);
  nor (_22640_, _22639_, _22626_);
  nor (_22641_, _22640_, _04733_);
  nor (_22642_, _22641_, _22638_);
  nor (_22643_, _22642_, _03854_);
  nor (_22644_, _22628_, _03855_);
  or (_22646_, _22644_, _07927_);
  or (_22647_, _22646_, _22643_);
  and (_22648_, _06964_, _05475_);
  nor (_22649_, _22626_, _03738_);
  not (_22650_, _22649_);
  nor (_22651_, _22650_, _22648_);
  and (_22652_, _22640_, _08474_);
  or (_22653_, _22652_, _03455_);
  nor (_22654_, _22653_, _22651_);
  and (_22655_, _22654_, _22647_);
  nor (_22657_, _12775_, _09595_);
  nor (_22658_, _22657_, _22626_);
  nor (_22659_, _22658_, _03820_);
  or (_22660_, _22659_, _22655_);
  and (_22661_, _22660_, _04778_);
  and (_22662_, _05475_, _06345_);
  nor (_22663_, _22662_, _22626_);
  nor (_22664_, _22663_, _04778_);
  or (_22665_, _22664_, _22661_);
  and (_22666_, _22665_, _04790_);
  and (_22668_, _12789_, _05475_);
  nor (_22669_, _22668_, _22626_);
  nor (_22670_, _22669_, _04790_);
  or (_22671_, _22670_, _22666_);
  and (_22672_, _22671_, _04792_);
  and (_22673_, _10491_, _05475_);
  nor (_22674_, _22673_, _22626_);
  nor (_22675_, _22674_, _04792_);
  nor (_22676_, _22675_, _22672_);
  nor (_22677_, _22676_, _03908_);
  nor (_22679_, _22626_, _05622_);
  not (_22680_, _22679_);
  nor (_22681_, _22663_, _03909_);
  and (_22682_, _22681_, _22680_);
  nor (_22683_, _22682_, _22677_);
  nor (_22684_, _22683_, _04027_);
  nor (_22685_, _22628_, _04785_);
  and (_22686_, _22685_, _22680_);
  or (_22687_, _22686_, _22684_);
  and (_22688_, _22687_, _06567_);
  nor (_22690_, _12788_, _09595_);
  nor (_22691_, _22690_, _22626_);
  nor (_22692_, _22691_, _06567_);
  or (_22693_, _22692_, _22688_);
  and (_22694_, _22693_, _06572_);
  nor (_22695_, _08742_, _09595_);
  nor (_22696_, _22695_, _22626_);
  nor (_22697_, _22696_, _06572_);
  or (_22698_, _22697_, _03773_);
  nor (_22699_, _22698_, _22694_);
  and (_22701_, _22635_, _03773_);
  or (_22702_, _22701_, _03772_);
  nor (_22703_, _22702_, _22699_);
  and (_22704_, _12848_, _05475_);
  nor (_22705_, _22704_, _22626_);
  nor (_22706_, _22705_, _04060_);
  or (_22707_, _22706_, _22703_);
  or (_22708_, _22707_, _43156_);
  or (_22709_, _43152_, \oc8051_golden_model_1.TMOD [3]);
  and (_22710_, _22709_, _41894_);
  and (_43467_, _22710_, _22708_);
  not (_22712_, \oc8051_golden_model_1.TMOD [4]);
  nor (_22713_, _05475_, _22712_);
  and (_22714_, _05475_, \oc8051_golden_model_1.ACC [4]);
  nor (_22715_, _22714_, _22713_);
  nor (_22716_, _22715_, _04708_);
  nor (_22717_, _04707_, _22712_);
  or (_22718_, _22717_, _22716_);
  and (_22719_, _22718_, _04722_);
  nor (_22720_, _12891_, _09595_);
  nor (_22722_, _22720_, _22713_);
  nor (_22723_, _22722_, _04722_);
  or (_22724_, _22723_, _22719_);
  and (_22725_, _22724_, _04733_);
  and (_22726_, _05950_, _05475_);
  nor (_22727_, _22726_, _22713_);
  nor (_22728_, _22727_, _04733_);
  nor (_22729_, _22728_, _22725_);
  nor (_22730_, _22729_, _03854_);
  nor (_22731_, _22715_, _03855_);
  or (_22733_, _22731_, _07927_);
  or (_22734_, _22733_, _22730_);
  and (_22735_, _06969_, _05475_);
  nor (_22736_, _22713_, _03738_);
  not (_22737_, _22736_);
  nor (_22738_, _22737_, _22735_);
  and (_22739_, _22727_, _08474_);
  or (_22740_, _22739_, _03455_);
  nor (_22741_, _22740_, _22738_);
  and (_22742_, _22741_, _22734_);
  nor (_22744_, _12982_, _09595_);
  nor (_22745_, _22744_, _22713_);
  nor (_22746_, _22745_, _03820_);
  or (_22747_, _22746_, _22742_);
  and (_22748_, _22747_, _04778_);
  and (_22749_, _06456_, _05475_);
  nor (_22750_, _22749_, _22713_);
  nor (_22751_, _22750_, _04778_);
  or (_22752_, _22751_, _22748_);
  nor (_22753_, _22752_, _03897_);
  and (_22755_, _12997_, _05475_);
  or (_22756_, _22713_, _04790_);
  nor (_22757_, _22756_, _22755_);
  or (_22758_, _22757_, _04018_);
  nor (_22759_, _22758_, _22753_);
  and (_22760_, _08741_, _05475_);
  nor (_22761_, _22760_, _22713_);
  nor (_22762_, _22761_, _04792_);
  nor (_22763_, _22762_, _22759_);
  nor (_22764_, _22763_, _03908_);
  nor (_22766_, _22713_, _08336_);
  not (_22767_, _22766_);
  nor (_22768_, _22750_, _03909_);
  and (_22769_, _22768_, _22767_);
  nor (_22770_, _22769_, _22764_);
  nor (_22771_, _22770_, _04027_);
  nor (_22772_, _22715_, _04785_);
  and (_22773_, _22772_, _22767_);
  or (_22774_, _22773_, _22771_);
  and (_22775_, _22774_, _06567_);
  nor (_22777_, _12996_, _09595_);
  nor (_22778_, _22777_, _22713_);
  nor (_22779_, _22778_, _06567_);
  or (_22780_, _22779_, _22775_);
  and (_22781_, _22780_, _06572_);
  nor (_22782_, _08740_, _09595_);
  nor (_22783_, _22782_, _22713_);
  nor (_22784_, _22783_, _06572_);
  or (_22785_, _22784_, _03773_);
  nor (_22786_, _22785_, _22781_);
  and (_22788_, _22722_, _03773_);
  or (_22789_, _22788_, _03772_);
  nor (_22790_, _22789_, _22786_);
  and (_22791_, _13056_, _05475_);
  nor (_22792_, _22791_, _22713_);
  nor (_22793_, _22792_, _04060_);
  or (_22794_, _22793_, _22790_);
  or (_22795_, _22794_, _43156_);
  or (_22796_, _43152_, \oc8051_golden_model_1.TMOD [4]);
  and (_22797_, _22796_, _41894_);
  and (_43468_, _22797_, _22795_);
  not (_22799_, \oc8051_golden_model_1.TMOD [5]);
  nor (_22800_, _05475_, _22799_);
  nor (_22801_, _13090_, _09595_);
  nor (_22802_, _22801_, _22800_);
  nor (_22803_, _22802_, _04722_);
  nor (_22804_, _04707_, _22799_);
  and (_22805_, _05475_, \oc8051_golden_model_1.ACC [5]);
  nor (_22806_, _22805_, _22800_);
  nor (_22807_, _22806_, _04708_);
  nor (_22809_, _22807_, _22804_);
  nor (_22810_, _22809_, _03850_);
  or (_22811_, _22810_, _22803_);
  and (_22812_, _22811_, _04733_);
  and (_22813_, _05857_, _05475_);
  nor (_22814_, _22813_, _22800_);
  nor (_22815_, _22814_, _04733_);
  or (_22816_, _22815_, _22812_);
  and (_22817_, _22816_, _03855_);
  nor (_22818_, _22806_, _03855_);
  or (_22820_, _22818_, _07927_);
  or (_22821_, _22820_, _22817_);
  and (_22822_, _06968_, _05475_);
  nor (_22823_, _22800_, _03738_);
  not (_22824_, _22823_);
  nor (_22825_, _22824_, _22822_);
  and (_22826_, _22814_, _08474_);
  or (_22827_, _22826_, _03455_);
  nor (_22828_, _22827_, _22825_);
  and (_22829_, _22828_, _22821_);
  nor (_22831_, _13182_, _09595_);
  nor (_22832_, _22831_, _22800_);
  nor (_22833_, _22832_, _03820_);
  or (_22834_, _22833_, _22829_);
  and (_22835_, _22834_, _04778_);
  and (_22836_, _06447_, _05475_);
  nor (_22837_, _22836_, _22800_);
  nor (_22838_, _22837_, _04778_);
  or (_22839_, _22838_, _22835_);
  and (_22840_, _22839_, _04790_);
  and (_22842_, _13196_, _05475_);
  nor (_22843_, _22842_, _22800_);
  nor (_22844_, _22843_, _04790_);
  or (_22845_, _22844_, _22840_);
  and (_22846_, _22845_, _04792_);
  and (_22847_, _10493_, _05475_);
  nor (_22848_, _22847_, _22800_);
  nor (_22849_, _22848_, _04792_);
  nor (_22850_, _22849_, _22846_);
  nor (_22851_, _22850_, _03908_);
  nor (_22853_, _22800_, _08335_);
  not (_22854_, _22853_);
  nor (_22855_, _22837_, _03909_);
  and (_22856_, _22855_, _22854_);
  nor (_22857_, _22856_, _22851_);
  nor (_22858_, _22857_, _04027_);
  nor (_22859_, _22806_, _04785_);
  and (_22860_, _22859_, _22854_);
  nor (_22861_, _22860_, _03914_);
  not (_22862_, _22861_);
  nor (_22864_, _22862_, _22858_);
  nor (_22865_, _13195_, _09595_);
  or (_22866_, _22800_, _06567_);
  nor (_22867_, _22866_, _22865_);
  or (_22868_, _22867_, _04011_);
  nor (_22869_, _22868_, _22864_);
  nor (_22870_, _08738_, _09595_);
  nor (_22871_, _22870_, _22800_);
  nor (_22872_, _22871_, _06572_);
  nor (_22873_, _22872_, _22869_);
  nor (_22875_, _22873_, _03773_);
  nor (_22876_, _22802_, _03774_);
  or (_22877_, _22876_, _03772_);
  nor (_22878_, _22877_, _22875_);
  and (_22879_, _13255_, _05475_);
  nor (_22880_, _22879_, _22800_);
  and (_22881_, _22880_, _03772_);
  nor (_22882_, _22881_, _22878_);
  or (_22883_, _22882_, _43156_);
  or (_22884_, _43152_, \oc8051_golden_model_1.TMOD [5]);
  and (_22885_, _22884_, _41894_);
  and (_43469_, _22885_, _22883_);
  not (_22886_, \oc8051_golden_model_1.TMOD [6]);
  nor (_22887_, _05475_, _22886_);
  and (_22888_, _05475_, \oc8051_golden_model_1.ACC [6]);
  nor (_22889_, _22888_, _22887_);
  nor (_22890_, _22889_, _04708_);
  nor (_22891_, _04707_, _22886_);
  or (_22892_, _22891_, _22890_);
  and (_22893_, _22892_, _04722_);
  nor (_22896_, _13293_, _09595_);
  nor (_22897_, _22896_, _22887_);
  nor (_22898_, _22897_, _04722_);
  or (_22899_, _22898_, _22893_);
  and (_22900_, _22899_, _04733_);
  and (_22901_, _06065_, _05475_);
  nor (_22902_, _22901_, _22887_);
  nor (_22903_, _22902_, _04733_);
  nor (_22904_, _22903_, _22900_);
  nor (_22905_, _22904_, _03854_);
  nor (_22907_, _22889_, _03855_);
  or (_22908_, _22907_, _07927_);
  or (_22909_, _22908_, _22905_);
  and (_22910_, _06641_, _05475_);
  nor (_22911_, _22887_, _03738_);
  not (_22912_, _22911_);
  nor (_22913_, _22912_, _22910_);
  and (_22914_, _22902_, _08474_);
  or (_22915_, _22914_, _03455_);
  nor (_22916_, _22915_, _22913_);
  and (_22917_, _22916_, _22909_);
  nor (_22918_, _13387_, _09595_);
  nor (_22919_, _22918_, _22887_);
  nor (_22920_, _22919_, _03820_);
  or (_22921_, _22920_, _22917_);
  and (_22922_, _22921_, _04778_);
  and (_22923_, _13394_, _05475_);
  nor (_22924_, _22923_, _22887_);
  nor (_22925_, _22924_, _04778_);
  or (_22926_, _22925_, _22922_);
  nor (_22929_, _22926_, _03897_);
  and (_22930_, _13402_, _05475_);
  or (_22931_, _22887_, _04790_);
  nor (_22932_, _22931_, _22930_);
  or (_22933_, _22932_, _04018_);
  nor (_22934_, _22933_, _22929_);
  and (_22935_, _08736_, _05475_);
  nor (_22936_, _22935_, _22887_);
  nor (_22937_, _22936_, _04792_);
  nor (_22938_, _22937_, _22934_);
  nor (_22940_, _22938_, _03908_);
  nor (_22941_, _22887_, _08322_);
  not (_22942_, _22941_);
  nor (_22943_, _22924_, _03909_);
  and (_22944_, _22943_, _22942_);
  nor (_22945_, _22944_, _22940_);
  nor (_22946_, _22945_, _04027_);
  nor (_22947_, _22889_, _04785_);
  and (_22948_, _22947_, _22942_);
  or (_22949_, _22948_, _22946_);
  and (_22950_, _22949_, _06567_);
  nor (_22951_, _13401_, _09595_);
  nor (_22952_, _22951_, _22887_);
  nor (_22953_, _22952_, _06567_);
  or (_22954_, _22953_, _22950_);
  and (_22955_, _22954_, _06572_);
  nor (_22956_, _08735_, _09595_);
  nor (_22957_, _22956_, _22887_);
  nor (_22958_, _22957_, _06572_);
  or (_22959_, _22958_, _03773_);
  nor (_22962_, _22959_, _22955_);
  and (_22963_, _22897_, _03773_);
  or (_22964_, _22963_, _03772_);
  nor (_22965_, _22964_, _22962_);
  nor (_22966_, _13460_, _09595_);
  nor (_22967_, _22966_, _22887_);
  nor (_22968_, _22967_, _04060_);
  or (_22969_, _22968_, _22965_);
  or (_22970_, _22969_, _43156_);
  or (_22971_, _43152_, \oc8051_golden_model_1.TMOD [6]);
  and (_22973_, _22971_, _41894_);
  and (_43470_, _22973_, _22970_);
  not (_22974_, \oc8051_golden_model_1.IE [0]);
  nor (_22975_, _05494_, _22974_);
  and (_22976_, _05716_, _05494_);
  nor (_22977_, _22976_, _22975_);
  nor (_22978_, _22977_, _04060_);
  nand (_22979_, _08753_, _05494_);
  nor (_22980_, _22975_, _04785_);
  and (_22981_, _22980_, _22979_);
  and (_22982_, _05494_, \oc8051_golden_model_1.ACC [0]);
  nor (_22983_, _22982_, _22975_);
  nor (_22984_, _22983_, _04708_);
  nor (_22985_, _04707_, _22974_);
  or (_22986_, _22985_, _22984_);
  and (_22987_, _22986_, _04722_);
  nor (_22988_, _22977_, _04722_);
  or (_22989_, _22988_, _22987_);
  and (_22990_, _22989_, _03764_);
  nor (_22991_, _06103_, _22974_);
  and (_22994_, _12064_, _06103_);
  nor (_22995_, _22994_, _22991_);
  nor (_22996_, _22995_, _03764_);
  nor (_22997_, _22996_, _22990_);
  nor (_22998_, _22997_, _03848_);
  and (_22999_, _05494_, _04700_);
  nor (_23000_, _22999_, _22975_);
  nor (_23001_, _23000_, _04733_);
  or (_23002_, _23001_, _22998_);
  and (_23003_, _23002_, _03855_);
  nor (_23005_, _22983_, _03855_);
  or (_23006_, _23005_, _23003_);
  and (_23007_, _23006_, _03760_);
  and (_23008_, _22975_, _03759_);
  or (_23009_, _23008_, _23007_);
  and (_23010_, _23009_, _03753_);
  nor (_23011_, _22977_, _03753_);
  or (_23012_, _23011_, _23010_);
  and (_23013_, _23012_, _03747_);
  nor (_23014_, _22991_, _14237_);
  or (_23015_, _23014_, _03747_);
  nor (_23016_, _23015_, _22995_);
  or (_23017_, _23016_, _07927_);
  or (_23018_, _23017_, _23013_);
  and (_23019_, _06962_, _05494_);
  nor (_23020_, _22975_, _03738_);
  not (_23021_, _23020_);
  nor (_23022_, _23021_, _23019_);
  and (_23023_, _23000_, _08474_);
  or (_23024_, _23023_, _03455_);
  nor (_23027_, _23024_, _23022_);
  and (_23028_, _23027_, _23018_);
  nor (_23029_, _12164_, _09694_);
  nor (_23030_, _23029_, _22975_);
  nor (_23031_, _23030_, _03820_);
  or (_23032_, _23031_, _23028_);
  and (_23033_, _23032_, _04778_);
  and (_23034_, _05494_, _06479_);
  nor (_23035_, _23034_, _22975_);
  nor (_23036_, _23035_, _04778_);
  or (_23038_, _23036_, _23033_);
  and (_23039_, _23038_, _04790_);
  and (_23040_, _12178_, _05494_);
  nor (_23041_, _23040_, _22975_);
  nor (_23042_, _23041_, _04790_);
  or (_23043_, _23042_, _23039_);
  and (_23044_, _23043_, _04792_);
  nor (_23045_, _10488_, _09694_);
  nor (_23046_, _23045_, _22975_);
  nand (_23047_, _22979_, _04018_);
  nor (_23048_, _23047_, _23046_);
  nor (_23049_, _23048_, _23044_);
  nor (_23050_, _23049_, _03908_);
  nor (_23051_, _23035_, _03909_);
  not (_23052_, _23051_);
  nor (_23053_, _23052_, _22976_);
  nor (_23054_, _23053_, _04027_);
  not (_23055_, _23054_);
  nor (_23056_, _23055_, _23050_);
  nor (_23057_, _23056_, _22981_);
  and (_23060_, _23057_, _06567_);
  nor (_23061_, _12177_, _09694_);
  nor (_23062_, _23061_, _22975_);
  nor (_23063_, _23062_, _06567_);
  or (_23064_, _23063_, _23060_);
  and (_23065_, _23064_, _06572_);
  nor (_23066_, _23046_, _06572_);
  or (_23067_, _23066_, _03773_);
  or (_23068_, _23067_, _23065_);
  nand (_23069_, _22977_, _03773_);
  and (_23071_, _23069_, _23068_);
  nor (_23072_, _23071_, _03374_);
  nor (_23073_, _22975_, _03375_);
  nor (_23074_, _23073_, _23072_);
  and (_23075_, _23074_, _04060_);
  nor (_23076_, _23075_, _22978_);
  nand (_23077_, _23076_, _43152_);
  or (_23078_, _43152_, \oc8051_golden_model_1.IE [0]);
  and (_23079_, _23078_, _41894_);
  and (_43473_, _23079_, _23077_);
  and (_23080_, _05494_, _04595_);
  not (_23081_, _23080_);
  nor (_23082_, _05494_, \oc8051_golden_model_1.IE [1]);
  nor (_23083_, _23082_, _04778_);
  and (_23084_, _23083_, _23081_);
  not (_23085_, \oc8051_golden_model_1.IE [1]);
  nor (_23086_, _05494_, _23085_);
  and (_23087_, _05494_, \oc8051_golden_model_1.ACC [1]);
  nor (_23088_, _23087_, _23086_);
  nor (_23089_, _23088_, _04708_);
  nor (_23092_, _04707_, _23085_);
  or (_23093_, _23092_, _23089_);
  and (_23094_, _23093_, _04722_);
  and (_23095_, _12262_, _05494_);
  nor (_23096_, _23095_, _23082_);
  and (_23097_, _23096_, _03850_);
  or (_23098_, _23097_, _23094_);
  and (_23099_, _23098_, _03764_);
  nor (_23100_, _06103_, _23085_);
  and (_23101_, _12249_, _06103_);
  nor (_23103_, _23101_, _23100_);
  nor (_23104_, _23103_, _03764_);
  or (_23105_, _23104_, _23099_);
  and (_23106_, _23105_, _04733_);
  and (_23107_, _05494_, _04900_);
  nor (_23108_, _23107_, _23086_);
  nor (_23109_, _23108_, _04733_);
  or (_23110_, _23109_, _23106_);
  and (_23111_, _23110_, _03855_);
  nor (_23112_, _23088_, _03855_);
  or (_23114_, _23112_, _23111_);
  and (_23115_, _23114_, _03760_);
  and (_23116_, _12252_, _06103_);
  nor (_23117_, _23116_, _23100_);
  nor (_23118_, _23117_, _03760_);
  or (_23119_, _23118_, _03752_);
  or (_23120_, _23119_, _23115_);
  and (_23121_, _23101_, _12248_);
  or (_23122_, _23100_, _03753_);
  or (_23123_, _23122_, _23121_);
  and (_23125_, _23123_, _03747_);
  and (_23126_, _23125_, _23120_);
  nor (_23127_, _12293_, _09680_);
  nor (_23128_, _23127_, _23100_);
  nor (_23129_, _23128_, _03747_);
  or (_23130_, _23129_, _07927_);
  or (_23131_, _23130_, _23126_);
  and (_23132_, _06961_, _05494_);
  nor (_23133_, _23086_, _03738_);
  not (_23134_, _23133_);
  nor (_23136_, _23134_, _23132_);
  and (_23137_, _23108_, _08474_);
  or (_23138_, _23137_, _03455_);
  nor (_23139_, _23138_, _23136_);
  and (_23140_, _23139_, _23131_);
  nor (_23141_, _12352_, _09694_);
  nor (_23142_, _23141_, _23086_);
  nor (_23143_, _23142_, _03820_);
  nor (_23144_, _23143_, _23140_);
  nor (_23145_, _23144_, _03903_);
  nor (_23147_, _23145_, _23084_);
  nor (_23148_, _23147_, _03897_);
  and (_23149_, _12366_, _05494_);
  or (_23150_, _23149_, _23086_);
  and (_23151_, _23150_, _03897_);
  nor (_23152_, _23151_, _23148_);
  nor (_23153_, _23152_, _04018_);
  nor (_23154_, _08751_, _09694_);
  nor (_23155_, _23154_, _23086_);
  and (_23156_, _08750_, _05494_);
  nor (_23158_, _23156_, _23155_);
  and (_23159_, _23158_, _04018_);
  or (_23160_, _23159_, _23153_);
  and (_23161_, _23160_, _03909_);
  and (_23162_, _12244_, _05494_);
  or (_23163_, _23162_, _23086_);
  and (_23164_, _23163_, _03908_);
  or (_23165_, _23164_, _23161_);
  and (_23166_, _23165_, _04785_);
  nor (_23167_, _23156_, _23086_);
  nor (_23169_, _23167_, _04785_);
  or (_23170_, _23169_, _23166_);
  and (_23171_, _23170_, _06567_);
  nor (_23172_, _12365_, _09694_);
  or (_23173_, _23172_, _23086_);
  and (_23174_, _23173_, _03914_);
  or (_23175_, _23174_, _23171_);
  and (_23176_, _23175_, _06572_);
  nor (_23177_, _23155_, _06572_);
  or (_23178_, _23177_, _23176_);
  and (_23180_, _23178_, _03774_);
  and (_23181_, _23096_, _03773_);
  or (_23182_, _23181_, _23180_);
  and (_23183_, _23182_, _03375_);
  nor (_23184_, _23117_, _03375_);
  nor (_23185_, _23184_, _03772_);
  not (_23186_, _23185_);
  nor (_23187_, _23186_, _23183_);
  nor (_23188_, _23095_, _23086_);
  and (_23189_, _23188_, _03772_);
  nor (_23191_, _23189_, _23187_);
  or (_23192_, _23191_, _43156_);
  or (_23193_, _43152_, \oc8051_golden_model_1.IE [1]);
  and (_23194_, _23193_, _41894_);
  and (_43474_, _23194_, _23192_);
  not (_23195_, \oc8051_golden_model_1.IE [2]);
  nor (_23196_, _05494_, _23195_);
  and (_23197_, _05494_, \oc8051_golden_model_1.ACC [2]);
  nor (_23198_, _23197_, _23196_);
  nor (_23199_, _23198_, _04708_);
  nor (_23201_, _04707_, _23195_);
  or (_23202_, _23201_, _23199_);
  and (_23203_, _23202_, _04722_);
  nor (_23204_, _12471_, _09694_);
  nor (_23205_, _23204_, _23196_);
  nor (_23206_, _23205_, _04722_);
  or (_23207_, _23206_, _23203_);
  and (_23208_, _23207_, _03764_);
  nor (_23209_, _06103_, _23195_);
  and (_23210_, _12464_, _06103_);
  nor (_23212_, _23210_, _23209_);
  nor (_23213_, _23212_, _03764_);
  or (_23214_, _23213_, _23208_);
  and (_23215_, _23214_, _04733_);
  and (_23216_, _05494_, _05307_);
  nor (_23217_, _23216_, _23196_);
  nor (_23218_, _23217_, _04733_);
  or (_23219_, _23218_, _23215_);
  and (_23220_, _23219_, _03855_);
  nor (_23221_, _23198_, _03855_);
  or (_23223_, _23221_, _23220_);
  and (_23224_, _23223_, _03760_);
  and (_23225_, _12467_, _06103_);
  nor (_23226_, _23225_, _23209_);
  nor (_23227_, _23226_, _03760_);
  or (_23228_, _23227_, _03752_);
  or (_23229_, _23228_, _23224_);
  and (_23230_, _23210_, _12463_);
  or (_23231_, _23209_, _03753_);
  or (_23232_, _23231_, _23230_);
  and (_23234_, _23232_, _03747_);
  and (_23235_, _23234_, _23229_);
  nor (_23236_, _12514_, _09680_);
  nor (_23237_, _23236_, _23209_);
  nor (_23238_, _23237_, _03747_);
  or (_23239_, _23238_, _07927_);
  or (_23240_, _23239_, _23235_);
  and (_23241_, _06965_, _05494_);
  nor (_23242_, _23196_, _03738_);
  not (_23243_, _23242_);
  nor (_23245_, _23243_, _23241_);
  and (_23246_, _23217_, _08474_);
  or (_23247_, _23246_, _03455_);
  nor (_23248_, _23247_, _23245_);
  and (_23249_, _23248_, _23240_);
  nor (_23250_, _12572_, _09694_);
  nor (_23251_, _23250_, _23196_);
  nor (_23252_, _23251_, _03820_);
  or (_23253_, _23252_, _23249_);
  and (_23254_, _23253_, _04778_);
  and (_23256_, _05494_, _06495_);
  nor (_23257_, _23256_, _23196_);
  nor (_23258_, _23257_, _04778_);
  or (_23259_, _23258_, _23254_);
  and (_23260_, _23259_, _04790_);
  and (_23261_, _12586_, _05494_);
  nor (_23262_, _23261_, _23196_);
  nor (_23263_, _23262_, _04790_);
  or (_23264_, _23263_, _23260_);
  and (_23265_, _23264_, _04792_);
  and (_23267_, _08748_, _05494_);
  nor (_23268_, _23267_, _23196_);
  nor (_23269_, _23268_, _04792_);
  nor (_23270_, _23269_, _23265_);
  nor (_23271_, _23270_, _03908_);
  nor (_23272_, _23196_, _05765_);
  not (_23273_, _23272_);
  nor (_23274_, _23257_, _03909_);
  and (_23275_, _23274_, _23273_);
  nor (_23276_, _23275_, _23271_);
  nor (_23278_, _23276_, _04027_);
  nor (_23279_, _23198_, _04785_);
  and (_23280_, _23279_, _23273_);
  or (_23281_, _23280_, _23278_);
  and (_23282_, _23281_, _06567_);
  nor (_23283_, _12585_, _09694_);
  nor (_23284_, _23283_, _23196_);
  nor (_23285_, _23284_, _06567_);
  or (_23286_, _23285_, _23282_);
  and (_23287_, _23286_, _06572_);
  nor (_23289_, _08747_, _09694_);
  nor (_23290_, _23289_, _23196_);
  nor (_23291_, _23290_, _06572_);
  or (_23292_, _23291_, _23287_);
  and (_23293_, _23292_, _03774_);
  nor (_23294_, _23205_, _03774_);
  or (_23295_, _23294_, _23293_);
  and (_23296_, _23295_, _03375_);
  nor (_23297_, _23226_, _03375_);
  or (_23298_, _23297_, _23296_);
  and (_23300_, _23298_, _04060_);
  and (_23301_, _12642_, _05494_);
  nor (_23302_, _23301_, _23196_);
  nor (_23303_, _23302_, _04060_);
  or (_23304_, _23303_, _23300_);
  or (_23305_, _23304_, _43156_);
  or (_23306_, _43152_, \oc8051_golden_model_1.IE [2]);
  and (_23307_, _23306_, _41894_);
  and (_43475_, _23307_, _23305_);
  not (_23308_, \oc8051_golden_model_1.IE [3]);
  nor (_23310_, _05494_, _23308_);
  and (_23311_, _05494_, \oc8051_golden_model_1.ACC [3]);
  nor (_23312_, _23311_, _23310_);
  nor (_23313_, _23312_, _04708_);
  nor (_23314_, _04707_, _23308_);
  or (_23315_, _23314_, _23313_);
  and (_23316_, _23315_, _04722_);
  nor (_23317_, _12681_, _09694_);
  nor (_23318_, _23317_, _23310_);
  nor (_23319_, _23318_, _04722_);
  or (_23321_, _23319_, _23316_);
  and (_23322_, _23321_, _03764_);
  nor (_23323_, _06103_, _23308_);
  and (_23324_, _12674_, _06103_);
  nor (_23325_, _23324_, _23323_);
  nor (_23326_, _23325_, _03764_);
  or (_23327_, _23326_, _03848_);
  or (_23328_, _23327_, _23322_);
  and (_23329_, _05494_, _05119_);
  nor (_23330_, _23329_, _23310_);
  nand (_23332_, _23330_, _03848_);
  and (_23333_, _23332_, _23328_);
  and (_23334_, _23333_, _03855_);
  nor (_23335_, _23312_, _03855_);
  or (_23336_, _23335_, _23334_);
  and (_23337_, _23336_, _03760_);
  and (_23338_, _12667_, _06103_);
  nor (_23339_, _23338_, _23323_);
  nor (_23340_, _23339_, _03760_);
  or (_23341_, _23340_, _03752_);
  or (_23343_, _23341_, _23337_);
  nor (_23344_, _23323_, _12673_);
  nor (_23345_, _23344_, _23325_);
  or (_23346_, _23345_, _03753_);
  and (_23347_, _23346_, _03747_);
  and (_23348_, _23347_, _23343_);
  nor (_23349_, _12668_, _09680_);
  nor (_23350_, _23349_, _23323_);
  nor (_23351_, _23350_, _03747_);
  or (_23352_, _23351_, _07927_);
  or (_23354_, _23352_, _23348_);
  and (_23355_, _06964_, _05494_);
  nor (_23356_, _23310_, _03738_);
  not (_23357_, _23356_);
  nor (_23358_, _23357_, _23355_);
  and (_23359_, _23330_, _08474_);
  or (_23360_, _23359_, _03455_);
  nor (_23361_, _23360_, _23358_);
  and (_23362_, _23361_, _23354_);
  nor (_23363_, _12775_, _09694_);
  nor (_23365_, _23363_, _23310_);
  nor (_23366_, _23365_, _03820_);
  or (_23367_, _23366_, _23362_);
  and (_23368_, _23367_, _04778_);
  and (_23369_, _05494_, _06345_);
  nor (_23370_, _23369_, _23310_);
  nor (_23371_, _23370_, _04778_);
  or (_23372_, _23371_, _23368_);
  and (_23373_, _23372_, _04790_);
  and (_23374_, _12789_, _05494_);
  nor (_23376_, _23374_, _23310_);
  nor (_23377_, _23376_, _04790_);
  or (_23378_, _23377_, _23373_);
  and (_23379_, _23378_, _04792_);
  and (_23380_, _10491_, _05494_);
  nor (_23381_, _23380_, _23310_);
  nor (_23382_, _23381_, _04792_);
  nor (_23383_, _23382_, _23379_);
  nor (_23384_, _23383_, _03908_);
  nor (_23385_, _23310_, _05622_);
  not (_23387_, _23385_);
  nor (_23388_, _23370_, _03909_);
  and (_23389_, _23388_, _23387_);
  nor (_23390_, _23389_, _23384_);
  nor (_23391_, _23390_, _04027_);
  nor (_23392_, _23312_, _04785_);
  and (_23393_, _23392_, _23387_);
  or (_23394_, _23393_, _23391_);
  and (_23395_, _23394_, _06567_);
  nor (_23396_, _12788_, _09694_);
  nor (_23398_, _23396_, _23310_);
  nor (_23399_, _23398_, _06567_);
  or (_23400_, _23399_, _23395_);
  and (_23401_, _23400_, _06572_);
  nor (_23402_, _08742_, _09694_);
  nor (_23403_, _23402_, _23310_);
  nor (_23404_, _23403_, _06572_);
  or (_23405_, _23404_, _23401_);
  and (_23406_, _23405_, _03774_);
  nor (_23407_, _23318_, _03774_);
  or (_23409_, _23407_, _23406_);
  and (_23410_, _23409_, _03375_);
  nor (_23411_, _23339_, _03375_);
  or (_23412_, _23411_, _23410_);
  and (_23413_, _23412_, _04060_);
  and (_23414_, _12848_, _05494_);
  nor (_23415_, _23414_, _23310_);
  nor (_23416_, _23415_, _04060_);
  or (_23417_, _23416_, _23413_);
  or (_23418_, _23417_, _43156_);
  or (_23420_, _43152_, \oc8051_golden_model_1.IE [3]);
  and (_23421_, _23420_, _41894_);
  and (_43476_, _23421_, _23418_);
  not (_23422_, \oc8051_golden_model_1.IE [4]);
  nor (_23423_, _05494_, _23422_);
  and (_23424_, _05494_, \oc8051_golden_model_1.ACC [4]);
  nor (_23425_, _23424_, _23423_);
  nor (_23426_, _23425_, _04708_);
  nor (_23427_, _04707_, _23422_);
  or (_23428_, _23427_, _23426_);
  and (_23430_, _23428_, _04722_);
  nor (_23431_, _12891_, _09694_);
  nor (_23432_, _23431_, _23423_);
  nor (_23433_, _23432_, _04722_);
  or (_23434_, _23433_, _23430_);
  and (_23435_, _23434_, _03764_);
  nor (_23436_, _06103_, _23422_);
  and (_23437_, _12875_, _06103_);
  nor (_23438_, _23437_, _23436_);
  nor (_23439_, _23438_, _03764_);
  or (_23441_, _23439_, _03848_);
  or (_23442_, _23441_, _23435_);
  and (_23443_, _05950_, _05494_);
  nor (_23444_, _23443_, _23423_);
  nand (_23445_, _23444_, _03848_);
  and (_23446_, _23445_, _23442_);
  and (_23447_, _23446_, _03855_);
  nor (_23448_, _23425_, _03855_);
  or (_23449_, _23448_, _23447_);
  and (_23450_, _23449_, _03760_);
  and (_23452_, _12870_, _06103_);
  nor (_23453_, _23452_, _23436_);
  nor (_23454_, _23453_, _03760_);
  or (_23455_, _23454_, _03752_);
  or (_23456_, _23455_, _23450_);
  nor (_23457_, _23436_, _12874_);
  nor (_23458_, _23457_, _23438_);
  or (_23459_, _23458_, _03753_);
  and (_23460_, _23459_, _03747_);
  and (_23461_, _23460_, _23456_);
  nor (_23463_, _12872_, _09680_);
  nor (_23464_, _23463_, _23436_);
  nor (_23465_, _23464_, _03747_);
  or (_23466_, _23465_, _07927_);
  or (_23467_, _23466_, _23461_);
  and (_23468_, _06969_, _05494_);
  nor (_23469_, _23423_, _03738_);
  not (_23470_, _23469_);
  nor (_23471_, _23470_, _23468_);
  and (_23472_, _23444_, _08474_);
  or (_23474_, _23472_, _03455_);
  nor (_23475_, _23474_, _23471_);
  and (_23476_, _23475_, _23467_);
  nor (_23477_, _12982_, _09694_);
  nor (_23478_, _23477_, _23423_);
  nor (_23479_, _23478_, _03820_);
  or (_23480_, _23479_, _23476_);
  and (_23481_, _23480_, _04778_);
  and (_23482_, _06456_, _05494_);
  nor (_23483_, _23482_, _23423_);
  nor (_23485_, _23483_, _04778_);
  or (_23486_, _23485_, _23481_);
  and (_23487_, _23486_, _04790_);
  and (_23488_, _12997_, _05494_);
  nor (_23489_, _23488_, _23423_);
  nor (_23490_, _23489_, _04790_);
  or (_23491_, _23490_, _23487_);
  and (_23492_, _23491_, _04792_);
  and (_23493_, _08741_, _05494_);
  nor (_23494_, _23493_, _23423_);
  nor (_23496_, _23494_, _04792_);
  nor (_23497_, _23496_, _23492_);
  nor (_23498_, _23497_, _03908_);
  nor (_23499_, _23423_, _08336_);
  not (_23500_, _23499_);
  nor (_23501_, _23483_, _03909_);
  and (_23502_, _23501_, _23500_);
  nor (_23503_, _23502_, _23498_);
  nor (_23504_, _23503_, _04027_);
  nor (_23505_, _23425_, _04785_);
  and (_23507_, _23505_, _23500_);
  or (_23508_, _23507_, _23504_);
  and (_23509_, _23508_, _06567_);
  nor (_23510_, _12996_, _09694_);
  nor (_23511_, _23510_, _23423_);
  nor (_23512_, _23511_, _06567_);
  or (_23513_, _23512_, _23509_);
  and (_23514_, _23513_, _06572_);
  nor (_23515_, _08740_, _09694_);
  nor (_23516_, _23515_, _23423_);
  nor (_23518_, _23516_, _06572_);
  or (_23519_, _23518_, _23514_);
  and (_23520_, _23519_, _03774_);
  nor (_23521_, _23432_, _03774_);
  or (_23522_, _23521_, _23520_);
  and (_23523_, _23522_, _03375_);
  nor (_23524_, _23453_, _03375_);
  or (_23525_, _23524_, _23523_);
  and (_23526_, _23525_, _04060_);
  and (_23527_, _13056_, _05494_);
  nor (_23529_, _23527_, _23423_);
  nor (_23530_, _23529_, _04060_);
  or (_23531_, _23530_, _23526_);
  or (_23532_, _23531_, _43156_);
  or (_23533_, _43152_, \oc8051_golden_model_1.IE [4]);
  and (_23534_, _23533_, _41894_);
  and (_43477_, _23534_, _23532_);
  not (_23535_, \oc8051_golden_model_1.IE [5]);
  nor (_23536_, _05494_, _23535_);
  and (_23537_, _05494_, \oc8051_golden_model_1.ACC [5]);
  nor (_23539_, _23537_, _23536_);
  nor (_23540_, _23539_, _04708_);
  nor (_23541_, _04707_, _23535_);
  or (_23542_, _23541_, _23540_);
  and (_23543_, _23542_, _04722_);
  nor (_23544_, _13090_, _09694_);
  nor (_23545_, _23544_, _23536_);
  nor (_23546_, _23545_, _04722_);
  or (_23547_, _23546_, _23543_);
  and (_23548_, _23547_, _03764_);
  nor (_23550_, _06103_, _23535_);
  and (_23551_, _13094_, _06103_);
  nor (_23552_, _23551_, _23550_);
  nor (_23553_, _23552_, _03764_);
  or (_23554_, _23553_, _03848_);
  or (_23555_, _23554_, _23548_);
  and (_23556_, _05857_, _05494_);
  nor (_23557_, _23556_, _23536_);
  nand (_23558_, _23557_, _03848_);
  and (_23559_, _23558_, _23555_);
  and (_23561_, _23559_, _03855_);
  nor (_23562_, _23539_, _03855_);
  or (_23563_, _23562_, _23561_);
  and (_23564_, _23563_, _03760_);
  and (_23565_, _13071_, _06103_);
  nor (_23566_, _23565_, _23550_);
  nor (_23567_, _23566_, _03760_);
  or (_23568_, _23567_, _03752_);
  or (_23569_, _23568_, _23564_);
  nor (_23570_, _23550_, _13109_);
  nor (_23572_, _23570_, _23552_);
  or (_23573_, _23572_, _03753_);
  and (_23574_, _23573_, _03747_);
  and (_23575_, _23574_, _23569_);
  nor (_23576_, _13073_, _09680_);
  nor (_23577_, _23576_, _23550_);
  nor (_23578_, _23577_, _03747_);
  or (_23579_, _23578_, _07927_);
  or (_23580_, _23579_, _23575_);
  and (_23581_, _06968_, _05494_);
  nor (_23583_, _23536_, _03738_);
  not (_23584_, _23583_);
  nor (_23585_, _23584_, _23581_);
  and (_23586_, _23557_, _08474_);
  or (_23587_, _23586_, _03455_);
  nor (_23588_, _23587_, _23585_);
  and (_23589_, _23588_, _23580_);
  nor (_23590_, _13182_, _09694_);
  nor (_23591_, _23590_, _23536_);
  nor (_23592_, _23591_, _03820_);
  or (_23594_, _23592_, _23589_);
  and (_23595_, _23594_, _04778_);
  and (_23596_, _06447_, _05494_);
  nor (_23597_, _23596_, _23536_);
  nor (_23598_, _23597_, _04778_);
  or (_23599_, _23598_, _23595_);
  and (_23600_, _23599_, _04790_);
  and (_23601_, _13196_, _05494_);
  nor (_23602_, _23601_, _23536_);
  nor (_23603_, _23602_, _04790_);
  or (_23605_, _23603_, _23600_);
  and (_23606_, _23605_, _04792_);
  and (_23607_, _10493_, _05494_);
  nor (_23608_, _23607_, _23536_);
  nor (_23609_, _23608_, _04792_);
  nor (_23610_, _23609_, _23606_);
  nor (_23611_, _23610_, _03908_);
  nor (_23612_, _23536_, _08335_);
  not (_23613_, _23612_);
  nor (_23614_, _23597_, _03909_);
  and (_23616_, _23614_, _23613_);
  nor (_23617_, _23616_, _23611_);
  nor (_23618_, _23617_, _04027_);
  nor (_23619_, _23539_, _04785_);
  and (_23620_, _23619_, _23613_);
  or (_23621_, _23620_, _23618_);
  and (_23622_, _23621_, _06567_);
  nor (_23623_, _13195_, _09694_);
  nor (_23624_, _23623_, _23536_);
  nor (_23625_, _23624_, _06567_);
  or (_23627_, _23625_, _23622_);
  and (_23628_, _23627_, _06572_);
  nor (_23629_, _08738_, _09694_);
  nor (_23630_, _23629_, _23536_);
  nor (_23631_, _23630_, _06572_);
  or (_23632_, _23631_, _23628_);
  and (_23633_, _23632_, _03774_);
  nor (_23634_, _23545_, _03774_);
  or (_23635_, _23634_, _23633_);
  and (_23636_, _23635_, _03375_);
  nor (_23638_, _23566_, _03375_);
  or (_23639_, _23638_, _23636_);
  and (_23640_, _23639_, _04060_);
  and (_23641_, _13255_, _05494_);
  nor (_23642_, _23641_, _23536_);
  nor (_23643_, _23642_, _04060_);
  or (_23644_, _23643_, _23640_);
  or (_23645_, _23644_, _43156_);
  or (_23646_, _43152_, \oc8051_golden_model_1.IE [5]);
  and (_23647_, _23646_, _41894_);
  and (_43478_, _23647_, _23645_);
  not (_23649_, \oc8051_golden_model_1.IE [6]);
  nor (_23650_, _05494_, _23649_);
  and (_23651_, _05494_, \oc8051_golden_model_1.ACC [6]);
  nor (_23652_, _23651_, _23650_);
  nor (_23653_, _23652_, _04708_);
  nor (_23654_, _04707_, _23649_);
  or (_23655_, _23654_, _23653_);
  and (_23656_, _23655_, _04722_);
  nor (_23657_, _13293_, _09694_);
  nor (_23659_, _23657_, _23650_);
  nor (_23660_, _23659_, _04722_);
  or (_23661_, _23660_, _23656_);
  and (_23662_, _23661_, _03764_);
  nor (_23663_, _06103_, _23649_);
  and (_23664_, _13297_, _06103_);
  nor (_23665_, _23664_, _23663_);
  nor (_23666_, _23665_, _03764_);
  or (_23667_, _23666_, _03848_);
  or (_23668_, _23667_, _23662_);
  and (_23670_, _06065_, _05494_);
  nor (_23671_, _23670_, _23650_);
  nand (_23672_, _23671_, _03848_);
  and (_23673_, _23672_, _23668_);
  and (_23674_, _23673_, _03855_);
  nor (_23675_, _23652_, _03855_);
  or (_23676_, _23675_, _23674_);
  and (_23677_, _23676_, _03760_);
  and (_23678_, _13277_, _06103_);
  nor (_23679_, _23678_, _23663_);
  nor (_23681_, _23679_, _03760_);
  or (_23682_, _23681_, _23677_);
  and (_23683_, _23682_, _03753_);
  nor (_23684_, _23663_, _13312_);
  nor (_23685_, _23684_, _23665_);
  and (_23686_, _23685_, _03752_);
  or (_23687_, _23686_, _23683_);
  and (_23688_, _23687_, _03747_);
  nor (_23689_, _13279_, _09680_);
  nor (_23690_, _23689_, _23663_);
  nor (_23692_, _23690_, _03747_);
  or (_23693_, _23692_, _07927_);
  or (_23694_, _23693_, _23688_);
  and (_23695_, _06641_, _05494_);
  nor (_23696_, _23650_, _03738_);
  not (_23697_, _23696_);
  nor (_23698_, _23697_, _23695_);
  and (_23699_, _23671_, _08474_);
  or (_23700_, _23699_, _03455_);
  nor (_23701_, _23700_, _23698_);
  and (_23703_, _23701_, _23694_);
  nor (_23704_, _13387_, _09694_);
  nor (_23705_, _23704_, _23650_);
  nor (_23706_, _23705_, _03820_);
  or (_23707_, _23706_, _23703_);
  and (_23708_, _23707_, _04778_);
  and (_23709_, _13394_, _05494_);
  nor (_23710_, _23709_, _23650_);
  nor (_23711_, _23710_, _04778_);
  or (_23712_, _23711_, _23708_);
  nor (_23714_, _23712_, _03897_);
  and (_23715_, _13402_, _05494_);
  or (_23716_, _23650_, _04790_);
  nor (_23717_, _23716_, _23715_);
  or (_23718_, _23717_, _04018_);
  nor (_23719_, _23718_, _23714_);
  and (_23720_, _08736_, _05494_);
  nor (_23721_, _23720_, _23650_);
  nor (_23722_, _23721_, _04792_);
  nor (_23723_, _23722_, _23719_);
  nor (_23725_, _23723_, _03908_);
  nor (_23726_, _23650_, _08322_);
  not (_23727_, _23726_);
  nor (_23728_, _23710_, _03909_);
  and (_23729_, _23728_, _23727_);
  nor (_23730_, _23729_, _23725_);
  nor (_23731_, _23730_, _04027_);
  nor (_23732_, _23652_, _04785_);
  and (_23733_, _23732_, _23727_);
  or (_23734_, _23733_, _23731_);
  and (_23736_, _23734_, _06567_);
  nor (_23737_, _13401_, _09694_);
  nor (_23738_, _23737_, _23650_);
  nor (_23739_, _23738_, _06567_);
  or (_23740_, _23739_, _23736_);
  and (_23741_, _23740_, _06572_);
  nor (_23742_, _08735_, _09694_);
  nor (_23743_, _23742_, _23650_);
  nor (_23744_, _23743_, _06572_);
  or (_23745_, _23744_, _23741_);
  and (_23747_, _23745_, _03774_);
  nor (_23748_, _23659_, _03774_);
  or (_23749_, _23748_, _23747_);
  and (_23750_, _23749_, _03375_);
  nor (_23751_, _23679_, _03375_);
  or (_23752_, _23751_, _23750_);
  and (_23753_, _23752_, _04060_);
  nor (_23754_, _13460_, _09694_);
  nor (_23755_, _23754_, _23650_);
  nor (_23756_, _23755_, _04060_);
  or (_23758_, _23756_, _23753_);
  or (_23759_, _23758_, _43156_);
  or (_23760_, _43152_, \oc8051_golden_model_1.IE [6]);
  and (_23761_, _23760_, _41894_);
  and (_43479_, _23761_, _23759_);
  not (_23762_, \oc8051_golden_model_1.IP [0]);
  nor (_23763_, _05437_, _23762_);
  and (_23764_, _05716_, _05437_);
  nor (_23765_, _23764_, _23763_);
  nor (_23766_, _23765_, _04060_);
  nand (_23768_, _08753_, _05437_);
  nor (_23769_, _23763_, _04785_);
  and (_23770_, _23769_, _23768_);
  and (_23771_, _06962_, _05437_);
  nor (_23772_, _23763_, _03738_);
  not (_23773_, _23772_);
  nor (_23774_, _23773_, _23771_);
  nor (_23775_, _23765_, _04722_);
  nor (_23776_, _04707_, _23762_);
  and (_23777_, _05437_, \oc8051_golden_model_1.ACC [0]);
  nor (_23778_, _23777_, _23763_);
  nor (_23779_, _23778_, _04708_);
  nor (_23780_, _23779_, _23776_);
  nor (_23781_, _23780_, _03850_);
  or (_23782_, _23781_, _03763_);
  nor (_23783_, _23782_, _23775_);
  and (_23784_, _12064_, _06091_);
  nor (_23785_, _06091_, _23762_);
  or (_23786_, _23785_, _03764_);
  nor (_23787_, _23786_, _23784_);
  nor (_23789_, _23787_, _23783_);
  and (_23790_, _23789_, _04733_);
  and (_23791_, _05437_, _04700_);
  nor (_23792_, _23791_, _23763_);
  nor (_23793_, _23792_, _04733_);
  or (_23794_, _23793_, _23790_);
  and (_23795_, _23794_, _03855_);
  nor (_23796_, _23778_, _03855_);
  or (_23797_, _23796_, _23795_);
  and (_23798_, _23797_, _03760_);
  and (_23800_, _23763_, _03759_);
  or (_23801_, _23800_, _23798_);
  and (_23802_, _23801_, _03753_);
  nor (_23803_, _23765_, _03753_);
  or (_23804_, _23803_, _23802_);
  and (_23805_, _23804_, _03747_);
  and (_23806_, _23784_, _14237_);
  nor (_23807_, _23806_, _23785_);
  nor (_23808_, _23807_, _03747_);
  or (_23809_, _23808_, _07927_);
  nor (_23810_, _23809_, _23805_);
  and (_23811_, _23792_, _08474_);
  or (_23812_, _23811_, _03455_);
  or (_23813_, _23812_, _23810_);
  nor (_23814_, _23813_, _23774_);
  nor (_23815_, _12164_, _09799_);
  nor (_23816_, _23815_, _23763_);
  nor (_23817_, _23816_, _03820_);
  or (_23818_, _23817_, _23814_);
  and (_23819_, _23818_, _04778_);
  and (_23820_, _05437_, _06479_);
  nor (_23821_, _23820_, _23763_);
  nor (_23822_, _23821_, _04778_);
  or (_23823_, _23822_, _23819_);
  and (_23824_, _23823_, _04790_);
  and (_23825_, _12178_, _05437_);
  nor (_23826_, _23825_, _23763_);
  nor (_23827_, _23826_, _04790_);
  or (_23828_, _23827_, _23824_);
  and (_23829_, _23828_, _04792_);
  nor (_23830_, _10488_, _09799_);
  nor (_23831_, _23830_, _23763_);
  nand (_23832_, _23768_, _04018_);
  nor (_23833_, _23832_, _23831_);
  nor (_23834_, _23833_, _23829_);
  nor (_23835_, _23834_, _03908_);
  nor (_23836_, _23821_, _03909_);
  not (_23837_, _23836_);
  nor (_23838_, _23837_, _23764_);
  nor (_23839_, _23838_, _04027_);
  not (_23840_, _23839_);
  nor (_23841_, _23840_, _23835_);
  nor (_23842_, _23841_, _23770_);
  and (_23843_, _23842_, _06567_);
  nor (_23844_, _12177_, _09799_);
  nor (_23845_, _23844_, _23763_);
  nor (_23846_, _23845_, _06567_);
  or (_23847_, _23846_, _23843_);
  and (_23848_, _23847_, _06572_);
  nor (_23849_, _23831_, _06572_);
  or (_23850_, _23849_, _03773_);
  or (_23851_, _23850_, _23848_);
  nand (_23852_, _23765_, _03773_);
  and (_23853_, _23852_, _23851_);
  nor (_23854_, _23853_, _03374_);
  nor (_23855_, _23763_, _03375_);
  nor (_23856_, _23855_, _23854_);
  and (_23857_, _23856_, _04060_);
  nor (_23858_, _23857_, _23766_);
  nand (_23859_, _23858_, _43152_);
  or (_23861_, _43152_, \oc8051_golden_model_1.IP [0]);
  and (_23862_, _23861_, _41894_);
  and (_43480_, _23862_, _23859_);
  not (_23863_, \oc8051_golden_model_1.IP [1]);
  nor (_23864_, _05437_, _23863_);
  and (_23865_, _05437_, \oc8051_golden_model_1.ACC [1]);
  nor (_23866_, _23865_, _23864_);
  nor (_23867_, _23866_, _04708_);
  nor (_23868_, _04707_, _23863_);
  or (_23869_, _23868_, _23867_);
  and (_23871_, _23869_, _04722_);
  nor (_23872_, _05437_, \oc8051_golden_model_1.IP [1]);
  and (_23873_, _12262_, _05437_);
  nor (_23874_, _23873_, _23872_);
  and (_23875_, _23874_, _03850_);
  or (_23876_, _23875_, _23871_);
  and (_23877_, _23876_, _03764_);
  nor (_23878_, _06091_, _23863_);
  and (_23879_, _12249_, _06091_);
  nor (_23880_, _23879_, _23878_);
  nor (_23881_, _23880_, _03764_);
  or (_23882_, _23881_, _23877_);
  and (_23883_, _23882_, _04733_);
  and (_23884_, _05437_, _04900_);
  nor (_23885_, _23884_, _23864_);
  nor (_23886_, _23885_, _04733_);
  or (_23887_, _23886_, _23883_);
  and (_23888_, _23887_, _03855_);
  nor (_23889_, _23866_, _03855_);
  or (_23890_, _23889_, _23888_);
  and (_23892_, _23890_, _03760_);
  and (_23893_, _12252_, _06091_);
  nor (_23894_, _23893_, _23878_);
  nor (_23895_, _23894_, _03760_);
  or (_23896_, _23895_, _03752_);
  or (_23897_, _23896_, _23892_);
  and (_23898_, _23879_, _12248_);
  or (_23899_, _23878_, _03753_);
  or (_23900_, _23899_, _23898_);
  and (_23901_, _23900_, _03747_);
  and (_23903_, _23901_, _23897_);
  nor (_23904_, _12293_, _09785_);
  nor (_23905_, _23904_, _23878_);
  nor (_23906_, _23905_, _03747_);
  or (_23907_, _23906_, _07927_);
  or (_23908_, _23907_, _23903_);
  and (_23909_, _06961_, _05437_);
  nor (_23910_, _23864_, _03738_);
  not (_23911_, _23910_);
  nor (_23912_, _23911_, _23909_);
  and (_23914_, _23885_, _08474_);
  or (_23915_, _23914_, _03455_);
  nor (_23916_, _23915_, _23912_);
  and (_23917_, _23916_, _23908_);
  nor (_23918_, _12352_, _09799_);
  nor (_23919_, _23918_, _23864_);
  nor (_23920_, _23919_, _03820_);
  nor (_23921_, _23920_, _23917_);
  nor (_23922_, _23921_, _03903_);
  and (_23923_, _05437_, _04595_);
  not (_23925_, _23923_);
  nor (_23926_, _23872_, _04778_);
  and (_23927_, _23926_, _23925_);
  nor (_23928_, _23927_, _23922_);
  nor (_23929_, _23928_, _03897_);
  and (_23930_, _12366_, _05437_);
  or (_23931_, _23930_, _23864_);
  and (_23932_, _23931_, _03897_);
  nor (_23933_, _23932_, _23929_);
  nor (_23934_, _23933_, _04018_);
  nor (_23935_, _08751_, _09799_);
  nor (_23936_, _23935_, _23864_);
  and (_23937_, _08750_, _05437_);
  nor (_23938_, _23937_, _23936_);
  and (_23939_, _23938_, _04018_);
  or (_23940_, _23939_, _23934_);
  and (_23941_, _23940_, _03909_);
  and (_23942_, _12244_, _05437_);
  or (_23943_, _23942_, _23864_);
  and (_23944_, _23943_, _03908_);
  or (_23946_, _23944_, _23941_);
  and (_23947_, _23946_, _04785_);
  nor (_23948_, _23937_, _23864_);
  nor (_23949_, _23948_, _04785_);
  or (_23950_, _23949_, _23947_);
  and (_23951_, _23950_, _06567_);
  nor (_23952_, _12365_, _09799_);
  or (_23953_, _23952_, _23864_);
  and (_23954_, _23953_, _03914_);
  or (_23955_, _23954_, _23951_);
  and (_23957_, _23955_, _06572_);
  nor (_23958_, _23936_, _06572_);
  or (_23959_, _23958_, _23957_);
  and (_23960_, _23959_, _03774_);
  and (_23961_, _23874_, _03773_);
  or (_23962_, _23961_, _23960_);
  and (_23963_, _23962_, _03375_);
  nor (_23964_, _23894_, _03375_);
  or (_23965_, _23964_, _23963_);
  and (_23966_, _23965_, _04060_);
  nor (_23968_, _23873_, _23864_);
  nor (_23969_, _23968_, _04060_);
  or (_23970_, _23969_, _23966_);
  or (_23971_, _23970_, _43156_);
  or (_23972_, _43152_, \oc8051_golden_model_1.IP [1]);
  and (_23973_, _23972_, _41894_);
  and (_43483_, _23973_, _23971_);
  not (_23974_, \oc8051_golden_model_1.IP [2]);
  nor (_23975_, _05437_, _23974_);
  and (_23976_, _05437_, \oc8051_golden_model_1.ACC [2]);
  nor (_23978_, _23976_, _23975_);
  nor (_23979_, _23978_, _04708_);
  nor (_23980_, _04707_, _23974_);
  or (_23981_, _23980_, _23979_);
  and (_23982_, _23981_, _04722_);
  nor (_23983_, _12471_, _09799_);
  nor (_23984_, _23983_, _23975_);
  nor (_23985_, _23984_, _04722_);
  or (_23986_, _23985_, _23982_);
  and (_23987_, _23986_, _03764_);
  nor (_23989_, _06091_, _23974_);
  and (_23990_, _12464_, _06091_);
  nor (_23991_, _23990_, _23989_);
  nor (_23992_, _23991_, _03764_);
  or (_23993_, _23992_, _23987_);
  and (_23994_, _23993_, _04733_);
  and (_23995_, _05437_, _05307_);
  nor (_23996_, _23995_, _23975_);
  nor (_23997_, _23996_, _04733_);
  or (_23998_, _23997_, _23994_);
  and (_23999_, _23998_, _03855_);
  nor (_24000_, _23978_, _03855_);
  or (_24001_, _24000_, _23999_);
  and (_24002_, _24001_, _03760_);
  and (_24003_, _12467_, _06091_);
  nor (_24004_, _24003_, _23989_);
  nor (_24005_, _24004_, _03760_);
  or (_24006_, _24005_, _03752_);
  or (_24007_, _24006_, _24002_);
  and (_24008_, _23990_, _12463_);
  or (_24010_, _23989_, _03753_);
  or (_24011_, _24010_, _24008_);
  and (_24012_, _24011_, _03747_);
  and (_24013_, _24012_, _24007_);
  nor (_24014_, _12514_, _09785_);
  nor (_24015_, _24014_, _23989_);
  nor (_24016_, _24015_, _03747_);
  or (_24017_, _24016_, _07927_);
  or (_24018_, _24017_, _24013_);
  and (_24019_, _06965_, _05437_);
  nor (_24021_, _23975_, _03738_);
  not (_24022_, _24021_);
  nor (_24023_, _24022_, _24019_);
  and (_24024_, _23996_, _08474_);
  or (_24025_, _24024_, _03455_);
  nor (_24026_, _24025_, _24023_);
  and (_24027_, _24026_, _24018_);
  nor (_24028_, _12572_, _09799_);
  nor (_24029_, _24028_, _23975_);
  nor (_24030_, _24029_, _03820_);
  or (_24032_, _24030_, _24027_);
  and (_24033_, _24032_, _04778_);
  and (_24034_, _05437_, _06495_);
  nor (_24035_, _24034_, _23975_);
  nor (_24036_, _24035_, _04778_);
  or (_24037_, _24036_, _24033_);
  and (_24038_, _24037_, _04790_);
  and (_24039_, _12586_, _05437_);
  nor (_24040_, _24039_, _23975_);
  nor (_24041_, _24040_, _04790_);
  or (_24043_, _24041_, _24038_);
  and (_24044_, _24043_, _04792_);
  and (_24045_, _08748_, _05437_);
  nor (_24046_, _24045_, _23975_);
  nor (_24047_, _24046_, _04792_);
  nor (_24048_, _24047_, _24044_);
  nor (_24049_, _24048_, _03908_);
  nor (_24050_, _23975_, _05765_);
  not (_24051_, _24050_);
  nor (_24052_, _24035_, _03909_);
  and (_24054_, _24052_, _24051_);
  nor (_24055_, _24054_, _24049_);
  nor (_24056_, _24055_, _04027_);
  nor (_24057_, _23978_, _04785_);
  and (_24058_, _24057_, _24051_);
  nor (_24059_, _24058_, _03914_);
  not (_24060_, _24059_);
  nor (_24061_, _24060_, _24056_);
  nor (_24062_, _12585_, _09799_);
  or (_24063_, _23975_, _06567_);
  nor (_24065_, _24063_, _24062_);
  or (_24066_, _24065_, _04011_);
  nor (_24067_, _24066_, _24061_);
  nor (_24068_, _08747_, _09799_);
  nor (_24069_, _24068_, _23975_);
  nor (_24070_, _24069_, _06572_);
  or (_24071_, _24070_, _24067_);
  and (_24072_, _24071_, _03774_);
  nor (_24073_, _23984_, _03774_);
  or (_24074_, _24073_, _24072_);
  and (_24076_, _24074_, _03375_);
  nor (_24077_, _24004_, _03375_);
  or (_24078_, _24077_, _24076_);
  and (_24079_, _24078_, _04060_);
  and (_24080_, _12642_, _05437_);
  nor (_24081_, _24080_, _23975_);
  nor (_24082_, _24081_, _04060_);
  or (_24083_, _24082_, _24079_);
  or (_24084_, _24083_, _43156_);
  or (_24085_, _43152_, \oc8051_golden_model_1.IP [2]);
  and (_24088_, _24085_, _41894_);
  and (_43484_, _24088_, _24084_);
  not (_24089_, \oc8051_golden_model_1.IP [3]);
  nor (_24090_, _05437_, _24089_);
  and (_24091_, _05437_, \oc8051_golden_model_1.ACC [3]);
  nor (_24092_, _24091_, _24090_);
  nor (_24093_, _24092_, _04708_);
  nor (_24094_, _04707_, _24089_);
  or (_24095_, _24094_, _24093_);
  and (_24096_, _24095_, _04722_);
  nor (_24099_, _12681_, _09799_);
  nor (_24100_, _24099_, _24090_);
  nor (_24101_, _24100_, _04722_);
  or (_24102_, _24101_, _24096_);
  and (_24103_, _24102_, _03764_);
  nor (_24104_, _06091_, _24089_);
  and (_24105_, _12674_, _06091_);
  nor (_24106_, _24105_, _24104_);
  nor (_24107_, _24106_, _03764_);
  or (_24108_, _24107_, _03848_);
  or (_24111_, _24108_, _24103_);
  and (_24112_, _05437_, _05119_);
  nor (_24113_, _24112_, _24090_);
  nand (_24114_, _24113_, _03848_);
  and (_24115_, _24114_, _24111_);
  and (_24116_, _24115_, _03855_);
  nor (_24117_, _24092_, _03855_);
  or (_24118_, _24117_, _24116_);
  and (_24119_, _24118_, _03760_);
  and (_24120_, _12667_, _06091_);
  nor (_24123_, _24120_, _24104_);
  nor (_24124_, _24123_, _03760_);
  or (_24125_, _24124_, _24119_);
  and (_24126_, _24125_, _03753_);
  nor (_24127_, _24104_, _12673_);
  nor (_24128_, _24127_, _24106_);
  and (_24129_, _24128_, _03752_);
  or (_24130_, _24129_, _24126_);
  and (_24131_, _24130_, _03747_);
  nor (_24132_, _12668_, _09785_);
  nor (_24135_, _24132_, _24104_);
  nor (_24136_, _24135_, _03747_);
  or (_24137_, _24136_, _07927_);
  or (_24138_, _24137_, _24131_);
  and (_24139_, _06964_, _05437_);
  nor (_24140_, _24090_, _03738_);
  not (_24141_, _24140_);
  nor (_24142_, _24141_, _24139_);
  and (_24143_, _24113_, _08474_);
  or (_24144_, _24143_, _03455_);
  nor (_24146_, _24144_, _24142_);
  and (_24147_, _24146_, _24138_);
  nor (_24148_, _12775_, _09799_);
  nor (_24149_, _24148_, _24090_);
  nor (_24150_, _24149_, _03820_);
  or (_24151_, _24150_, _24147_);
  and (_24152_, _24151_, _04778_);
  and (_24153_, _05437_, _06345_);
  nor (_24154_, _24153_, _24090_);
  nor (_24155_, _24154_, _04778_);
  or (_24157_, _24155_, _24152_);
  nor (_24158_, _24157_, _03897_);
  and (_24159_, _12789_, _05437_);
  or (_24160_, _24090_, _04790_);
  nor (_24161_, _24160_, _24159_);
  or (_24162_, _24161_, _04018_);
  nor (_24163_, _24162_, _24158_);
  and (_24164_, _10491_, _05437_);
  nor (_24165_, _24164_, _24090_);
  nor (_24166_, _24165_, _04792_);
  nor (_24168_, _24166_, _24163_);
  nor (_24169_, _24168_, _03908_);
  nor (_24170_, _24090_, _05622_);
  not (_24171_, _24170_);
  nor (_24172_, _24154_, _03909_);
  and (_24173_, _24172_, _24171_);
  nor (_24174_, _24173_, _24169_);
  nor (_24175_, _24174_, _04027_);
  nor (_24176_, _24092_, _04785_);
  and (_24177_, _24176_, _24171_);
  or (_24179_, _24177_, _24175_);
  and (_24180_, _24179_, _06567_);
  nor (_24181_, _12788_, _09799_);
  nor (_24182_, _24181_, _24090_);
  nor (_24183_, _24182_, _06567_);
  or (_24184_, _24183_, _24180_);
  and (_24185_, _24184_, _06572_);
  nor (_24186_, _08742_, _09799_);
  nor (_24187_, _24186_, _24090_);
  nor (_24188_, _24187_, _06572_);
  or (_24190_, _24188_, _24185_);
  and (_24191_, _24190_, _03774_);
  nor (_24192_, _24100_, _03774_);
  or (_24193_, _24192_, _24191_);
  and (_24194_, _24193_, _03375_);
  nor (_24195_, _24123_, _03375_);
  or (_24196_, _24195_, _24194_);
  and (_24197_, _24196_, _04060_);
  and (_24198_, _12848_, _05437_);
  nor (_24199_, _24198_, _24090_);
  nor (_24200_, _24199_, _04060_);
  or (_24201_, _24200_, _24197_);
  or (_24202_, _24201_, _43156_);
  or (_24203_, _43152_, \oc8051_golden_model_1.IP [3]);
  and (_24204_, _24203_, _41894_);
  and (_43485_, _24204_, _24202_);
  not (_24205_, \oc8051_golden_model_1.IP [4]);
  nor (_24206_, _05437_, _24205_);
  and (_24207_, _05437_, \oc8051_golden_model_1.ACC [4]);
  nor (_24208_, _24207_, _24206_);
  nor (_24210_, _24208_, _04708_);
  nor (_24211_, _04707_, _24205_);
  or (_24212_, _24211_, _24210_);
  and (_24213_, _24212_, _04722_);
  nor (_24214_, _12891_, _09799_);
  nor (_24215_, _24214_, _24206_);
  nor (_24216_, _24215_, _04722_);
  or (_24217_, _24216_, _24213_);
  and (_24218_, _24217_, _03764_);
  nor (_24219_, _06091_, _24205_);
  and (_24221_, _12875_, _06091_);
  nor (_24222_, _24221_, _24219_);
  nor (_24223_, _24222_, _03764_);
  or (_24224_, _24223_, _03848_);
  or (_24225_, _24224_, _24218_);
  and (_24226_, _05950_, _05437_);
  nor (_24227_, _24226_, _24206_);
  nand (_24228_, _24227_, _03848_);
  and (_24229_, _24228_, _24225_);
  and (_24230_, _24229_, _03855_);
  nor (_24232_, _24208_, _03855_);
  or (_24233_, _24232_, _24230_);
  and (_24234_, _24233_, _03760_);
  and (_24235_, _12870_, _06091_);
  nor (_24236_, _24235_, _24219_);
  nor (_24237_, _24236_, _03760_);
  or (_24238_, _24237_, _24234_);
  and (_24239_, _24238_, _03753_);
  nor (_24240_, _24219_, _12874_);
  nor (_24241_, _24240_, _24222_);
  and (_24243_, _24241_, _03752_);
  or (_24244_, _24243_, _24239_);
  and (_24245_, _24244_, _03747_);
  nor (_24246_, _12872_, _09785_);
  nor (_24247_, _24246_, _24219_);
  nor (_24248_, _24247_, _03747_);
  or (_24249_, _24248_, _07927_);
  or (_24250_, _24249_, _24245_);
  and (_24251_, _06969_, _05437_);
  nor (_24252_, _24206_, _03738_);
  not (_24254_, _24252_);
  nor (_24255_, _24254_, _24251_);
  and (_24256_, _24227_, _08474_);
  or (_24257_, _24256_, _03455_);
  nor (_24258_, _24257_, _24255_);
  and (_24259_, _24258_, _24250_);
  nor (_24260_, _12982_, _09799_);
  nor (_24261_, _24260_, _24206_);
  nor (_24262_, _24261_, _03820_);
  or (_24263_, _24262_, _24259_);
  and (_24265_, _24263_, _04778_);
  and (_24266_, _06456_, _05437_);
  nor (_24267_, _24266_, _24206_);
  nor (_24268_, _24267_, _04778_);
  or (_24269_, _24268_, _24265_);
  nor (_24270_, _24269_, _03897_);
  and (_24271_, _12997_, _05437_);
  or (_24272_, _24206_, _04790_);
  nor (_24273_, _24272_, _24271_);
  or (_24274_, _24273_, _04018_);
  nor (_24276_, _24274_, _24270_);
  and (_24277_, _08741_, _05437_);
  nor (_24278_, _24277_, _24206_);
  nor (_24279_, _24278_, _04792_);
  nor (_24280_, _24279_, _24276_);
  nor (_24281_, _24280_, _03908_);
  nor (_24282_, _24206_, _08336_);
  not (_24283_, _24282_);
  nor (_24284_, _24267_, _03909_);
  and (_24285_, _24284_, _24283_);
  nor (_24286_, _24285_, _24281_);
  nor (_24287_, _24286_, _04027_);
  nor (_24288_, _24208_, _04785_);
  and (_24289_, _24288_, _24283_);
  or (_24290_, _24289_, _24287_);
  and (_24291_, _24290_, _06567_);
  nor (_24292_, _12996_, _09799_);
  nor (_24293_, _24292_, _24206_);
  nor (_24294_, _24293_, _06567_);
  or (_24295_, _24294_, _24291_);
  and (_24297_, _24295_, _06572_);
  nor (_24298_, _08740_, _09799_);
  nor (_24299_, _24298_, _24206_);
  nor (_24300_, _24299_, _06572_);
  or (_24301_, _24300_, _24297_);
  and (_24302_, _24301_, _03774_);
  nor (_24303_, _24215_, _03774_);
  or (_24304_, _24303_, _24302_);
  and (_24305_, _24304_, _03375_);
  nor (_24306_, _24236_, _03375_);
  or (_24308_, _24306_, _24305_);
  and (_24309_, _24308_, _04060_);
  and (_24310_, _13056_, _05437_);
  nor (_24311_, _24310_, _24206_);
  nor (_24312_, _24311_, _04060_);
  or (_24313_, _24312_, _24309_);
  or (_24314_, _24313_, _43156_);
  or (_24315_, _43152_, \oc8051_golden_model_1.IP [4]);
  and (_24316_, _24315_, _41894_);
  and (_43486_, _24316_, _24314_);
  not (_24318_, \oc8051_golden_model_1.IP [5]);
  nor (_24319_, _05437_, _24318_);
  nor (_24320_, _13090_, _09799_);
  nor (_24321_, _24320_, _24319_);
  nor (_24322_, _24321_, _04722_);
  nor (_24323_, _04707_, _24318_);
  and (_24324_, _05437_, \oc8051_golden_model_1.ACC [5]);
  nor (_24325_, _24324_, _24319_);
  nor (_24326_, _24325_, _04708_);
  nor (_24327_, _24326_, _24323_);
  nor (_24329_, _24327_, _03850_);
  or (_24330_, _24329_, _03857_);
  or (_24331_, _24330_, _24322_);
  nor (_24332_, _06091_, _24318_);
  and (_24333_, _13094_, _06091_);
  nor (_24334_, _24333_, _24332_);
  and (_24335_, _24334_, _03763_);
  and (_24336_, _05857_, _05437_);
  nor (_24337_, _24336_, _24319_);
  and (_24338_, _24337_, _03848_);
  nor (_24340_, _24338_, _24335_);
  and (_24341_, _24340_, _24331_);
  and (_24342_, _24341_, _03855_);
  nor (_24343_, _24325_, _03855_);
  or (_24344_, _24343_, _24342_);
  and (_24345_, _24344_, _03760_);
  and (_24346_, _13071_, _06091_);
  nor (_24347_, _24346_, _24332_);
  nor (_24348_, _24347_, _03760_);
  or (_24349_, _24348_, _24345_);
  and (_24350_, _24349_, _03753_);
  nor (_24351_, _24332_, _13109_);
  nor (_24352_, _24351_, _24334_);
  and (_24353_, _24352_, _03752_);
  or (_24354_, _24353_, _24350_);
  and (_24355_, _24354_, _03747_);
  nor (_24356_, _13073_, _09785_);
  nor (_24357_, _24356_, _24332_);
  nor (_24358_, _24357_, _03747_);
  or (_24359_, _24358_, _07927_);
  or (_24361_, _24359_, _24355_);
  and (_24362_, _06968_, _05437_);
  nor (_24363_, _24319_, _03738_);
  not (_24364_, _24363_);
  nor (_24365_, _24364_, _24362_);
  and (_24366_, _24337_, _08474_);
  or (_24367_, _24366_, _03455_);
  nor (_24368_, _24367_, _24365_);
  and (_24369_, _24368_, _24361_);
  nor (_24370_, _13182_, _09799_);
  nor (_24372_, _24370_, _24319_);
  nor (_24373_, _24372_, _03820_);
  or (_24374_, _24373_, _24369_);
  and (_24375_, _24374_, _04778_);
  and (_24376_, _06447_, _05437_);
  nor (_24377_, _24376_, _24319_);
  nor (_24378_, _24377_, _04778_);
  or (_24379_, _24378_, _24375_);
  and (_24380_, _24379_, _04790_);
  and (_24381_, _13196_, _05437_);
  nor (_24383_, _24381_, _24319_);
  nor (_24384_, _24383_, _04790_);
  or (_24385_, _24384_, _24380_);
  and (_24386_, _24385_, _04792_);
  and (_24387_, _10493_, _05437_);
  nor (_24388_, _24387_, _24319_);
  nor (_24389_, _24388_, _04792_);
  nor (_24390_, _24389_, _24386_);
  nor (_24391_, _24390_, _03908_);
  nor (_24392_, _24319_, _08335_);
  not (_24394_, _24392_);
  nor (_24395_, _24377_, _03909_);
  and (_24396_, _24395_, _24394_);
  nor (_24397_, _24396_, _24391_);
  nor (_24398_, _24397_, _04027_);
  nor (_24399_, _24325_, _04785_);
  and (_24400_, _24399_, _24394_);
  or (_24401_, _24400_, _24398_);
  and (_24402_, _24401_, _06567_);
  nor (_24403_, _13195_, _09799_);
  nor (_24405_, _24403_, _24319_);
  nor (_24406_, _24405_, _06567_);
  or (_24407_, _24406_, _24402_);
  and (_24408_, _24407_, _06572_);
  nor (_24409_, _08738_, _09799_);
  nor (_24410_, _24409_, _24319_);
  nor (_24411_, _24410_, _06572_);
  or (_24412_, _24411_, _24408_);
  and (_24413_, _24412_, _03774_);
  nor (_24414_, _24321_, _03774_);
  or (_24416_, _24414_, _24413_);
  and (_24417_, _24416_, _03375_);
  nor (_24418_, _24347_, _03375_);
  or (_24419_, _24418_, _24417_);
  and (_24420_, _24419_, _04060_);
  and (_24421_, _13255_, _05437_);
  nor (_24422_, _24421_, _24319_);
  nor (_24423_, _24422_, _04060_);
  or (_24424_, _24423_, _24420_);
  or (_24425_, _24424_, _43156_);
  or (_24427_, _43152_, \oc8051_golden_model_1.IP [5]);
  and (_24428_, _24427_, _41894_);
  and (_43487_, _24428_, _24425_);
  not (_24429_, \oc8051_golden_model_1.IP [6]);
  nor (_24430_, _05437_, _24429_);
  and (_24431_, _05437_, \oc8051_golden_model_1.ACC [6]);
  nor (_24432_, _24431_, _24430_);
  nor (_24433_, _24432_, _04708_);
  nor (_24434_, _04707_, _24429_);
  or (_24435_, _24434_, _24433_);
  and (_24437_, _24435_, _04722_);
  nor (_24438_, _13293_, _09799_);
  nor (_24439_, _24438_, _24430_);
  nor (_24440_, _24439_, _04722_);
  or (_24441_, _24440_, _24437_);
  and (_24442_, _24441_, _03764_);
  nor (_24443_, _06091_, _24429_);
  and (_24444_, _13297_, _06091_);
  nor (_24445_, _24444_, _24443_);
  nor (_24446_, _24445_, _03764_);
  or (_24448_, _24446_, _03848_);
  or (_24449_, _24448_, _24442_);
  and (_24450_, _06065_, _05437_);
  nor (_24451_, _24450_, _24430_);
  nand (_24452_, _24451_, _03848_);
  and (_24453_, _24452_, _24449_);
  and (_24454_, _24453_, _03855_);
  nor (_24455_, _24432_, _03855_);
  or (_24456_, _24455_, _24454_);
  and (_24457_, _24456_, _03760_);
  and (_24459_, _13277_, _06091_);
  nor (_24460_, _24459_, _24443_);
  nor (_24461_, _24460_, _03760_);
  or (_24462_, _24461_, _24457_);
  and (_24463_, _24462_, _03753_);
  nor (_24464_, _24443_, _13312_);
  nor (_24465_, _24464_, _24445_);
  and (_24466_, _24465_, _03752_);
  or (_24467_, _24466_, _24463_);
  and (_24468_, _24467_, _03747_);
  nor (_24470_, _13279_, _09785_);
  nor (_24471_, _24470_, _24443_);
  nor (_24472_, _24471_, _03747_);
  or (_24473_, _24472_, _07927_);
  or (_24474_, _24473_, _24468_);
  and (_24475_, _06641_, _05437_);
  nor (_24476_, _24430_, _03738_);
  not (_24477_, _24476_);
  nor (_24478_, _24477_, _24475_);
  and (_24479_, _24451_, _08474_);
  or (_24481_, _24479_, _03455_);
  nor (_24482_, _24481_, _24478_);
  and (_24483_, _24482_, _24474_);
  nor (_24484_, _13387_, _09799_);
  nor (_24485_, _24484_, _24430_);
  nor (_24486_, _24485_, _03820_);
  or (_24487_, _24486_, _24483_);
  and (_24488_, _24487_, _04778_);
  and (_24489_, _13394_, _05437_);
  nor (_24490_, _24489_, _24430_);
  nor (_24492_, _24490_, _04778_);
  or (_24493_, _24492_, _24488_);
  nor (_24494_, _24493_, _03897_);
  and (_24495_, _13402_, _05437_);
  or (_24496_, _24430_, _04790_);
  nor (_24497_, _24496_, _24495_);
  or (_24498_, _24497_, _04018_);
  nor (_24499_, _24498_, _24494_);
  and (_24500_, _08736_, _05437_);
  nor (_24501_, _24500_, _24430_);
  nor (_24504_, _24501_, _04792_);
  nor (_24505_, _24504_, _24499_);
  nor (_24506_, _24505_, _03908_);
  nor (_24507_, _24430_, _08322_);
  not (_24508_, _24507_);
  nor (_24509_, _24490_, _03909_);
  and (_24510_, _24509_, _24508_);
  nor (_24511_, _24510_, _24506_);
  nor (_24512_, _24511_, _04027_);
  nor (_24513_, _24432_, _04785_);
  and (_24515_, _24513_, _24508_);
  or (_24516_, _24515_, _24512_);
  and (_24517_, _24516_, _06567_);
  nor (_24518_, _13401_, _09799_);
  nor (_24519_, _24518_, _24430_);
  nor (_24520_, _24519_, _06567_);
  or (_24521_, _24520_, _24517_);
  and (_24522_, _24521_, _06572_);
  nor (_24523_, _08735_, _09799_);
  nor (_24524_, _24523_, _24430_);
  nor (_24526_, _24524_, _06572_);
  or (_24527_, _24526_, _24522_);
  and (_24528_, _24527_, _03774_);
  nor (_24529_, _24439_, _03774_);
  or (_24530_, _24529_, _24528_);
  and (_24531_, _24530_, _03375_);
  nor (_24532_, _24460_, _03375_);
  or (_24533_, _24532_, _24531_);
  and (_24534_, _24533_, _04060_);
  nor (_24535_, _13460_, _09799_);
  nor (_24537_, _24535_, _24430_);
  nor (_24538_, _24537_, _04060_);
  or (_24539_, _24538_, _24534_);
  or (_24540_, _24539_, _43156_);
  or (_24541_, _43152_, \oc8051_golden_model_1.IP [6]);
  and (_24542_, _24541_, _41894_);
  and (_43488_, _24542_, _24540_);
  not (_24543_, \oc8051_golden_model_1.DPL [0]);
  nor (_24544_, _43152_, _24543_);
  and (_24545_, _06962_, _05513_);
  nor (_24547_, _05513_, _24543_);
  or (_24548_, _24547_, _03738_);
  or (_24549_, _24548_, _24545_);
  and (_24550_, _05513_, _04700_);
  or (_24551_, _24550_, _24547_);
  or (_24552_, _24551_, _07925_);
  and (_24553_, _05513_, \oc8051_golden_model_1.ACC [0]);
  or (_24554_, _24553_, _24547_);
  or (_24555_, _24554_, _03855_);
  and (_24556_, _05716_, _05513_);
  or (_24558_, _24556_, _24547_);
  or (_24559_, _24558_, _04722_);
  and (_24560_, _24554_, _04707_);
  nor (_24561_, _04707_, _24543_);
  or (_24562_, _24561_, _03850_);
  or (_24563_, _24562_, _24560_);
  and (_24564_, _24563_, _04733_);
  and (_24565_, _24564_, _24559_);
  and (_24566_, _24551_, _03848_);
  or (_24567_, _24566_, _03854_);
  or (_24569_, _24567_, _24565_);
  and (_24570_, _24569_, _24555_);
  or (_24571_, _24570_, _09878_);
  nand (_24572_, _09878_, \oc8051_golden_model_1.DPL [0]);
  and (_24573_, _24572_, _09861_);
  and (_24574_, _24573_, _24571_);
  nor (_24575_, _04382_, _09861_);
  or (_24576_, _24575_, _07927_);
  or (_24577_, _24576_, _24574_);
  and (_24578_, _24577_, _24552_);
  and (_24580_, _24578_, _24549_);
  or (_24581_, _24580_, _03455_);
  nor (_24582_, _12164_, _09905_);
  or (_24583_, _24547_, _03820_);
  or (_24584_, _24583_, _24582_);
  and (_24585_, _24584_, _04778_);
  and (_24586_, _24585_, _24581_);
  and (_24587_, _05513_, _06479_);
  or (_24588_, _24587_, _24547_);
  and (_24589_, _24588_, _03903_);
  or (_24591_, _24589_, _03897_);
  or (_24592_, _24591_, _24586_);
  and (_24593_, _12178_, _05513_);
  or (_24594_, _24593_, _24547_);
  or (_24595_, _24594_, _04790_);
  and (_24596_, _24595_, _04792_);
  and (_24597_, _24596_, _24592_);
  nor (_24598_, _10488_, _09905_);
  or (_24599_, _24598_, _24547_);
  nand (_24600_, _08753_, _05513_);
  and (_24602_, _24600_, _04018_);
  and (_24603_, _24602_, _24599_);
  or (_24604_, _24603_, _24597_);
  and (_24605_, _24604_, _03909_);
  nand (_24606_, _24588_, _03908_);
  nor (_24607_, _24606_, _24556_);
  or (_24608_, _24607_, _04027_);
  or (_24609_, _24608_, _24605_);
  nor (_24610_, _24547_, _04785_);
  nand (_24611_, _24610_, _24600_);
  and (_24613_, _24611_, _24609_);
  or (_24614_, _24613_, _03914_);
  nor (_24615_, _12177_, _09905_);
  or (_24616_, _24547_, _06567_);
  or (_24617_, _24616_, _24615_);
  and (_24618_, _24617_, _06572_);
  and (_24619_, _24618_, _24614_);
  and (_24620_, _24599_, _04011_);
  or (_24621_, _24620_, _17157_);
  or (_24622_, _24621_, _24619_);
  or (_24624_, _24558_, _04144_);
  and (_24625_, _24624_, _43152_);
  and (_24626_, _24625_, _24622_);
  or (_24627_, _24626_, _24544_);
  and (_43491_, _24627_, _41894_);
  not (_24628_, \oc8051_golden_model_1.DPL [1]);
  nor (_24629_, _43152_, _24628_);
  nor (_24630_, _05513_, _24628_);
  and (_24631_, _05513_, _04900_);
  or (_24632_, _24631_, _24630_);
  or (_24634_, _24632_, _04733_);
  or (_24635_, _05513_, \oc8051_golden_model_1.DPL [1]);
  and (_24636_, _12262_, _05513_);
  not (_24637_, _24636_);
  and (_24638_, _24637_, _24635_);
  and (_24639_, _24638_, _03850_);
  nor (_24640_, _04707_, _24628_);
  and (_24641_, _05513_, \oc8051_golden_model_1.ACC [1]);
  or (_24642_, _24641_, _24630_);
  and (_24643_, _24642_, _04707_);
  or (_24645_, _24643_, _24640_);
  and (_24646_, _24645_, _04722_);
  or (_24647_, _24646_, _03848_);
  or (_24648_, _24647_, _24639_);
  and (_24649_, _24648_, _24634_);
  or (_24650_, _24649_, _03854_);
  or (_24651_, _24642_, _03855_);
  and (_24652_, _24651_, _09879_);
  and (_24653_, _24652_, _24650_);
  nor (_24654_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_24656_, _24654_, _09883_);
  and (_24657_, _24656_, _09878_);
  or (_24658_, _24657_, _24653_);
  and (_24659_, _24658_, _09861_);
  nor (_24660_, _04595_, _09861_);
  or (_24661_, _24660_, _07927_);
  or (_24662_, _24661_, _24659_);
  and (_24663_, _06961_, _05513_);
  or (_24664_, _24630_, _03738_);
  or (_24665_, _24664_, _24663_);
  or (_24667_, _24632_, _07925_);
  and (_24668_, _24667_, _03820_);
  and (_24669_, _24668_, _24665_);
  and (_24670_, _24669_, _24662_);
  nor (_24671_, _12352_, _09905_);
  or (_24672_, _24671_, _24630_);
  and (_24673_, _24672_, _03455_);
  or (_24674_, _24673_, _24670_);
  and (_24675_, _24674_, _04778_);
  nand (_24676_, _05513_, _04595_);
  and (_24678_, _24635_, _03903_);
  and (_24679_, _24678_, _24676_);
  or (_24680_, _24679_, _24675_);
  and (_24681_, _24680_, _04790_);
  or (_24682_, _12366_, _09905_);
  and (_24683_, _24635_, _03897_);
  and (_24684_, _24683_, _24682_);
  or (_24685_, _24684_, _04018_);
  or (_24686_, _24685_, _24681_);
  nor (_24687_, _08751_, _09905_);
  or (_24689_, _24687_, _24630_);
  nand (_24690_, _08750_, _05513_);
  and (_24691_, _24690_, _24689_);
  or (_24692_, _24691_, _04792_);
  and (_24693_, _24692_, _03909_);
  and (_24694_, _24693_, _24686_);
  or (_24695_, _12244_, _09905_);
  and (_24696_, _24635_, _03908_);
  and (_24697_, _24696_, _24695_);
  or (_24698_, _24697_, _04027_);
  or (_24700_, _24698_, _24694_);
  nor (_24701_, _24630_, _04785_);
  nand (_24702_, _24701_, _24690_);
  and (_24703_, _24702_, _06567_);
  and (_24704_, _24703_, _24700_);
  or (_24705_, _24676_, _08366_);
  and (_24706_, _24635_, _03914_);
  and (_24707_, _24706_, _24705_);
  or (_24708_, _24707_, _04011_);
  or (_24709_, _24708_, _24704_);
  or (_24711_, _24689_, _06572_);
  and (_24712_, _24711_, _03774_);
  and (_24713_, _24712_, _24709_);
  and (_24714_, _24638_, _03773_);
  or (_24715_, _24714_, _03772_);
  or (_24716_, _24715_, _24713_);
  or (_24717_, _24630_, _04060_);
  or (_24718_, _24717_, _24636_);
  and (_24719_, _24718_, _43152_);
  and (_24720_, _24719_, _24716_);
  or (_24722_, _24720_, _24629_);
  and (_43492_, _24722_, _41894_);
  or (_24723_, _43152_, \oc8051_golden_model_1.DPL [2]);
  and (_24724_, _24723_, _41894_);
  and (_24725_, _09905_, \oc8051_golden_model_1.DPL [2]);
  and (_24726_, _05513_, _06495_);
  or (_24727_, _24726_, _24725_);
  or (_24728_, _24727_, _04778_);
  nor (_24729_, _09883_, \oc8051_golden_model_1.DPL [2]);
  nor (_24730_, _24729_, _09884_);
  and (_24732_, _24730_, _09878_);
  nor (_24733_, _12471_, _09905_);
  or (_24734_, _24733_, _24725_);
  or (_24735_, _24734_, _04722_);
  and (_24736_, _05513_, \oc8051_golden_model_1.ACC [2]);
  or (_24737_, _24736_, _24725_);
  and (_24738_, _24737_, _04707_);
  and (_24739_, _04708_, \oc8051_golden_model_1.DPL [2]);
  or (_24740_, _24739_, _03850_);
  or (_24741_, _24740_, _24738_);
  and (_24743_, _24741_, _04733_);
  and (_24744_, _24743_, _24735_);
  and (_24745_, _05513_, _05307_);
  or (_24746_, _24745_, _24725_);
  and (_24747_, _24746_, _03848_);
  or (_24748_, _24747_, _03854_);
  or (_24749_, _24748_, _24744_);
  or (_24750_, _24737_, _03855_);
  and (_24751_, _24750_, _09879_);
  and (_24752_, _24751_, _24749_);
  or (_24754_, _24752_, _24732_);
  and (_24755_, _24754_, _09861_);
  nor (_24756_, _04180_, _09861_);
  or (_24757_, _24756_, _07927_);
  or (_24758_, _24757_, _24755_);
  and (_24759_, _06965_, _05513_);
  or (_24760_, _24725_, _03738_);
  or (_24761_, _24760_, _24759_);
  or (_24762_, _24746_, _07925_);
  and (_24763_, _24762_, _03820_);
  and (_24765_, _24763_, _24761_);
  and (_24766_, _24765_, _24758_);
  nor (_24767_, _12572_, _09905_);
  or (_24768_, _24767_, _24725_);
  and (_24769_, _24768_, _03455_);
  or (_24770_, _24769_, _03903_);
  or (_24771_, _24770_, _24766_);
  and (_24772_, _24771_, _24728_);
  or (_24773_, _24772_, _03897_);
  and (_24774_, _12586_, _05513_);
  or (_24776_, _24774_, _24725_);
  or (_24777_, _24776_, _04790_);
  and (_24778_, _24777_, _04792_);
  and (_24779_, _24778_, _24773_);
  and (_24780_, _08748_, _05513_);
  or (_24781_, _24780_, _24725_);
  and (_24782_, _24781_, _04018_);
  or (_24783_, _24782_, _24779_);
  and (_24784_, _24783_, _03909_);
  or (_24785_, _24725_, _05765_);
  and (_24787_, _24727_, _03908_);
  and (_24788_, _24787_, _24785_);
  or (_24789_, _24788_, _24784_);
  and (_24790_, _24789_, _04785_);
  and (_24791_, _24737_, _04027_);
  and (_24792_, _24791_, _24785_);
  or (_24793_, _24792_, _03914_);
  or (_24794_, _24793_, _24790_);
  nor (_24795_, _12585_, _09905_);
  or (_24796_, _24725_, _06567_);
  or (_24798_, _24796_, _24795_);
  and (_24799_, _24798_, _06572_);
  and (_24800_, _24799_, _24794_);
  nor (_24801_, _08747_, _09905_);
  or (_24802_, _24801_, _24725_);
  and (_24803_, _24802_, _04011_);
  or (_24804_, _24803_, _03773_);
  or (_24805_, _24804_, _24800_);
  or (_24806_, _24734_, _03774_);
  and (_24807_, _24806_, _04060_);
  and (_24809_, _24807_, _24805_);
  and (_24810_, _12642_, _05513_);
  or (_24811_, _24810_, _24725_);
  and (_24812_, _24811_, _03772_);
  or (_24813_, _24812_, _43156_);
  or (_24814_, _24813_, _24809_);
  and (_43493_, _24814_, _24724_);
  or (_24815_, _43152_, \oc8051_golden_model_1.DPL [3]);
  and (_24816_, _24815_, _41894_);
  and (_24817_, _09905_, \oc8051_golden_model_1.DPL [3]);
  and (_24819_, _05513_, _06345_);
  or (_24820_, _24819_, _24817_);
  or (_24821_, _24820_, _04778_);
  nor (_24822_, _09884_, \oc8051_golden_model_1.DPL [3]);
  nor (_24823_, _24822_, _09885_);
  and (_24824_, _24823_, _09878_);
  nor (_24825_, _12681_, _09905_);
  or (_24826_, _24825_, _24817_);
  or (_24827_, _24826_, _04722_);
  and (_24828_, _05513_, \oc8051_golden_model_1.ACC [3]);
  or (_24830_, _24828_, _24817_);
  and (_24831_, _24830_, _04707_);
  and (_24832_, _04708_, \oc8051_golden_model_1.DPL [3]);
  or (_24833_, _24832_, _03850_);
  or (_24834_, _24833_, _24831_);
  and (_24835_, _24834_, _04733_);
  and (_24836_, _24835_, _24827_);
  and (_24837_, _05513_, _05119_);
  or (_24838_, _24837_, _24817_);
  and (_24839_, _24838_, _03848_);
  or (_24841_, _24839_, _03854_);
  or (_24842_, _24841_, _24836_);
  or (_24843_, _24830_, _03855_);
  and (_24844_, _24843_, _09879_);
  and (_24845_, _24844_, _24842_);
  or (_24846_, _24845_, _24824_);
  and (_24847_, _24846_, _09861_);
  nor (_24848_, _04005_, _09861_);
  or (_24849_, _24848_, _07927_);
  or (_24850_, _24849_, _24847_);
  and (_24852_, _06964_, _05513_);
  or (_24853_, _24817_, _03738_);
  or (_24854_, _24853_, _24852_);
  or (_24855_, _24838_, _07925_);
  and (_24856_, _24855_, _03820_);
  and (_24857_, _24856_, _24854_);
  and (_24858_, _24857_, _24850_);
  nor (_24859_, _12775_, _09905_);
  or (_24860_, _24859_, _24817_);
  and (_24861_, _24860_, _03455_);
  or (_24863_, _24861_, _03903_);
  or (_24864_, _24863_, _24858_);
  and (_24865_, _24864_, _24821_);
  or (_24866_, _24865_, _03897_);
  and (_24867_, _12789_, _05513_);
  or (_24868_, _24867_, _24817_);
  or (_24869_, _24868_, _04790_);
  and (_24870_, _24869_, _04792_);
  and (_24871_, _24870_, _24866_);
  and (_24872_, _10491_, _05513_);
  or (_24874_, _24872_, _24817_);
  and (_24875_, _24874_, _04018_);
  or (_24876_, _24875_, _24871_);
  and (_24877_, _24876_, _03909_);
  or (_24878_, _24817_, _05622_);
  and (_24879_, _24820_, _03908_);
  and (_24880_, _24879_, _24878_);
  or (_24881_, _24880_, _24877_);
  and (_24882_, _24881_, _04785_);
  and (_24883_, _24830_, _04027_);
  and (_24885_, _24883_, _24878_);
  or (_24886_, _24885_, _03914_);
  or (_24887_, _24886_, _24882_);
  nor (_24888_, _12788_, _09905_);
  or (_24889_, _24817_, _06567_);
  or (_24890_, _24889_, _24888_);
  and (_24891_, _24890_, _06572_);
  and (_24892_, _24891_, _24887_);
  nor (_24893_, _08742_, _09905_);
  or (_24894_, _24893_, _24817_);
  and (_24896_, _24894_, _04011_);
  or (_24897_, _24896_, _03773_);
  or (_24898_, _24897_, _24892_);
  or (_24899_, _24826_, _03774_);
  and (_24900_, _24899_, _04060_);
  and (_24901_, _24900_, _24898_);
  and (_24902_, _12848_, _05513_);
  or (_24903_, _24902_, _24817_);
  and (_24904_, _24903_, _03772_);
  or (_24905_, _24904_, _43156_);
  or (_24907_, _24905_, _24901_);
  and (_43494_, _24907_, _24816_);
  or (_24908_, _43152_, \oc8051_golden_model_1.DPL [4]);
  and (_24909_, _24908_, _41894_);
  and (_24910_, _09905_, \oc8051_golden_model_1.DPL [4]);
  and (_24911_, _06456_, _05513_);
  or (_24912_, _24911_, _24910_);
  or (_24913_, _24912_, _04778_);
  nor (_24914_, _12891_, _09905_);
  or (_24915_, _24914_, _24910_);
  or (_24917_, _24915_, _04722_);
  and (_24918_, _05513_, \oc8051_golden_model_1.ACC [4]);
  or (_24919_, _24918_, _24910_);
  and (_24920_, _24919_, _04707_);
  and (_24921_, _04708_, \oc8051_golden_model_1.DPL [4]);
  or (_24922_, _24921_, _03850_);
  or (_24923_, _24922_, _24920_);
  and (_24924_, _24923_, _04733_);
  and (_24925_, _24924_, _24917_);
  and (_24926_, _05950_, _05513_);
  or (_24928_, _24926_, _24910_);
  and (_24929_, _24928_, _03848_);
  or (_24930_, _24929_, _03854_);
  or (_24931_, _24930_, _24925_);
  or (_24932_, _24919_, _03855_);
  and (_24933_, _24932_, _09879_);
  and (_24934_, _24933_, _24931_);
  nor (_24935_, _09885_, \oc8051_golden_model_1.DPL [4]);
  nor (_24936_, _24935_, _09886_);
  and (_24937_, _24936_, _09878_);
  or (_24939_, _24937_, _24934_);
  and (_24940_, _24939_, _09861_);
  nor (_24941_, _06442_, _09861_);
  or (_24942_, _24941_, _07927_);
  or (_24943_, _24942_, _24940_);
  and (_24944_, _06969_, _05513_);
  or (_24945_, _24910_, _03738_);
  or (_24946_, _24945_, _24944_);
  or (_24947_, _24928_, _07925_);
  and (_24948_, _24947_, _03820_);
  and (_24950_, _24948_, _24946_);
  and (_24951_, _24950_, _24943_);
  nor (_24952_, _12982_, _09905_);
  or (_24953_, _24952_, _24910_);
  and (_24954_, _24953_, _03455_);
  or (_24955_, _24954_, _03903_);
  or (_24956_, _24955_, _24951_);
  and (_24957_, _24956_, _24913_);
  or (_24958_, _24957_, _03897_);
  and (_24959_, _12997_, _05513_);
  or (_24961_, _24910_, _04790_);
  or (_24962_, _24961_, _24959_);
  and (_24963_, _24962_, _04792_);
  and (_24964_, _24963_, _24958_);
  and (_24965_, _08741_, _05513_);
  or (_24966_, _24965_, _24910_);
  and (_24967_, _24966_, _04018_);
  or (_24968_, _24967_, _24964_);
  and (_24969_, _24968_, _03909_);
  or (_24970_, _24910_, _08336_);
  and (_24972_, _24912_, _03908_);
  and (_24973_, _24972_, _24970_);
  or (_24974_, _24973_, _24969_);
  and (_24975_, _24974_, _04785_);
  and (_24976_, _24919_, _04027_);
  and (_24977_, _24976_, _24970_);
  or (_24978_, _24977_, _03914_);
  or (_24979_, _24978_, _24975_);
  nor (_24980_, _12996_, _09905_);
  or (_24981_, _24910_, _06567_);
  or (_24982_, _24981_, _24980_);
  and (_24983_, _24982_, _06572_);
  and (_24984_, _24983_, _24979_);
  nor (_24985_, _08740_, _09905_);
  or (_24986_, _24985_, _24910_);
  and (_24987_, _24986_, _04011_);
  or (_24988_, _24987_, _03773_);
  or (_24989_, _24988_, _24984_);
  or (_24990_, _24915_, _03774_);
  and (_24991_, _24990_, _04060_);
  and (_24994_, _24991_, _24989_);
  and (_24995_, _13056_, _05513_);
  or (_24996_, _24995_, _24910_);
  and (_24997_, _24996_, _03772_);
  or (_24998_, _24997_, _43156_);
  or (_24999_, _24998_, _24994_);
  and (_43495_, _24999_, _24909_);
  and (_25000_, _43156_, \oc8051_golden_model_1.DPL [5]);
  and (_25001_, _09905_, \oc8051_golden_model_1.DPL [5]);
  and (_25002_, _06447_, _05513_);
  or (_25004_, _25002_, _25001_);
  or (_25005_, _25004_, _04778_);
  nor (_25006_, _13090_, _09905_);
  or (_25007_, _25006_, _25001_);
  or (_25008_, _25007_, _04722_);
  and (_25009_, _05513_, \oc8051_golden_model_1.ACC [5]);
  or (_25010_, _25009_, _25001_);
  and (_25011_, _25010_, _04707_);
  and (_25012_, _04708_, \oc8051_golden_model_1.DPL [5]);
  or (_25013_, _25012_, _03850_);
  or (_25015_, _25013_, _25011_);
  and (_25016_, _25015_, _04733_);
  and (_25017_, _25016_, _25008_);
  and (_25018_, _05857_, _05513_);
  or (_25019_, _25018_, _25001_);
  and (_25020_, _25019_, _03848_);
  or (_25021_, _25020_, _03854_);
  or (_25022_, _25021_, _25017_);
  or (_25023_, _25010_, _03855_);
  and (_25024_, _25023_, _09879_);
  and (_25025_, _25024_, _25022_);
  nor (_25026_, _09886_, \oc8051_golden_model_1.DPL [5]);
  nor (_25027_, _25026_, _09887_);
  and (_25028_, _25027_, _09878_);
  or (_25029_, _25028_, _25025_);
  and (_25030_, _25029_, _09861_);
  nor (_25031_, _06411_, _09861_);
  or (_25032_, _25031_, _07927_);
  or (_25033_, _25032_, _25030_);
  and (_25034_, _06968_, _05513_);
  or (_25037_, _25001_, _03738_);
  or (_25038_, _25037_, _25034_);
  or (_25039_, _25019_, _07925_);
  and (_25040_, _25039_, _03820_);
  and (_25041_, _25040_, _25038_);
  and (_25042_, _25041_, _25033_);
  nor (_25043_, _13182_, _09905_);
  or (_25044_, _25043_, _25001_);
  and (_25045_, _25044_, _03455_);
  or (_25046_, _25045_, _03903_);
  or (_25048_, _25046_, _25042_);
  and (_25049_, _25048_, _25005_);
  or (_25050_, _25049_, _03897_);
  and (_25051_, _13196_, _05513_);
  or (_25052_, _25001_, _04790_);
  or (_25053_, _25052_, _25051_);
  and (_25054_, _25053_, _04792_);
  and (_25055_, _25054_, _25050_);
  and (_25056_, _10493_, _05513_);
  or (_25057_, _25056_, _25001_);
  and (_25058_, _25057_, _04018_);
  or (_25059_, _25058_, _25055_);
  and (_25060_, _25059_, _03909_);
  or (_25061_, _25001_, _08335_);
  and (_25062_, _25004_, _03908_);
  and (_25063_, _25062_, _25061_);
  or (_25064_, _25063_, _25060_);
  and (_25065_, _25064_, _04785_);
  and (_25066_, _25010_, _04027_);
  and (_25067_, _25066_, _25061_);
  or (_25070_, _25067_, _03914_);
  or (_25071_, _25070_, _25065_);
  nor (_25072_, _13195_, _09905_);
  or (_25073_, _25001_, _06567_);
  or (_25074_, _25073_, _25072_);
  and (_25075_, _25074_, _06572_);
  and (_25076_, _25075_, _25071_);
  nor (_25077_, _08738_, _09905_);
  or (_25078_, _25077_, _25001_);
  and (_25079_, _25078_, _04011_);
  or (_25081_, _25079_, _25076_);
  and (_25082_, _25081_, _03774_);
  and (_25083_, _25007_, _03773_);
  or (_25084_, _25083_, _03772_);
  or (_25085_, _25084_, _25082_);
  and (_25086_, _13255_, _05513_);
  or (_25087_, _25001_, _04060_);
  or (_25088_, _25087_, _25086_);
  and (_25089_, _25088_, _43152_);
  and (_25090_, _25089_, _25085_);
  or (_25092_, _25090_, _25000_);
  and (_43496_, _25092_, _41894_);
  or (_25093_, _43152_, \oc8051_golden_model_1.DPL [6]);
  and (_25094_, _25093_, _41894_);
  and (_25095_, _09905_, \oc8051_golden_model_1.DPL [6]);
  and (_25096_, _13394_, _05513_);
  or (_25097_, _25096_, _25095_);
  or (_25098_, _25097_, _04778_);
  nor (_25099_, _13293_, _09905_);
  or (_25100_, _25099_, _25095_);
  or (_25102_, _25100_, _04722_);
  and (_25103_, _05513_, \oc8051_golden_model_1.ACC [6]);
  or (_25104_, _25103_, _25095_);
  and (_25105_, _25104_, _04707_);
  and (_25106_, _04708_, \oc8051_golden_model_1.DPL [6]);
  or (_25107_, _25106_, _03850_);
  or (_25108_, _25107_, _25105_);
  and (_25109_, _25108_, _04733_);
  and (_25110_, _25109_, _25102_);
  and (_25111_, _06065_, _05513_);
  or (_25112_, _25111_, _25095_);
  and (_25113_, _25112_, _03848_);
  or (_25114_, _25113_, _03854_);
  or (_25115_, _25114_, _25110_);
  or (_25116_, _25104_, _03855_);
  and (_25117_, _25116_, _09879_);
  and (_25118_, _25117_, _25115_);
  nor (_25119_, _09887_, \oc8051_golden_model_1.DPL [6]);
  nor (_25120_, _25119_, _09888_);
  and (_25121_, _25120_, _09878_);
  or (_25124_, _25121_, _25118_);
  and (_25125_, _25124_, _09861_);
  nor (_25126_, _06379_, _09861_);
  or (_25127_, _25126_, _07927_);
  or (_25128_, _25127_, _25125_);
  and (_25129_, _06641_, _05513_);
  or (_25130_, _25095_, _03738_);
  or (_25131_, _25130_, _25129_);
  or (_25132_, _25112_, _07925_);
  and (_25133_, _25132_, _03820_);
  and (_25135_, _25133_, _25131_);
  and (_25136_, _25135_, _25128_);
  nor (_25137_, _13387_, _09905_);
  or (_25138_, _25137_, _25095_);
  and (_25139_, _25138_, _03455_);
  or (_25140_, _25139_, _03903_);
  or (_25141_, _25140_, _25136_);
  and (_25142_, _25141_, _25098_);
  or (_25143_, _25142_, _03897_);
  and (_25144_, _13402_, _05513_);
  or (_25146_, _25144_, _25095_);
  or (_25147_, _25146_, _04790_);
  and (_25148_, _25147_, _04792_);
  and (_25149_, _25148_, _25143_);
  and (_25150_, _08736_, _05513_);
  or (_25151_, _25150_, _25095_);
  and (_25152_, _25151_, _04018_);
  or (_25153_, _25152_, _25149_);
  and (_25154_, _25153_, _03909_);
  or (_25155_, _25095_, _08322_);
  and (_25157_, _25097_, _03908_);
  and (_25158_, _25157_, _25155_);
  or (_25159_, _25158_, _25154_);
  and (_25160_, _25159_, _04785_);
  and (_25161_, _25104_, _04027_);
  and (_25162_, _25161_, _25155_);
  or (_25163_, _25162_, _03914_);
  or (_25164_, _25163_, _25160_);
  nor (_25165_, _13401_, _09905_);
  or (_25166_, _25095_, _06567_);
  or (_25168_, _25166_, _25165_);
  and (_25169_, _25168_, _06572_);
  and (_25170_, _25169_, _25164_);
  nor (_25171_, _08735_, _09905_);
  or (_25172_, _25171_, _25095_);
  and (_25173_, _25172_, _04011_);
  or (_25174_, _25173_, _03773_);
  or (_25175_, _25174_, _25170_);
  or (_25176_, _25100_, _03774_);
  and (_25177_, _25176_, _04060_);
  and (_25179_, _25177_, _25175_);
  nor (_25180_, _13460_, _09905_);
  or (_25181_, _25180_, _25095_);
  and (_25182_, _25181_, _03772_);
  or (_25183_, _25182_, _43156_);
  or (_25184_, _25183_, _25179_);
  and (_43497_, _25184_, _25094_);
  nor (_25185_, _43152_, _10585_);
  nand (_25186_, _08753_, _05509_);
  nor (_25187_, _05509_, _10585_);
  nor (_25189_, _25187_, _04785_);
  nand (_25190_, _25189_, _25186_);
  and (_25191_, _06962_, _05509_);
  or (_25192_, _25187_, _03738_);
  or (_25193_, _25192_, _25191_);
  and (_25194_, _05509_, _04700_);
  or (_25195_, _25194_, _25187_);
  or (_25196_, _25195_, _07925_);
  nor (_25197_, _09890_, \oc8051_golden_model_1.DPH [0]);
  nor (_25198_, _25197_, _09977_);
  and (_25200_, _25198_, _09878_);
  and (_25201_, _05716_, _05509_);
  or (_25202_, _25201_, _25187_);
  or (_25203_, _25202_, _04722_);
  and (_25204_, _05509_, \oc8051_golden_model_1.ACC [0]);
  or (_25205_, _25204_, _25187_);
  and (_25206_, _25205_, _04707_);
  nor (_25207_, _04707_, _10585_);
  or (_25208_, _25207_, _03850_);
  or (_25209_, _25208_, _25206_);
  and (_25211_, _25209_, _04733_);
  and (_25212_, _25211_, _25203_);
  and (_25213_, _25195_, _03848_);
  or (_25214_, _25213_, _03854_);
  or (_25215_, _25214_, _25212_);
  or (_25216_, _25205_, _03855_);
  and (_25217_, _25216_, _09879_);
  and (_25218_, _25217_, _25215_);
  or (_25219_, _25218_, _25200_);
  and (_25220_, _25219_, _09861_);
  nor (_25222_, _03715_, _09861_);
  or (_25223_, _25222_, _07927_);
  or (_25224_, _25223_, _25220_);
  and (_25225_, _25224_, _25196_);
  and (_25226_, _25225_, _25193_);
  or (_25227_, _25226_, _03455_);
  nor (_25228_, _12164_, _10000_);
  or (_25229_, _25187_, _03820_);
  or (_25230_, _25229_, _25228_);
  and (_25231_, _25230_, _04778_);
  and (_25233_, _25231_, _25227_);
  and (_25234_, _05509_, _06479_);
  or (_25235_, _25234_, _25187_);
  and (_25236_, _25235_, _03903_);
  or (_25237_, _25236_, _03897_);
  or (_25238_, _25237_, _25233_);
  and (_25239_, _12178_, _05509_);
  or (_25240_, _25239_, _25187_);
  or (_25241_, _25240_, _04790_);
  and (_25242_, _25241_, _04792_);
  and (_25243_, _25242_, _25238_);
  nor (_25244_, _10488_, _10000_);
  or (_25245_, _25244_, _25187_);
  and (_25246_, _25186_, _04018_);
  and (_25247_, _25246_, _25245_);
  or (_25248_, _25247_, _25243_);
  and (_25249_, _25248_, _03909_);
  nand (_25250_, _25235_, _03908_);
  nor (_25251_, _25250_, _25201_);
  or (_25252_, _25251_, _04027_);
  or (_25255_, _25252_, _25249_);
  and (_25256_, _25255_, _25190_);
  or (_25257_, _25256_, _03914_);
  nor (_25258_, _12177_, _10000_);
  or (_25259_, _25187_, _06567_);
  or (_25260_, _25259_, _25258_);
  and (_25261_, _25260_, _06572_);
  and (_25262_, _25261_, _25257_);
  and (_25263_, _25245_, _04011_);
  or (_25264_, _25263_, _17157_);
  or (_25266_, _25264_, _25262_);
  or (_25267_, _25202_, _04144_);
  and (_25268_, _25267_, _43152_);
  and (_25269_, _25268_, _25266_);
  or (_25270_, _25269_, _25185_);
  and (_43498_, _25270_, _41894_);
  not (_25271_, \oc8051_golden_model_1.DPH [1]);
  nor (_25272_, _43152_, _25271_);
  nand (_25273_, _05509_, _04595_);
  or (_25274_, _05509_, \oc8051_golden_model_1.DPH [1]);
  and (_25276_, _25274_, _03903_);
  and (_25277_, _25276_, _25273_);
  nor (_25278_, _09977_, \oc8051_golden_model_1.DPH [1]);
  nor (_25279_, _25278_, _09978_);
  and (_25280_, _25279_, _09878_);
  and (_25281_, _12262_, _05509_);
  not (_25282_, _25281_);
  and (_25283_, _25282_, _25274_);
  or (_25284_, _25283_, _04722_);
  nor (_25285_, _05509_, _25271_);
  and (_25287_, _05509_, \oc8051_golden_model_1.ACC [1]);
  or (_25288_, _25287_, _25285_);
  and (_25289_, _25288_, _04707_);
  nor (_25290_, _04707_, _25271_);
  or (_25291_, _25290_, _03850_);
  or (_25292_, _25291_, _25289_);
  and (_25293_, _25292_, _04733_);
  and (_25294_, _25293_, _25284_);
  and (_25295_, _05509_, _04900_);
  or (_25296_, _25295_, _25285_);
  and (_25298_, _25296_, _03848_);
  or (_25299_, _25298_, _03854_);
  or (_25300_, _25299_, _25294_);
  or (_25301_, _25288_, _03855_);
  and (_25302_, _25301_, _09879_);
  and (_25303_, _25302_, _25300_);
  or (_25304_, _25303_, _25280_);
  and (_25305_, _25304_, _09861_);
  nor (_25306_, _04563_, _09861_);
  or (_25307_, _25306_, _07927_);
  or (_25309_, _25307_, _25305_);
  and (_25310_, _06961_, _05509_);
  or (_25311_, _25285_, _03738_);
  or (_25312_, _25311_, _25310_);
  or (_25313_, _25296_, _07925_);
  and (_25314_, _25313_, _03820_);
  and (_25315_, _25314_, _25312_);
  and (_25316_, _25315_, _25309_);
  nor (_25317_, _12352_, _10000_);
  or (_25318_, _25317_, _25285_);
  and (_25320_, _25318_, _03455_);
  or (_25321_, _25320_, _25316_);
  and (_25322_, _25321_, _04778_);
  or (_25323_, _25322_, _25277_);
  and (_25324_, _25323_, _04790_);
  or (_25325_, _12366_, _10000_);
  and (_25326_, _25274_, _03897_);
  and (_25327_, _25326_, _25325_);
  or (_25328_, _25327_, _04018_);
  or (_25329_, _25328_, _25324_);
  and (_25331_, _08752_, _05509_);
  or (_25332_, _25331_, _25285_);
  or (_25333_, _25332_, _04792_);
  and (_25334_, _25333_, _03909_);
  and (_25335_, _25334_, _25329_);
  or (_25336_, _12244_, _10000_);
  and (_25337_, _25274_, _03908_);
  and (_25338_, _25337_, _25336_);
  or (_25339_, _25338_, _04027_);
  or (_25340_, _25339_, _25335_);
  and (_25342_, _08750_, _05509_);
  or (_25343_, _25285_, _04785_);
  or (_25344_, _25343_, _25342_);
  and (_25345_, _25344_, _06567_);
  and (_25346_, _25345_, _25340_);
  or (_25347_, _25273_, _08366_);
  and (_25348_, _25274_, _03914_);
  and (_25349_, _25348_, _25347_);
  or (_25350_, _25349_, _04011_);
  or (_25351_, _25350_, _25346_);
  nor (_25353_, _08751_, _10000_);
  or (_25354_, _25353_, _25285_);
  or (_25355_, _25354_, _06572_);
  and (_25356_, _25355_, _03774_);
  and (_25357_, _25356_, _25351_);
  and (_25358_, _25283_, _03773_);
  or (_25359_, _25358_, _03772_);
  or (_25360_, _25359_, _25357_);
  or (_25361_, _25285_, _04060_);
  or (_25362_, _25361_, _25281_);
  and (_25364_, _25362_, _43152_);
  and (_25365_, _25364_, _25360_);
  or (_25366_, _25365_, _25272_);
  and (_43499_, _25366_, _41894_);
  or (_25367_, _43152_, \oc8051_golden_model_1.DPH [2]);
  and (_25368_, _25367_, _41894_);
  and (_25369_, _10000_, \oc8051_golden_model_1.DPH [2]);
  and (_25370_, _05509_, _06495_);
  or (_25371_, _25370_, _25369_);
  or (_25372_, _25371_, _04778_);
  or (_25374_, _09978_, \oc8051_golden_model_1.DPH [2]);
  nor (_25375_, _09979_, _09879_);
  and (_25376_, _25375_, _25374_);
  nor (_25377_, _12471_, _10000_);
  or (_25378_, _25377_, _25369_);
  or (_25379_, _25378_, _04722_);
  and (_25380_, _05509_, \oc8051_golden_model_1.ACC [2]);
  or (_25381_, _25380_, _25369_);
  and (_25382_, _25381_, _04707_);
  and (_25383_, _04708_, \oc8051_golden_model_1.DPH [2]);
  or (_25385_, _25383_, _03850_);
  or (_25386_, _25385_, _25382_);
  and (_25387_, _25386_, _04733_);
  and (_25388_, _25387_, _25379_);
  and (_25389_, _05509_, _05307_);
  or (_25390_, _25389_, _25369_);
  and (_25391_, _25390_, _03848_);
  or (_25392_, _25391_, _03854_);
  or (_25393_, _25392_, _25388_);
  or (_25394_, _25381_, _03855_);
  and (_25396_, _25394_, _09879_);
  and (_25397_, _25396_, _25393_);
  or (_25398_, _25397_, _25376_);
  and (_25399_, _25398_, _09861_);
  nor (_25400_, _04139_, _09861_);
  or (_25401_, _25400_, _07927_);
  or (_25402_, _25401_, _25399_);
  and (_25403_, _06965_, _05509_);
  or (_25404_, _25369_, _03738_);
  or (_25405_, _25404_, _25403_);
  or (_25407_, _25390_, _07925_);
  and (_25408_, _25407_, _03820_);
  and (_25409_, _25408_, _25405_);
  and (_25410_, _25409_, _25402_);
  nor (_25411_, _12572_, _10000_);
  or (_25412_, _25411_, _25369_);
  and (_25413_, _25412_, _03455_);
  or (_25414_, _25413_, _03903_);
  or (_25415_, _25414_, _25410_);
  and (_25416_, _25415_, _25372_);
  or (_25417_, _25416_, _03897_);
  and (_25418_, _12586_, _05509_);
  or (_25419_, _25369_, _04790_);
  or (_25420_, _25419_, _25418_);
  and (_25421_, _25420_, _04792_);
  and (_25422_, _25421_, _25417_);
  and (_25423_, _08748_, _05509_);
  or (_25424_, _25423_, _25369_);
  and (_25425_, _25424_, _04018_);
  or (_25426_, _25425_, _25422_);
  and (_25429_, _25426_, _03909_);
  or (_25430_, _25369_, _05765_);
  and (_25431_, _25371_, _03908_);
  and (_25432_, _25431_, _25430_);
  or (_25433_, _25432_, _25429_);
  and (_25434_, _25433_, _04785_);
  and (_25435_, _25381_, _04027_);
  and (_25436_, _25435_, _25430_);
  or (_25437_, _25436_, _03914_);
  or (_25438_, _25437_, _25434_);
  nor (_25440_, _12585_, _10000_);
  or (_25441_, _25369_, _06567_);
  or (_25442_, _25441_, _25440_);
  and (_25443_, _25442_, _06572_);
  and (_25444_, _25443_, _25438_);
  nor (_25445_, _08747_, _10000_);
  or (_25446_, _25445_, _25369_);
  and (_25447_, _25446_, _04011_);
  or (_25448_, _25447_, _03773_);
  or (_25449_, _25448_, _25444_);
  or (_25451_, _25378_, _03774_);
  and (_25452_, _25451_, _04060_);
  and (_25453_, _25452_, _25449_);
  and (_25454_, _12642_, _05509_);
  or (_25455_, _25454_, _25369_);
  and (_25456_, _25455_, _03772_);
  or (_25457_, _25456_, _43156_);
  or (_25458_, _25457_, _25453_);
  and (_43500_, _25458_, _25368_);
  or (_25459_, _43152_, \oc8051_golden_model_1.DPH [3]);
  and (_25461_, _25459_, _41894_);
  not (_25462_, \oc8051_golden_model_1.DPH [3]);
  nor (_25463_, _05509_, _25462_);
  and (_25464_, _05509_, _06345_);
  or (_25465_, _25464_, _25463_);
  or (_25466_, _25465_, _04778_);
  nor (_25467_, _12681_, _10000_);
  or (_25468_, _25467_, _25463_);
  or (_25469_, _25468_, _04722_);
  and (_25470_, _05509_, \oc8051_golden_model_1.ACC [3]);
  or (_25472_, _25470_, _25463_);
  and (_25473_, _25472_, _04707_);
  nor (_25474_, _04707_, _25462_);
  or (_25475_, _25474_, _03850_);
  or (_25476_, _25475_, _25473_);
  and (_25477_, _25476_, _04733_);
  and (_25478_, _25477_, _25469_);
  and (_25479_, _05509_, _05119_);
  or (_25480_, _25479_, _25463_);
  and (_25481_, _25480_, _03848_);
  or (_25483_, _25481_, _03854_);
  or (_25484_, _25483_, _25478_);
  or (_25485_, _25472_, _03855_);
  and (_25486_, _25485_, _09879_);
  and (_25487_, _25486_, _25484_);
  or (_25488_, _09979_, \oc8051_golden_model_1.DPH [3]);
  nor (_25489_, _09980_, _09879_);
  and (_25490_, _25489_, _25488_);
  or (_25491_, _25490_, _25487_);
  and (_25492_, _25491_, _09861_);
  nor (_25494_, _09861_, _03678_);
  or (_25495_, _25494_, _07927_);
  or (_25496_, _25495_, _25492_);
  and (_25497_, _06964_, _05509_);
  or (_25498_, _25463_, _03738_);
  or (_25499_, _25498_, _25497_);
  or (_25500_, _25480_, _07925_);
  and (_25501_, _25500_, _03820_);
  and (_25502_, _25501_, _25499_);
  and (_25503_, _25502_, _25496_);
  nor (_25505_, _12775_, _10000_);
  or (_25506_, _25505_, _25463_);
  and (_25507_, _25506_, _03455_);
  or (_25508_, _25507_, _03903_);
  or (_25509_, _25508_, _25503_);
  and (_25510_, _25509_, _25466_);
  or (_25511_, _25510_, _03897_);
  and (_25512_, _12789_, _05509_);
  or (_25513_, _25512_, _25463_);
  or (_25514_, _25513_, _04790_);
  and (_25516_, _25514_, _04792_);
  and (_25517_, _25516_, _25511_);
  and (_25518_, _10491_, _05509_);
  or (_25519_, _25518_, _25463_);
  and (_25520_, _25519_, _04018_);
  or (_25521_, _25520_, _25517_);
  and (_25522_, _25521_, _03909_);
  or (_25523_, _25463_, _05622_);
  and (_25524_, _25465_, _03908_);
  and (_25525_, _25524_, _25523_);
  or (_25527_, _25525_, _25522_);
  and (_25528_, _25527_, _04785_);
  and (_25529_, _25472_, _04027_);
  and (_25530_, _25529_, _25523_);
  or (_25531_, _25530_, _03914_);
  or (_25532_, _25531_, _25528_);
  nor (_25533_, _12788_, _10000_);
  or (_25534_, _25463_, _06567_);
  or (_25535_, _25534_, _25533_);
  and (_25536_, _25535_, _06572_);
  and (_25538_, _25536_, _25532_);
  nor (_25539_, _08742_, _10000_);
  or (_25540_, _25539_, _25463_);
  and (_25541_, _25540_, _04011_);
  or (_25542_, _25541_, _03773_);
  or (_25543_, _25542_, _25538_);
  or (_25544_, _25468_, _03774_);
  and (_25545_, _25544_, _04060_);
  and (_25546_, _25545_, _25543_);
  and (_25547_, _12848_, _05509_);
  or (_25549_, _25547_, _25463_);
  and (_25550_, _25549_, _03772_);
  or (_25551_, _25550_, _43156_);
  or (_25552_, _25551_, _25546_);
  and (_43503_, _25552_, _25461_);
  or (_25553_, _43152_, \oc8051_golden_model_1.DPH [4]);
  and (_25554_, _25553_, _41894_);
  not (_25555_, \oc8051_golden_model_1.DPH [4]);
  nor (_25556_, _05509_, _25555_);
  and (_25557_, _06456_, _05509_);
  or (_25559_, _25557_, _25556_);
  or (_25560_, _25559_, _04778_);
  nor (_25561_, _12891_, _10000_);
  or (_25562_, _25561_, _25556_);
  or (_25563_, _25562_, _04722_);
  and (_25564_, _05509_, \oc8051_golden_model_1.ACC [4]);
  or (_25565_, _25564_, _25556_);
  and (_25566_, _25565_, _04707_);
  nor (_25567_, _04707_, _25555_);
  or (_25568_, _25567_, _03850_);
  or (_25570_, _25568_, _25566_);
  and (_25571_, _25570_, _04733_);
  and (_25572_, _25571_, _25563_);
  and (_25573_, _05950_, _05509_);
  or (_25574_, _25573_, _25556_);
  and (_25575_, _25574_, _03848_);
  or (_25576_, _25575_, _03854_);
  or (_25577_, _25576_, _25572_);
  or (_25578_, _25565_, _03855_);
  and (_25579_, _25578_, _09879_);
  and (_25581_, _25579_, _25577_);
  or (_25582_, _09980_, \oc8051_golden_model_1.DPH [4]);
  nor (_25583_, _09981_, _09879_);
  and (_25584_, _25583_, _25582_);
  or (_25585_, _25584_, _25581_);
  and (_25586_, _25585_, _09861_);
  nor (_25587_, _04526_, _09861_);
  or (_25588_, _25587_, _07927_);
  or (_25589_, _25588_, _25586_);
  and (_25590_, _06969_, _05509_);
  or (_25592_, _25556_, _03738_);
  or (_25593_, _25592_, _25590_);
  or (_25594_, _25574_, _07925_);
  and (_25595_, _25594_, _03820_);
  and (_25596_, _25595_, _25593_);
  and (_25597_, _25596_, _25589_);
  nor (_25598_, _12982_, _10000_);
  or (_25599_, _25598_, _25556_);
  and (_25600_, _25599_, _03455_);
  or (_25601_, _25600_, _03903_);
  or (_25603_, _25601_, _25597_);
  and (_25604_, _25603_, _25560_);
  or (_25605_, _25604_, _03897_);
  and (_25606_, _12997_, _05509_);
  or (_25607_, _25606_, _25556_);
  or (_25608_, _25607_, _04790_);
  and (_25609_, _25608_, _04792_);
  and (_25610_, _25609_, _25605_);
  and (_25611_, _08741_, _05509_);
  or (_25612_, _25611_, _25556_);
  and (_25613_, _25612_, _04018_);
  or (_25614_, _25613_, _25610_);
  and (_25615_, _25614_, _03909_);
  or (_25616_, _25556_, _08336_);
  and (_25617_, _25559_, _03908_);
  and (_25618_, _25617_, _25616_);
  or (_25619_, _25618_, _25615_);
  and (_25620_, _25619_, _04785_);
  and (_25621_, _25565_, _04027_);
  and (_25622_, _25621_, _25616_);
  or (_25625_, _25622_, _03914_);
  or (_25626_, _25625_, _25620_);
  nor (_25627_, _12996_, _10000_);
  or (_25628_, _25556_, _06567_);
  or (_25629_, _25628_, _25627_);
  and (_25630_, _25629_, _06572_);
  and (_25631_, _25630_, _25626_);
  nor (_25632_, _08740_, _10000_);
  or (_25633_, _25632_, _25556_);
  and (_25634_, _25633_, _04011_);
  or (_25636_, _25634_, _03773_);
  or (_25637_, _25636_, _25631_);
  or (_25638_, _25562_, _03774_);
  and (_25639_, _25638_, _04060_);
  and (_25640_, _25639_, _25637_);
  and (_25641_, _13056_, _05509_);
  or (_25642_, _25641_, _25556_);
  and (_25643_, _25642_, _03772_);
  or (_25644_, _25643_, _43156_);
  or (_25645_, _25644_, _25640_);
  and (_43504_, _25645_, _25554_);
  not (_25647_, \oc8051_golden_model_1.DPH [5]);
  nor (_25648_, _43152_, _25647_);
  nor (_25649_, _05509_, _25647_);
  and (_25650_, _06447_, _05509_);
  or (_25651_, _25650_, _25649_);
  or (_25652_, _25651_, _04778_);
  nor (_25653_, _13090_, _10000_);
  or (_25654_, _25653_, _25649_);
  or (_25655_, _25654_, _04722_);
  and (_25657_, _05509_, \oc8051_golden_model_1.ACC [5]);
  or (_25658_, _25657_, _25649_);
  and (_25659_, _25658_, _04707_);
  nor (_25660_, _04707_, _25647_);
  or (_25661_, _25660_, _03850_);
  or (_25662_, _25661_, _25659_);
  and (_25663_, _25662_, _04733_);
  and (_25664_, _25663_, _25655_);
  and (_25665_, _05857_, _05509_);
  or (_25666_, _25665_, _25649_);
  and (_25668_, _25666_, _03848_);
  or (_25669_, _25668_, _03854_);
  or (_25670_, _25669_, _25664_);
  or (_25671_, _25658_, _03855_);
  and (_25672_, _25671_, _09879_);
  and (_25673_, _25672_, _25670_);
  or (_25674_, _09981_, \oc8051_golden_model_1.DPH [5]);
  and (_25675_, _09982_, _09878_);
  and (_25676_, _25675_, _25674_);
  or (_25677_, _25676_, _25673_);
  and (_25679_, _25677_, _09861_);
  nor (_25680_, _04093_, _09861_);
  or (_25681_, _25680_, _07927_);
  or (_25682_, _25681_, _25679_);
  and (_25683_, _06968_, _05509_);
  or (_25684_, _25649_, _03738_);
  or (_25685_, _25684_, _25683_);
  or (_25686_, _25666_, _07925_);
  and (_25687_, _25686_, _03820_);
  and (_25688_, _25687_, _25685_);
  and (_25690_, _25688_, _25682_);
  nor (_25691_, _13182_, _10000_);
  or (_25692_, _25691_, _25649_);
  and (_25693_, _25692_, _03455_);
  or (_25694_, _25693_, _03903_);
  or (_25695_, _25694_, _25690_);
  and (_25696_, _25695_, _25652_);
  or (_25697_, _25696_, _03897_);
  and (_25698_, _13196_, _05509_);
  or (_25699_, _25698_, _25649_);
  or (_25701_, _25699_, _04790_);
  and (_25702_, _25701_, _04792_);
  and (_25703_, _25702_, _25697_);
  and (_25704_, _10493_, _05509_);
  or (_25705_, _25704_, _25649_);
  and (_25706_, _25705_, _04018_);
  or (_25707_, _25706_, _25703_);
  and (_25708_, _25707_, _03909_);
  or (_25709_, _25649_, _08335_);
  and (_25710_, _25651_, _03908_);
  and (_25712_, _25710_, _25709_);
  or (_25713_, _25712_, _25708_);
  and (_25714_, _25713_, _04785_);
  and (_25715_, _25658_, _04027_);
  and (_25716_, _25715_, _25709_);
  or (_25717_, _25716_, _03914_);
  or (_25718_, _25717_, _25714_);
  nor (_25719_, _13195_, _10000_);
  or (_25720_, _25649_, _06567_);
  or (_25721_, _25720_, _25719_);
  and (_25723_, _25721_, _06572_);
  and (_25724_, _25723_, _25718_);
  nor (_25725_, _08738_, _10000_);
  or (_25726_, _25725_, _25649_);
  and (_25727_, _25726_, _04011_);
  or (_25728_, _25727_, _25724_);
  and (_25729_, _25728_, _03774_);
  and (_25730_, _25654_, _03773_);
  or (_25731_, _25730_, _03772_);
  or (_25732_, _25731_, _25729_);
  and (_25734_, _13255_, _05509_);
  or (_25735_, _25649_, _04060_);
  or (_25736_, _25735_, _25734_);
  and (_25737_, _25736_, _43152_);
  and (_25738_, _25737_, _25732_);
  or (_25739_, _25738_, _25648_);
  and (_43505_, _25739_, _41894_);
  or (_25740_, _43152_, \oc8051_golden_model_1.DPH [6]);
  and (_25741_, _25740_, _41894_);
  nor (_25742_, _05509_, _09976_);
  and (_25744_, _13394_, _05509_);
  or (_25745_, _25744_, _25742_);
  or (_25746_, _25745_, _04778_);
  nor (_25747_, _13293_, _10000_);
  or (_25748_, _25747_, _25742_);
  or (_25749_, _25748_, _04722_);
  and (_25750_, _05509_, \oc8051_golden_model_1.ACC [6]);
  or (_25751_, _25750_, _25742_);
  and (_25752_, _25751_, _04707_);
  nor (_25753_, _04707_, _09976_);
  or (_25755_, _25753_, _03850_);
  or (_25756_, _25755_, _25752_);
  and (_25757_, _25756_, _04733_);
  and (_25758_, _25757_, _25749_);
  and (_25759_, _06065_, _05509_);
  or (_25760_, _25759_, _25742_);
  and (_25761_, _25760_, _03848_);
  or (_25762_, _25761_, _03854_);
  or (_25763_, _25762_, _25758_);
  or (_25764_, _25751_, _03855_);
  and (_25766_, _25764_, _09879_);
  and (_25767_, _25766_, _25763_);
  nand (_25768_, _09982_, _09976_);
  nor (_25769_, _09983_, _09879_);
  and (_25770_, _25769_, _25768_);
  or (_25771_, _25770_, _25767_);
  and (_25772_, _25771_, _09861_);
  nor (_25773_, _09861_, _03810_);
  or (_25774_, _25773_, _07927_);
  or (_25775_, _25774_, _25772_);
  and (_25777_, _06641_, _05509_);
  or (_25778_, _25742_, _03738_);
  or (_25779_, _25778_, _25777_);
  or (_25780_, _25760_, _07925_);
  and (_25781_, _25780_, _03820_);
  and (_25782_, _25781_, _25779_);
  and (_25783_, _25782_, _25775_);
  nor (_25784_, _13387_, _10000_);
  or (_25785_, _25784_, _25742_);
  and (_25786_, _25785_, _03455_);
  or (_25788_, _25786_, _03903_);
  or (_25789_, _25788_, _25783_);
  and (_25790_, _25789_, _25746_);
  or (_25791_, _25790_, _03897_);
  and (_25792_, _13402_, _05509_);
  or (_25793_, _25742_, _04790_);
  or (_25794_, _25793_, _25792_);
  and (_25795_, _25794_, _04792_);
  and (_25796_, _25795_, _25791_);
  and (_25797_, _08736_, _05509_);
  or (_25799_, _25797_, _25742_);
  and (_25800_, _25799_, _04018_);
  or (_25801_, _25800_, _25796_);
  and (_25802_, _25801_, _03909_);
  or (_25803_, _25742_, _08322_);
  and (_25804_, _25745_, _03908_);
  and (_25805_, _25804_, _25803_);
  or (_25806_, _25805_, _25802_);
  and (_25807_, _25806_, _04785_);
  and (_25808_, _25751_, _04027_);
  and (_25810_, _25808_, _25803_);
  or (_25811_, _25810_, _03914_);
  or (_25812_, _25811_, _25807_);
  nor (_25813_, _13401_, _10000_);
  or (_25814_, _25742_, _06567_);
  or (_25815_, _25814_, _25813_);
  and (_25816_, _25815_, _06572_);
  and (_25817_, _25816_, _25812_);
  nor (_25818_, _08735_, _10000_);
  or (_25819_, _25818_, _25742_);
  and (_25821_, _25819_, _04011_);
  or (_25822_, _25821_, _03773_);
  or (_25823_, _25822_, _25817_);
  or (_25824_, _25748_, _03774_);
  and (_25825_, _25824_, _04060_);
  and (_25826_, _25825_, _25823_);
  nor (_25827_, _13460_, _10000_);
  or (_25828_, _25827_, _25742_);
  and (_25829_, _25828_, _03772_);
  or (_25830_, _25829_, _43156_);
  or (_25832_, _25830_, _25826_);
  and (_43506_, _25832_, _25741_);
  nor (_25833_, _03901_, _03413_);
  not (_25834_, _25833_);
  and (_25835_, _25834_, _04382_);
  and (_25836_, _10906_, \oc8051_golden_model_1.PC [0]);
  and (_25837_, _04382_, \oc8051_golden_model_1.PC [0]);
  nor (_25838_, _25837_, _10163_);
  nor (_25839_, _25838_, _10906_);
  nor (_25840_, _25839_, _25836_);
  and (_25842_, _25840_, _03374_);
  and (_25843_, _10936_, _10943_);
  nor (_25844_, _25843_, _03119_);
  and (_25845_, _10059_, _08773_);
  nor (_25846_, _25845_, _03119_);
  not (_25847_, _03388_);
  and (_25848_, _10654_, _03909_);
  nor (_25849_, _25848_, _03119_);
  not (_25850_, _03405_);
  and (_25851_, _10082_, _04790_);
  nor (_25853_, _25851_, _03119_);
  and (_25854_, _03903_, _03119_);
  nor (_25855_, _03921_, _03455_);
  and (_25856_, _25855_, _10556_);
  nor (_25857_, _25856_, _03119_);
  nor (_25858_, _04382_, _03428_);
  and (_25859_, _10249_, _03119_);
  not (_25860_, _25838_);
  nor (_25861_, _25860_, _10249_);
  or (_25862_, _25861_, _10444_);
  or (_25864_, _25862_, _25859_);
  and (_25865_, _10476_, _03119_);
  nor (_25866_, _25860_, _10476_);
  or (_25867_, _25866_, _25865_);
  or (_25868_, _25867_, _10441_);
  nand (_25869_, _04382_, _03768_);
  nor (_25870_, _05011_, _04263_);
  or (_25871_, _25870_, _03119_);
  nand (_25872_, _25870_, _03119_);
  and (_25873_, _25872_, _25871_);
  nand (_25875_, _10402_, _03770_);
  or (_25876_, _25875_, _25873_);
  or (_25877_, _10402_, _03119_);
  and (_25878_, _25877_, _04266_);
  and (_25879_, _25878_, _25876_);
  and (_25880_, _25879_, _25869_);
  and (_25881_, _03715_, _03119_);
  nor (_25882_, _25881_, _10324_);
  and (_25883_, _25882_, _10383_);
  and (_25884_, _06126_, _10380_);
  and (_25886_, _06951_, _06124_);
  and (_25887_, _25886_, _25884_);
  and (_25888_, _25887_, \oc8051_golden_model_1.PC [0]);
  or (_25889_, _25888_, _25883_);
  and (_25890_, _25889_, _04267_);
  or (_25891_, _25890_, _25880_);
  and (_25892_, _25891_, _04717_);
  and (_25893_, _04716_, _03119_);
  or (_25894_, _25893_, _25892_);
  and (_25895_, _25894_, _04722_);
  and (_25897_, _06152_, _05621_);
  and (_25898_, _05764_, _05669_);
  and (_25899_, _25898_, _10262_);
  and (_25900_, _25899_, _06070_);
  and (_25901_, _25900_, _25897_);
  nor (_25902_, _25860_, _25901_);
  and (_25903_, _10262_, _05669_);
  and (_25904_, _06154_, _25903_);
  and (_25905_, _06152_, _06070_);
  and (_25906_, _25905_, _25904_);
  and (_25908_, _25906_, _03119_);
  or (_25909_, _25908_, _25902_);
  and (_25910_, _25909_, _03850_);
  or (_25911_, _25910_, _10413_);
  or (_25912_, _25911_, _25895_);
  or (_25913_, _10412_, _03119_);
  and (_25914_, _25913_, _03431_);
  and (_25915_, _25914_, _25912_);
  or (_25916_, _04382_, _03431_);
  and (_25917_, _10431_, _10421_);
  nand (_25919_, _25917_, _25916_);
  or (_25920_, _25919_, _25915_);
  or (_25921_, _25917_, _03119_);
  and (_25922_, _25921_, _03434_);
  and (_25923_, _25922_, _25920_);
  nor (_25924_, _04382_, _03434_);
  or (_25925_, _25924_, _10442_);
  or (_25926_, _25925_, _25923_);
  and (_25927_, _25926_, _25868_);
  or (_25928_, _25927_, _03925_);
  and (_25930_, _25928_, _03918_);
  and (_25931_, _25930_, _25864_);
  nor (_25932_, _25860_, _10498_);
  and (_25933_, _10498_, _03119_);
  or (_25934_, _25933_, _25932_);
  and (_25935_, _25934_, _03868_);
  or (_25936_, _25935_, _25931_);
  and (_25937_, _25936_, _10486_);
  and (_25938_, _10515_, \oc8051_golden_model_1.PC [0]);
  and (_25939_, _10485_, _03119_);
  nor (_25941_, _25838_, _10515_);
  nor (_25942_, _25941_, _11857_);
  nor (_25943_, _25942_, _25939_);
  nor (_25944_, _25943_, _25938_);
  nor (_25945_, _25944_, _25937_);
  nor (_25946_, _25945_, _05049_);
  or (_25947_, _25946_, _10093_);
  nor (_25948_, _25947_, _25858_);
  not (_25949_, _03441_);
  nor (_25950_, _10092_, _03119_);
  nor (_25952_, _25950_, _25949_);
  not (_25953_, _25952_);
  nor (_25954_, _25953_, _25948_);
  nor (_25955_, _04382_, _03441_);
  and (_25956_, _10087_, _03426_);
  not (_25957_, _25956_);
  nor (_25958_, _25957_, _25955_);
  not (_25959_, _25958_);
  nor (_25960_, _25959_, _25954_);
  nor (_25961_, _25956_, _03119_);
  nor (_25962_, _25961_, _03456_);
  not (_25963_, _25962_);
  nor (_25964_, _25963_, _25960_);
  nor (_25965_, _04382_, _06141_);
  not (_25966_, _25856_);
  nor (_25967_, _25966_, _25965_);
  not (_25968_, _25967_);
  nor (_25969_, _25968_, _25964_);
  or (_25970_, _25969_, _03398_);
  nor (_25971_, _25970_, _25857_);
  nor (_25974_, _10564_, _03398_);
  not (_25975_, _25974_);
  nand (_25976_, _10565_, _04382_);
  and (_25977_, _25976_, _25975_);
  nor (_25978_, _25977_, _25971_);
  nor (_25979_, _25882_, _10565_);
  nor (_25980_, _25979_, _25978_);
  and (_25981_, _25980_, _04778_);
  or (_25982_, _25981_, _25854_);
  and (_25983_, _25982_, _10581_);
  and (_25985_, _10580_, _03491_);
  or (_25986_, _25985_, _25983_);
  and (_25987_, _25986_, _11641_);
  nor (_25988_, _04382_, _11641_);
  or (_25989_, _25988_, _25987_);
  and (_25990_, _25989_, _10621_);
  not (_25991_, _25851_);
  and (_25992_, _08826_, \oc8051_golden_model_1.PC [0]);
  and (_25993_, _25882_, _10627_);
  or (_25994_, _25993_, _25992_);
  and (_25996_, _25994_, _10620_);
  nor (_25997_, _25996_, _25991_);
  not (_25998_, _25997_);
  nor (_25999_, _25998_, _25990_);
  nor (_26000_, _25999_, _25853_);
  and (_26001_, _26000_, _25850_);
  nor (_26002_, _04382_, _25850_);
  or (_26003_, _26002_, _26001_);
  and (_26004_, _26003_, _10644_);
  not (_26005_, _25848_);
  nor (_26007_, _25882_, _10627_);
  nor (_26008_, _08826_, \oc8051_golden_model_1.PC [0]);
  nor (_26009_, _26008_, _10644_);
  not (_26010_, _26009_);
  nor (_26011_, _26010_, _26007_);
  nor (_26012_, _26011_, _26005_);
  not (_26013_, _26012_);
  nor (_26014_, _26013_, _26004_);
  nor (_26015_, _26014_, _25849_);
  and (_26016_, _26015_, _25847_);
  nor (_26018_, _04382_, _25847_);
  or (_26019_, _26018_, _26016_);
  and (_26020_, _26019_, _10075_);
  and (_26021_, _10072_, _06567_);
  not (_26022_, _26021_);
  nor (_26023_, _25882_, \oc8051_golden_model_1.PSW [7]);
  and (_26024_, \oc8051_golden_model_1.PSW [7], _03119_);
  nor (_26025_, _26024_, _10075_);
  not (_26026_, _26025_);
  nor (_26027_, _26026_, _26023_);
  nor (_26029_, _26027_, _26022_);
  not (_26030_, _26029_);
  nor (_26031_, _26030_, _26020_);
  nor (_26032_, _10063_, _03393_);
  not (_26033_, _26032_);
  nor (_26034_, _26021_, _03119_);
  or (_26035_, _26034_, _26033_);
  or (_26036_, _26035_, _26031_);
  nor (_26037_, _08435_, _03119_);
  and (_26038_, _08435_, _03119_);
  nor (_26040_, _26038_, _26037_);
  nor (_26041_, _26040_, _10064_);
  not (_26042_, _03393_);
  nor (_26043_, _04382_, _26042_);
  and (_26044_, _10061_, _08658_);
  not (_26045_, _26044_);
  or (_26046_, _26045_, _26043_);
  nor (_26047_, _26046_, _26041_);
  and (_26048_, _26047_, _26036_);
  nor (_26049_, _26044_, _03119_);
  nor (_26051_, _26049_, _04034_);
  not (_26052_, _26051_);
  nor (_26053_, _26052_, _26048_);
  and (_26054_, _06962_, _04034_);
  or (_26055_, _26054_, _26053_);
  and (_26056_, _26055_, _03384_);
  nor (_26057_, _04382_, _03384_);
  or (_26058_, _26057_, _26056_);
  and (_26059_, _26058_, _04097_);
  and (_26060_, _25860_, _10906_);
  nor (_26062_, _10906_, _03119_);
  or (_26063_, _26062_, _04097_);
  or (_26064_, _26063_, _26060_);
  and (_26065_, _26064_, _25845_);
  not (_26066_, _26065_);
  nor (_26067_, _26066_, _26059_);
  nor (_26068_, _26067_, _25846_);
  and (_26069_, _26068_, _03778_);
  and (_26070_, _06962_, _03777_);
  or (_26071_, _26070_, _26069_);
  and (_26072_, _26071_, _03411_);
  nor (_26073_, _04382_, _03411_);
  nor (_26074_, _26073_, _26072_);
  nor (_26075_, _26074_, _03775_);
  not (_26076_, _25843_);
  and (_26077_, _25840_, _03775_);
  nor (_26078_, _26077_, _26076_);
  not (_26079_, _26078_);
  nor (_26080_, _26079_, _26075_);
  nor (_26081_, _26080_, _25844_);
  nor (_26084_, _26081_, _05223_);
  and (_26085_, _05223_, _04382_);
  nor (_26086_, _26085_, _03374_);
  not (_26087_, _26086_);
  nor (_26088_, _26087_, _26084_);
  nor (_26089_, _26088_, _25842_);
  and (_26090_, _10958_, _10965_);
  not (_26091_, _26090_);
  or (_26092_, _26091_, _26089_);
  or (_26093_, _26090_, \oc8051_golden_model_1.PC [0]);
  and (_26095_, _26093_, _25833_);
  and (_26096_, _26095_, _26092_);
  or (_26097_, _26096_, _10042_);
  nor (_26098_, _26097_, _25835_);
  and (_26099_, _10042_, _03119_);
  nor (_26100_, _26099_, _26098_);
  nand (_26101_, _26100_, _43152_);
  or (_26102_, _43152_, \oc8051_golden_model_1.PC [0]);
  and (_26103_, _26102_, _41894_);
  and (_43509_, _26103_, _26101_);
  and (_26105_, _10042_, _03948_);
  and (_26106_, _03772_, _03087_);
  and (_26107_, _10906_, _03447_);
  nor (_26108_, _10165_, _10163_);
  nor (_26109_, _26108_, _10166_);
  not (_26110_, _26109_);
  nor (_26111_, _26110_, _10906_);
  nor (_26112_, _26111_, _26107_);
  nor (_26113_, _26112_, _03375_);
  nor (_26114_, _26112_, _03776_);
  nor (_26116_, _10059_, _03948_);
  nor (_26117_, _10072_, _03948_);
  nor (_26118_, _10654_, _03948_);
  nor (_26119_, _08502_, _03948_);
  and (_26120_, _03746_, \oc8051_golden_model_1.PC [1]);
  and (_26121_, _04595_, _25949_);
  or (_26122_, _26121_, _03878_);
  and (_26123_, _10476_, _03447_);
  nor (_26124_, _26110_, _10476_);
  or (_26125_, _26124_, _26123_);
  nor (_26127_, _26125_, _10441_);
  nor (_26128_, _04595_, _03431_);
  or (_26129_, _10417_, _03948_);
  nor (_26130_, _10326_, _10324_);
  nor (_26131_, _26130_, _10327_);
  and (_26132_, _26131_, _10383_);
  and (_26133_, _10382_, _03087_);
  nor (_26134_, _26133_, _26132_);
  nor (_26135_, _26134_, _04266_);
  nand (_26136_, _04595_, _03768_);
  nor (_26138_, _05011_, _04230_);
  nor (_26139_, _04707_, \oc8051_golden_model_1.PC [0]);
  nor (_26140_, _26139_, _26138_);
  and (_26141_, _26140_, \oc8051_golden_model_1.PC [1]);
  nor (_26142_, _26140_, \oc8051_golden_model_1.PC [1]);
  nor (_26143_, _26142_, _26141_);
  or (_26144_, _26143_, _25875_);
  nor (_26145_, _10402_, _03948_);
  nor (_26146_, _26145_, _04267_);
  and (_26147_, _26146_, _26144_);
  and (_26149_, _26147_, _26136_);
  not (_26150_, _26149_);
  nor (_26151_, _04716_, _03850_);
  nand (_26152_, _26151_, _26150_);
  or (_26153_, _26152_, _26135_);
  nor (_26154_, _26110_, _25901_);
  and (_26155_, _25906_, _03447_);
  or (_26156_, _26155_, _04722_);
  or (_26157_, _26156_, _26154_);
  and (_26158_, _26157_, _26153_);
  or (_26160_, _26158_, _10413_);
  and (_26161_, _26160_, _26129_);
  and (_26162_, _26161_, _03764_);
  and (_26163_, _03763_, _03087_);
  or (_26164_, _26163_, _26162_);
  and (_26165_, _26164_, _03431_);
  nor (_26166_, _26165_, _26128_);
  nor (_26167_, _26166_, _03848_);
  not (_26168_, _10421_);
  and (_26169_, _03848_, _03087_);
  nor (_26171_, _26169_, _26168_);
  not (_26172_, _26171_);
  nor (_26173_, _26172_, _26167_);
  nor (_26174_, _10421_, _03948_);
  nor (_26175_, _26174_, _03854_);
  not (_26176_, _26175_);
  nor (_26177_, _26176_, _26173_);
  and (_26178_, _03854_, _03087_);
  nor (_26179_, _26178_, _10434_);
  not (_26180_, _26179_);
  nor (_26182_, _26180_, _26177_);
  nor (_26183_, _10431_, _03948_);
  nor (_26184_, _26183_, _03759_);
  not (_26185_, _26184_);
  nor (_26186_, _26185_, _26182_);
  and (_26187_, _03759_, _03087_);
  nor (_26188_, _26187_, _26186_);
  or (_26189_, _26188_, _10255_);
  or (_26190_, _04595_, _03434_);
  and (_26191_, _26190_, _26189_);
  or (_26193_, _26191_, _03758_);
  and (_26194_, _03758_, _03087_);
  nor (_26195_, _26194_, _10442_);
  and (_26196_, _26195_, _26193_);
  or (_26197_, _26196_, _26127_);
  nand (_26198_, _26197_, _10444_);
  and (_26199_, _10249_, _03447_);
  nor (_26200_, _26110_, _10249_);
  or (_26201_, _26200_, _10444_);
  nor (_26202_, _26201_, _26199_);
  nor (_26204_, _26202_, _03868_);
  nand (_26205_, _26204_, _26198_);
  and (_26206_, _10498_, _03948_);
  nor (_26207_, _26109_, _10498_);
  or (_26208_, _26207_, _03918_);
  or (_26209_, _26208_, _26206_);
  nand (_26210_, _26209_, _26205_);
  nand (_26211_, _26210_, _10486_);
  and (_26212_, _10515_, _03447_);
  nor (_26213_, _26110_, _10515_);
  nor (_26215_, _26213_, _26212_);
  nor (_26216_, _26215_, _11857_);
  and (_26217_, _10485_, _03948_);
  nor (_26218_, _26217_, _26216_);
  and (_26219_, _26218_, _03753_);
  nand (_26220_, _26219_, _26211_);
  and (_26221_, _03752_, \oc8051_golden_model_1.PC [1]);
  nor (_26222_, _26221_, _05049_);
  nand (_26223_, _26222_, _26220_);
  nor (_26224_, _04595_, _03428_);
  nor (_26226_, _04320_, _03843_);
  and (_26227_, _26226_, _03838_);
  nor (_26228_, _08166_, _03440_);
  not (_26229_, _26228_);
  and (_26230_, _26229_, _03830_);
  and (_26231_, _26230_, _26227_);
  not (_26232_, _26231_);
  nor (_26233_, _26232_, _26224_);
  nand (_26234_, _26233_, _26223_);
  nor (_26235_, _26231_, _03087_);
  nor (_26237_, _26235_, _10089_);
  nand (_26238_, _26237_, _26234_);
  and (_26239_, _10091_, _03447_);
  or (_26240_, _26239_, _10092_);
  nand (_26241_, _26240_, _26238_);
  nor (_26242_, _10091_, _03948_);
  nor (_26243_, _26242_, _03879_);
  nand (_26244_, _26243_, _26241_);
  and (_26245_, _03879_, _03087_);
  nor (_26246_, _26245_, _25949_);
  and (_26248_, _26246_, _26244_);
  or (_26249_, _26248_, _26122_);
  and (_26250_, _03878_, _03087_);
  nor (_26251_, _26250_, _15018_);
  and (_26252_, _26251_, _26249_);
  nor (_26253_, _10087_, _03948_);
  or (_26254_, _26253_, _26252_);
  nand (_26255_, _26254_, _10085_);
  nor (_26256_, _10085_, _03087_);
  nor (_26257_, _26256_, _03425_);
  nand (_26259_, _26257_, _26255_);
  and (_26260_, _03948_, _03425_);
  nor (_26261_, _26260_, _03746_);
  and (_26262_, _26261_, _26259_);
  or (_26263_, _26262_, _26120_);
  nand (_26264_, _26263_, _06141_);
  and (_26265_, _04595_, _03456_);
  nor (_26266_, _26265_, _03921_);
  nand (_26267_, _26266_, _26264_);
  and (_26268_, _03921_, _03447_);
  nor (_26270_, _26268_, _07927_);
  nand (_26271_, _26270_, _26267_);
  nor (_26272_, _07926_, _03087_);
  nor (_26273_, _26272_, _03455_);
  nand (_26274_, _26273_, _26271_);
  and (_26275_, _03455_, _03447_);
  nor (_26276_, _26275_, _10558_);
  nand (_26277_, _26276_, _26274_);
  nor (_26278_, _10556_, _03948_);
  nor (_26279_, _26278_, _03816_);
  nand (_26281_, _26279_, _26277_);
  nor (_26282_, _03398_, _03087_);
  or (_26283_, _26282_, _10560_);
  nand (_26284_, _26283_, _26281_);
  and (_26285_, _04595_, _03398_);
  nor (_26286_, _26285_, _10564_);
  nand (_26287_, _26286_, _26284_);
  and (_26288_, _26131_, _10564_);
  nor (_26289_, _26288_, _06309_);
  nand (_26290_, _26289_, _26287_);
  nor (_26292_, _06138_, _03087_);
  nor (_26293_, _26292_, _03903_);
  nand (_26294_, _26293_, _26290_);
  and (_26295_, _03903_, _03447_);
  nor (_26296_, _26295_, _08492_);
  and (_26297_, _26296_, _26294_);
  and (_26298_, _08492_, \oc8051_golden_model_1.PC [1]);
  or (_26299_, _26298_, _26297_);
  nand (_26300_, _26299_, _10581_);
  nor (_26301_, _10581_, _03465_);
  nor (_26303_, _26301_, _03815_);
  and (_26304_, _26303_, _26300_);
  and (_26305_, _03815_, _03087_);
  or (_26306_, _26305_, _03401_);
  or (_26307_, _26306_, _26304_);
  and (_26308_, _04595_, _03401_);
  nor (_26309_, _26308_, _10620_);
  nand (_26310_, _26309_, _26307_);
  nor (_26311_, _26131_, _08826_);
  and (_26312_, _08826_, \oc8051_golden_model_1.PC [1]);
  nor (_26314_, _26312_, _10621_);
  not (_26315_, _26314_);
  nor (_26316_, _26315_, _26311_);
  nor (_26317_, _26316_, _08503_);
  and (_26318_, _26317_, _26310_);
  or (_26319_, _26318_, _26119_);
  and (_26320_, _16845_, _08514_);
  nand (_26321_, _26320_, _26319_);
  nor (_26322_, _26320_, _03948_);
  nor (_26323_, _26322_, _04401_);
  nand (_26325_, _26323_, _26321_);
  and (_26326_, _04401_, _03948_);
  nor (_26327_, _26326_, _10080_);
  nand (_26328_, _26327_, _26325_);
  nor (_26329_, _10079_, _03087_);
  nor (_26330_, _26329_, _03897_);
  and (_26331_, _26330_, _26328_);
  and (_26332_, _03897_, _03447_);
  or (_26333_, _26332_, _04018_);
  nor (_26334_, _26333_, _26331_);
  and (_26336_, _04018_, \oc8051_golden_model_1.PC [1]);
  or (_26337_, _26336_, _26334_);
  nand (_26338_, _26337_, _25850_);
  and (_26339_, _04595_, _03405_);
  nor (_26340_, _26339_, _10643_);
  nand (_26341_, _26340_, _26338_);
  nor (_26342_, _26131_, _10627_);
  nor (_26343_, _08826_, _03087_);
  nor (_26344_, _26343_, _10644_);
  not (_26345_, _26344_);
  nor (_26347_, _26345_, _26342_);
  nor (_26348_, _26347_, _10656_);
  and (_26349_, _26348_, _26341_);
  or (_26350_, _26349_, _26118_);
  nand (_26351_, _26350_, _10658_);
  nor (_26352_, _10658_, _03087_);
  nor (_26353_, _26352_, _03908_);
  and (_26354_, _26353_, _26351_);
  and (_26355_, _03908_, _03447_);
  or (_26356_, _26355_, _04027_);
  nor (_26358_, _26356_, _26354_);
  and (_26359_, _04027_, \oc8051_golden_model_1.PC [1]);
  or (_26360_, _26359_, _26358_);
  nand (_26361_, _26360_, _25847_);
  and (_26362_, _04595_, _03388_);
  nor (_26363_, _26362_, _10074_);
  nand (_26364_, _26363_, _26361_);
  nor (_26365_, _26131_, \oc8051_golden_model_1.PSW [7]);
  and (_26366_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor (_26367_, _26366_, _10075_);
  not (_26369_, _26367_);
  nor (_26370_, _26369_, _26365_);
  nor (_26371_, _26370_, _10670_);
  and (_26372_, _26371_, _26364_);
  or (_26373_, _26372_, _26117_);
  nand (_26374_, _26373_, _08581_);
  nor (_26375_, _08581_, _03087_);
  nor (_26376_, _26375_, _03914_);
  and (_26377_, _26376_, _26374_);
  and (_26378_, _03914_, _03447_);
  or (_26380_, _26378_, _04011_);
  nor (_26381_, _26380_, _26377_);
  and (_26382_, _04011_, \oc8051_golden_model_1.PC [1]);
  nor (_26383_, _26382_, _26381_);
  nand (_26384_, _26383_, _26032_);
  nor (_26385_, _26131_, _08297_);
  and (_26386_, _08297_, \oc8051_golden_model_1.PC [1]);
  nor (_26387_, _26386_, _10064_);
  not (_26388_, _26387_);
  nor (_26389_, _26388_, _26385_);
  nor (_26391_, _04595_, _26042_);
  nor (_26392_, _26391_, _10688_);
  not (_26393_, _26392_);
  nor (_26394_, _26393_, _26389_);
  and (_26395_, _26394_, _26384_);
  nor (_26396_, _10061_, _03948_);
  or (_26397_, _26396_, _26395_);
  nand (_26398_, _26397_, _08628_);
  nor (_26399_, _08628_, _03087_);
  nor (_26400_, _26399_, _08657_);
  nand (_26402_, _26400_, _26398_);
  and (_26403_, _08657_, _03948_);
  nor (_26404_, _26403_, _04034_);
  and (_26405_, _26404_, _26402_);
  and (_26406_, _06688_, _04034_);
  or (_26407_, _26406_, _26405_);
  nand (_26408_, _26407_, _03384_);
  and (_26409_, _04595_, _03383_);
  nor (_26410_, _26409_, _03913_);
  nand (_26411_, _26410_, _26408_);
  and (_26413_, _26110_, _10906_);
  nor (_26414_, _10906_, _03447_);
  or (_26415_, _26414_, _04097_);
  nor (_26416_, _26415_, _26413_);
  nor (_26417_, _26416_, _10712_);
  and (_26418_, _26417_, _26411_);
  or (_26419_, _26418_, _26116_);
  nand (_26420_, _26419_, _10056_);
  nor (_26421_, _10056_, _03087_);
  nor (_26422_, _26421_, _08772_);
  and (_26424_, _26422_, _26420_);
  and (_26425_, _08772_, _03948_);
  or (_26426_, _26425_, _03777_);
  nor (_26427_, _26426_, _26424_);
  and (_26428_, _06688_, _03777_);
  or (_26429_, _26428_, _26427_);
  nand (_26430_, _26429_, _03411_);
  and (_26431_, _04595_, _03410_);
  nor (_26432_, _26431_, _03775_);
  and (_26433_, _26432_, _26430_);
  or (_26435_, _26433_, _26114_);
  nand (_26436_, _26435_, _04468_);
  and (_26437_, _05054_, _04813_);
  nor (_26438_, _04468_, _03447_);
  not (_26439_, _26438_);
  and (_26440_, _26439_, _26437_);
  nand (_26441_, _26440_, _26436_);
  nor (_26442_, _26437_, _03948_);
  nor (_26443_, _26442_, _03773_);
  nand (_26444_, _26443_, _26441_);
  not (_26446_, _10943_);
  and (_26447_, _03773_, _03087_);
  nor (_26448_, _26447_, _26446_);
  and (_26449_, _26448_, _26444_);
  nor (_26450_, _10943_, _03948_);
  or (_26451_, _26450_, _26449_);
  nand (_26452_, _26451_, _04819_);
  and (_26453_, _05223_, _04595_);
  nor (_26454_, _26453_, _03374_);
  and (_26455_, _26454_, _26452_);
  or (_26457_, _26455_, _26113_);
  nand (_26458_, _26457_, _12835_);
  not (_26459_, _05038_);
  and (_26460_, _12834_, _03948_);
  nor (_26461_, _26460_, _26459_);
  nand (_26462_, _26461_, _26458_);
  nor (_26463_, _05038_, _03948_);
  nor (_26464_, _26463_, _03772_);
  and (_26465_, _26464_, _26462_);
  or (_26466_, _26465_, _26106_);
  nand (_26468_, _26466_, _10965_);
  nor (_26469_, _10965_, _03447_);
  nor (_26470_, _26469_, _25834_);
  nand (_26471_, _26470_, _26468_);
  and (_26472_, _25834_, _04595_);
  nor (_26473_, _26472_, _10042_);
  and (_26474_, _26473_, _26471_);
  or (_26475_, _26474_, _26105_);
  or (_26476_, _26475_, _43156_);
  or (_26477_, _43152_, \oc8051_golden_model_1.PC [1]);
  and (_26479_, _26477_, _41894_);
  and (_43510_, _26479_, _26476_);
  and (_26480_, _10042_, _03518_);
  and (_26481_, _03772_, _03510_);
  and (_26482_, _03773_, _03510_);
  nor (_26483_, _10059_, _03518_);
  nor (_26484_, _10061_, _03518_);
  nor (_26485_, _10072_, _03518_);
  nor (_26486_, _10654_, _03518_);
  nor (_26487_, _10082_, _03518_);
  and (_26489_, _07919_, _08164_);
  nor (_26490_, _26489_, _03720_);
  and (_26491_, _10159_, _03921_);
  not (_26492_, _26491_);
  and (_26493_, _03746_, _03511_);
  nor (_26494_, _26231_, _03510_);
  and (_26495_, _10170_, _10167_);
  nor (_26496_, _26495_, _10171_);
  nor (_26497_, _26496_, _25901_);
  and (_26498_, _25901_, _10160_);
  nor (_26500_, _26498_, _26497_);
  or (_26501_, _26500_, _04722_);
  nor (_26502_, _10402_, _03518_);
  nand (_26503_, _04230_, _03511_);
  not (_26504_, _04263_);
  nor (_26505_, _05011_, _03092_);
  or (_26506_, _26505_, _04707_);
  and (_26507_, _26506_, _26504_);
  and (_26508_, _05011_, _03518_);
  or (_26509_, _26508_, _26507_);
  and (_26511_, _26509_, _26503_);
  and (_26512_, _04263_, _03518_);
  nor (_26513_, _26512_, _26511_);
  nor (_26514_, _26513_, _03768_);
  not (_26515_, _26514_);
  not (_26516_, _10402_);
  nor (_26517_, _04180_, _03770_);
  nor (_26518_, _26517_, _26516_);
  and (_26519_, _26518_, _26515_);
  nor (_26520_, _26519_, _26502_);
  nor (_26521_, _26520_, _04267_);
  and (_26522_, _10382_, _03510_);
  not (_26523_, _26522_);
  and (_26524_, _10331_, _10328_);
  nor (_26525_, _26524_, _10332_);
  and (_26526_, _26525_, _10383_);
  nor (_26527_, _26526_, _04266_);
  and (_26528_, _26527_, _26523_);
  or (_26529_, _26528_, _26521_);
  nor (_26530_, _26529_, _04716_);
  and (_26533_, _04716_, _03518_);
  or (_26534_, _26533_, _03850_);
  or (_26535_, _26534_, _26530_);
  and (_26536_, _26535_, _26501_);
  nor (_26537_, _26536_, _10413_);
  nor (_26538_, _10412_, _03518_);
  nor (_26539_, _26538_, _03763_);
  not (_26540_, _26539_);
  nor (_26541_, _26540_, _26537_);
  and (_26542_, _03763_, _03510_);
  or (_26544_, _26542_, _26541_);
  and (_26545_, _26544_, _03431_);
  nor (_26546_, _04180_, _03431_);
  or (_26547_, _26546_, _26545_);
  and (_26548_, _26547_, _04733_);
  and (_26549_, _03848_, _03510_);
  nor (_26550_, _26549_, _26168_);
  not (_26551_, _26550_);
  nor (_26552_, _26551_, _26548_);
  nor (_26553_, _10421_, _03518_);
  nor (_26555_, _26553_, _03854_);
  not (_26556_, _26555_);
  nor (_26557_, _26556_, _26552_);
  and (_26558_, _03854_, _03510_);
  nor (_26559_, _26558_, _10434_);
  not (_26560_, _26559_);
  or (_26561_, _26560_, _26557_);
  nor (_26562_, _10431_, _03518_);
  nor (_26563_, _26562_, _03759_);
  nand (_26564_, _26563_, _26561_);
  and (_26566_, _03759_, _03510_);
  nor (_26567_, _26566_, _10255_);
  nand (_26568_, _26567_, _26564_);
  and (_26569_, _04180_, _10255_);
  nor (_26570_, _26569_, _03758_);
  nand (_26571_, _26570_, _26568_);
  nor (_26572_, _26489_, _03427_);
  and (_26573_, _03758_, _03510_);
  nor (_26574_, _26573_, _26572_);
  and (_26575_, _26574_, _26571_);
  not (_26577_, _04306_);
  nor (_26578_, _26496_, _10476_);
  and (_26579_, _10476_, _10160_);
  nor (_26580_, _26579_, _26578_);
  and (_26581_, _26580_, _26577_);
  nor (_26582_, _26581_, _10441_);
  or (_26583_, _26582_, _26575_);
  and (_26584_, _26580_, _04306_);
  nor (_26585_, _26584_, _03925_);
  nand (_26586_, _26585_, _26583_);
  and (_26588_, _10249_, _10159_);
  not (_26589_, _26496_);
  nor (_26590_, _26589_, _10249_);
  or (_26591_, _26590_, _26588_);
  nor (_26592_, _26591_, _10444_);
  nor (_26593_, _26592_, _03868_);
  nand (_26594_, _26593_, _26586_);
  nor (_26595_, _26496_, _10498_);
  and (_26596_, _10498_, _10160_);
  or (_26597_, _26596_, _03918_);
  or (_26599_, _26597_, _26595_);
  nand (_26600_, _26599_, _26594_);
  nand (_26601_, _26600_, _10486_);
  nor (_26602_, _26589_, _10515_);
  and (_26603_, _10515_, _10159_);
  nor (_26604_, _26603_, _26602_);
  nor (_26605_, _26604_, _11857_);
  and (_26606_, _10485_, _03518_);
  nor (_26607_, _26606_, _26605_);
  and (_26608_, _26607_, _03753_);
  nand (_26610_, _26608_, _26601_);
  and (_26611_, _03752_, _03511_);
  nor (_26612_, _26611_, _05049_);
  nand (_26613_, _26612_, _26610_);
  nor (_26614_, _04180_, _03428_);
  nor (_26615_, _26614_, _26232_);
  and (_26616_, _26615_, _26613_);
  or (_26617_, _26616_, _26494_);
  nand (_26618_, _26617_, _10092_);
  nor (_26619_, _10092_, _03518_);
  nor (_26621_, _26619_, _03879_);
  nand (_26622_, _26621_, _26618_);
  and (_26623_, _03879_, _03510_);
  nor (_26624_, _26623_, _25949_);
  nand (_26625_, _26624_, _26622_);
  and (_26626_, _04180_, _25949_);
  nor (_26627_, _26626_, _03878_);
  nand (_26628_, _26627_, _26625_);
  and (_26629_, _03878_, _03510_);
  nor (_26630_, _26629_, _15018_);
  and (_26632_, _26630_, _26628_);
  nor (_26633_, _10087_, _03518_);
  or (_26634_, _26633_, _26632_);
  nand (_26635_, _26634_, _10085_);
  nor (_26636_, _10085_, _03510_);
  nor (_26637_, _26636_, _03425_);
  nand (_26638_, _26637_, _26635_);
  and (_26639_, _03518_, _03425_);
  nor (_26640_, _26639_, _03746_);
  and (_26641_, _26640_, _26638_);
  or (_26643_, _26641_, _26493_);
  nand (_26644_, _26643_, _06141_);
  and (_26645_, _04180_, _03456_);
  nor (_26646_, _26645_, _03921_);
  nand (_26647_, _26646_, _26644_);
  and (_26648_, _26647_, _26492_);
  or (_26649_, _26648_, _26490_);
  and (_26650_, _03831_, _03397_);
  nor (_26651_, _03737_, _26650_);
  nand (_26652_, _26490_, _03510_);
  and (_26654_, _26652_, _26651_);
  nand (_26655_, _26654_, _26649_);
  nor (_26656_, _26651_, _03510_);
  nor (_26657_, _26656_, _03455_);
  nand (_26658_, _26657_, _26655_);
  and (_26659_, _10159_, _03455_);
  nor (_26660_, _26659_, _10558_);
  nand (_26661_, _26660_, _26658_);
  nor (_26662_, _10556_, _03518_);
  nor (_26663_, _26662_, _03816_);
  and (_26665_, _26663_, _26661_);
  and (_26666_, _03816_, _03510_);
  or (_26667_, _26666_, _03398_);
  nor (_26668_, _26667_, _26665_);
  and (_26669_, _04180_, _03398_);
  or (_26670_, _26669_, _26668_);
  nand (_26671_, _26670_, _10565_);
  nor (_26672_, _26525_, _10565_);
  not (_26673_, _03400_);
  nor (_26674_, _10439_, _26673_);
  nor (_26676_, _26674_, _26672_);
  nand (_26677_, _26676_, _26671_);
  and (_26678_, _26674_, _03510_);
  nor (_26679_, _05009_, _26673_);
  nor (_26680_, _26679_, _26678_);
  nand (_26681_, _26680_, _26677_);
  and (_26682_, _26679_, _03511_);
  nor (_26683_, _26682_, _03903_);
  and (_26684_, _26683_, _26681_);
  and (_26685_, _10159_, _03903_);
  or (_26687_, _26685_, _08492_);
  nor (_26688_, _26687_, _26684_);
  and (_26689_, _08492_, _03511_);
  or (_26690_, _26689_, _26688_);
  nand (_26691_, _26690_, _10581_);
  and (_26692_, _10580_, _03529_);
  nor (_26693_, _26692_, _03815_);
  nand (_26694_, _26693_, _26691_);
  and (_26695_, _03815_, _03510_);
  nor (_26696_, _26695_, _03401_);
  nand (_26698_, _26696_, _26694_);
  and (_26699_, _04180_, _03401_);
  nor (_26700_, _26699_, _10620_);
  nand (_26701_, _26700_, _26698_);
  and (_26702_, _08826_, _03510_);
  and (_26703_, _26525_, _10627_);
  or (_26704_, _26703_, _26702_);
  and (_26705_, _26704_, _10620_);
  nor (_26706_, _26705_, _10625_);
  and (_26707_, _26706_, _26701_);
  or (_26709_, _26707_, _26487_);
  nand (_26710_, _26709_, _10079_);
  nor (_26711_, _10079_, _03510_);
  nor (_26712_, _26711_, _03897_);
  and (_26713_, _26712_, _26710_);
  and (_26714_, _10159_, _03897_);
  or (_26715_, _26714_, _04018_);
  nor (_26716_, _26715_, _26713_);
  and (_26717_, _04018_, _03511_);
  or (_26718_, _26717_, _26716_);
  nand (_26720_, _26718_, _25850_);
  and (_26721_, _04180_, _03405_);
  nor (_26722_, _26721_, _10643_);
  nand (_26723_, _26722_, _26720_);
  nor (_26724_, _26525_, _10627_);
  nor (_26725_, _08826_, _03510_);
  nor (_26726_, _26725_, _10644_);
  not (_26727_, _26726_);
  nor (_26728_, _26727_, _26724_);
  nor (_26729_, _26728_, _10656_);
  and (_26731_, _26729_, _26723_);
  or (_26732_, _26731_, _26486_);
  nand (_26733_, _26732_, _10658_);
  nor (_26734_, _10658_, _03510_);
  nor (_26735_, _26734_, _03908_);
  and (_26736_, _26735_, _26733_);
  and (_26737_, _10159_, _03908_);
  or (_26738_, _26737_, _04027_);
  nor (_26739_, _26738_, _26736_);
  and (_26740_, _04027_, _03511_);
  or (_26742_, _26740_, _26739_);
  nand (_26743_, _26742_, _25847_);
  and (_26744_, _04180_, _03388_);
  nor (_26745_, _26744_, _10074_);
  nand (_26746_, _26745_, _26743_);
  nor (_26747_, _26525_, \oc8051_golden_model_1.PSW [7]);
  nor (_26748_, _03510_, _08297_);
  nor (_26749_, _26748_, _10075_);
  not (_26750_, _26749_);
  nor (_26751_, _26750_, _26747_);
  nor (_26753_, _26751_, _10670_);
  and (_26754_, _26753_, _26746_);
  or (_26755_, _26754_, _26485_);
  nand (_26756_, _26755_, _08581_);
  nor (_26757_, _08581_, _03510_);
  nor (_26758_, _26757_, _03914_);
  and (_26759_, _26758_, _26756_);
  and (_26760_, _10159_, _03914_);
  or (_26761_, _26760_, _04011_);
  nor (_26762_, _26761_, _26759_);
  and (_26764_, _04011_, _03511_);
  or (_26765_, _26764_, _26762_);
  nand (_26766_, _26765_, _26042_);
  and (_26767_, _04180_, _03393_);
  nor (_26768_, _26767_, _10063_);
  nand (_26769_, _26768_, _26766_);
  nor (_26770_, _26525_, _08297_);
  nor (_26771_, _03510_, \oc8051_golden_model_1.PSW [7]);
  nor (_26772_, _26771_, _10064_);
  not (_26773_, _26772_);
  nor (_26775_, _26773_, _26770_);
  nor (_26776_, _26775_, _10688_);
  and (_26777_, _26776_, _26769_);
  or (_26778_, _26777_, _26484_);
  nand (_26779_, _26778_, _08628_);
  nor (_26780_, _08628_, _03510_);
  nor (_26781_, _26780_, _08657_);
  and (_26782_, _26781_, _26779_);
  and (_26783_, _08657_, _03518_);
  or (_26784_, _26783_, _04034_);
  nor (_26786_, _26784_, _26782_);
  and (_26787_, _06824_, _04034_);
  or (_26788_, _26787_, _26786_);
  nand (_26789_, _26788_, _03384_);
  and (_26790_, _04180_, _03383_);
  nor (_26791_, _26790_, _03913_);
  nand (_26792_, _26791_, _26789_);
  nor (_26793_, _10159_, _10906_);
  and (_26794_, _26589_, _10906_);
  or (_26795_, _26794_, _04097_);
  nor (_26797_, _26795_, _26793_);
  nor (_26798_, _26797_, _10712_);
  and (_26799_, _26798_, _26792_);
  or (_26800_, _26799_, _26483_);
  nand (_26801_, _26800_, _10056_);
  nor (_26802_, _10056_, _03510_);
  nor (_26803_, _26802_, _08772_);
  nand (_26804_, _26803_, _26801_);
  and (_26805_, _08772_, _03518_);
  nor (_26806_, _26805_, _03777_);
  and (_26808_, _26806_, _26804_);
  and (_26809_, _06824_, _03777_);
  or (_26810_, _26809_, _26808_);
  nand (_26811_, _26810_, _03411_);
  and (_26812_, _04180_, _03410_);
  nor (_26813_, _26812_, _03775_);
  nand (_26814_, _26813_, _26811_);
  nor (_26815_, _26496_, _10906_);
  and (_26816_, _10160_, _10906_);
  nor (_26817_, _26816_, _26815_);
  and (_26818_, _26817_, _03775_);
  nor (_26819_, _26818_, _10937_);
  nand (_26820_, _26819_, _26814_);
  nor (_26821_, _10936_, _03518_);
  nor (_26822_, _26821_, _03773_);
  and (_26823_, _26822_, _26820_);
  or (_26824_, _26823_, _26482_);
  nand (_26825_, _26824_, _10943_);
  nor (_26826_, _10943_, _03935_);
  nor (_26827_, _26826_, _05223_);
  nand (_26830_, _26827_, _26825_);
  and (_26831_, _05223_, _04180_);
  nor (_26832_, _26831_, _03374_);
  nand (_26833_, _26832_, _26830_);
  and (_26834_, _26817_, _03374_);
  nor (_26835_, _26834_, _10959_);
  nand (_26836_, _26835_, _26833_);
  nor (_26837_, _10958_, _03518_);
  nor (_26838_, _26837_, _03772_);
  and (_26839_, _26838_, _26836_);
  or (_26841_, _26839_, _26481_);
  nand (_26842_, _26841_, _10965_);
  nor (_26843_, _10965_, _03935_);
  nor (_26844_, _26843_, _25834_);
  nand (_26845_, _26844_, _26842_);
  and (_26846_, _25834_, _04180_);
  nor (_26847_, _26846_, _10042_);
  and (_26848_, _26847_, _26845_);
  or (_26849_, _26848_, _26480_);
  or (_26850_, _26849_, _43156_);
  or (_26852_, _43152_, \oc8051_golden_model_1.PC [2]);
  and (_26853_, _26852_, _41894_);
  and (_43511_, _26853_, _26850_);
  and (_26854_, _10042_, _03559_);
  and (_26855_, _03772_, _03552_);
  and (_26856_, _03773_, _03552_);
  nor (_26857_, _10059_, _03559_);
  and (_26858_, _06779_, _04034_);
  nor (_26859_, _10061_, _03559_);
  nor (_26860_, _10072_, _03559_);
  nor (_26862_, _10654_, _03559_);
  nor (_26863_, _10082_, _03559_);
  and (_26864_, _08492_, _03938_);
  and (_26865_, _03746_, _03938_);
  nor (_26866_, _10087_, _03559_);
  nor (_26867_, _26231_, _03552_);
  and (_26868_, _10485_, _03559_);
  nor (_26869_, _26868_, _03752_);
  or (_26870_, _10321_, _10320_);
  and (_26871_, _26870_, _10333_);
  nor (_26873_, _26870_, _10333_);
  nor (_26874_, _26873_, _26871_);
  and (_26875_, _26874_, _10383_);
  and (_26876_, _25887_, _03552_);
  nor (_26877_, _26876_, _26875_);
  or (_26878_, _26877_, _04266_);
  and (_26879_, _04005_, _03768_);
  nand (_26880_, _04230_, _03938_);
  nor (_26881_, _05011_, _03082_);
  or (_26882_, _26881_, _04707_);
  and (_26884_, _26882_, _26504_);
  and (_26885_, _05011_, _03559_);
  or (_26886_, _26885_, _26884_);
  and (_26887_, _26886_, _26880_);
  and (_26888_, _04263_, _03559_);
  or (_26889_, _26888_, _25875_);
  nor (_26890_, _26889_, _26887_);
  nor (_26891_, _10402_, _03559_);
  or (_26892_, _26891_, _04267_);
  or (_26893_, _26892_, _26890_);
  or (_26895_, _26893_, _26879_);
  and (_26896_, _26895_, _04717_);
  and (_26897_, _26896_, _26878_);
  and (_26898_, _04716_, _03558_);
  nor (_26899_, _26898_, _26897_);
  and (_26900_, _26899_, _04722_);
  or (_26901_, _10157_, _10156_);
  and (_26902_, _26901_, _10172_);
  nor (_26903_, _26901_, _10172_);
  nor (_26904_, _26903_, _26902_);
  nor (_26906_, _26904_, _25901_);
  and (_26907_, _25901_, _10155_);
  or (_26908_, _26907_, _04722_);
  nor (_26909_, _26908_, _26906_);
  or (_26910_, _26909_, _10413_);
  nor (_26911_, _26910_, _26900_);
  nor (_26912_, _10412_, _03559_);
  nor (_26913_, _26912_, _03763_);
  not (_26914_, _26913_);
  nor (_26915_, _26914_, _26911_);
  and (_26917_, _03763_, _03552_);
  or (_26918_, _26917_, _26915_);
  and (_26919_, _26918_, _03431_);
  nor (_26920_, _04005_, _03431_);
  or (_26921_, _26920_, _26919_);
  and (_26922_, _26921_, _04733_);
  and (_26923_, _03848_, _03552_);
  nor (_26924_, _26923_, _26168_);
  not (_26925_, _26924_);
  nor (_26926_, _26925_, _26922_);
  nor (_26927_, _10421_, _03559_);
  nor (_26928_, _26927_, _03854_);
  not (_26929_, _26928_);
  nor (_26930_, _26929_, _26926_);
  and (_26931_, _03854_, _03552_);
  nor (_26932_, _26931_, _10434_);
  not (_26933_, _26932_);
  nor (_26934_, _26933_, _26930_);
  nor (_26935_, _10431_, _03559_);
  nor (_26936_, _26935_, _03759_);
  not (_26939_, _26936_);
  or (_26940_, _26939_, _26934_);
  and (_26941_, _03759_, _03552_);
  nor (_26942_, _26941_, _10255_);
  nand (_26943_, _26942_, _26940_);
  and (_26944_, _04005_, _10255_);
  nor (_26945_, _26944_, _03758_);
  nand (_26946_, _26945_, _26943_);
  and (_26947_, _03758_, _03552_);
  nor (_26948_, _26947_, _10442_);
  and (_26950_, _26948_, _26946_);
  and (_26951_, _10476_, _10154_);
  not (_26952_, _26904_);
  nor (_26953_, _26952_, _10476_);
  or (_26954_, _26953_, _26951_);
  nor (_26955_, _26954_, _10441_);
  or (_26956_, _26955_, _26950_);
  nand (_26957_, _26956_, _10444_);
  and (_26958_, _10249_, _10154_);
  nor (_26959_, _26952_, _10249_);
  or (_26961_, _26959_, _10444_);
  or (_26962_, _26961_, _26958_);
  and (_26963_, _26962_, _03918_);
  nand (_26964_, _26963_, _26957_);
  nor (_26965_, _26904_, _10498_);
  and (_26966_, _10498_, _10155_);
  or (_26967_, _26966_, _03918_);
  or (_26968_, _26967_, _26965_);
  nand (_26969_, _26968_, _26964_);
  and (_26970_, _26969_, _10486_);
  nor (_26972_, _26904_, _10515_);
  and (_26973_, _10515_, _10155_);
  or (_26974_, _26973_, _11857_);
  nor (_26975_, _26974_, _26972_);
  nor (_26976_, _26975_, _26970_);
  nand (_26977_, _26976_, _26869_);
  and (_26978_, _03752_, _03938_);
  nor (_26979_, _26978_, _05049_);
  nand (_26980_, _26979_, _26977_);
  nor (_26981_, _04005_, _03428_);
  nor (_26983_, _26981_, _26232_);
  and (_26984_, _26983_, _26980_);
  or (_26985_, _26984_, _26867_);
  nand (_26986_, _26985_, _10092_);
  nor (_26987_, _10092_, _03559_);
  nor (_26988_, _26987_, _03879_);
  nand (_26989_, _26988_, _26986_);
  and (_26990_, _03879_, _03552_);
  nor (_26991_, _26990_, _25949_);
  nand (_26992_, _26991_, _26989_);
  and (_26994_, _04005_, _25949_);
  nor (_26995_, _26994_, _03878_);
  nand (_26996_, _26995_, _26992_);
  and (_26997_, _03878_, _03552_);
  nor (_26998_, _26997_, _15018_);
  and (_26999_, _26998_, _26996_);
  or (_27000_, _26999_, _26866_);
  nand (_27001_, _27000_, _10085_);
  nor (_27002_, _10085_, _03552_);
  nor (_27003_, _27002_, _03425_);
  nand (_27005_, _27003_, _27001_);
  and (_27006_, _03425_, _03559_);
  nor (_27007_, _27006_, _03746_);
  and (_27008_, _27007_, _27005_);
  or (_27009_, _27008_, _26865_);
  nand (_27010_, _27009_, _06141_);
  and (_27011_, _04005_, _03456_);
  nor (_27012_, _27011_, _03921_);
  nand (_27013_, _27012_, _27010_);
  and (_27014_, _10154_, _03921_);
  nor (_27016_, _27014_, _07927_);
  nand (_27017_, _27016_, _27013_);
  nor (_27018_, _07926_, _03552_);
  nor (_27019_, _27018_, _03455_);
  nand (_27020_, _27019_, _27017_);
  and (_27021_, _10154_, _03455_);
  nor (_27022_, _27021_, _10558_);
  nand (_27023_, _27022_, _27020_);
  nor (_27024_, _10556_, _03559_);
  nor (_27025_, _27024_, _03816_);
  and (_27027_, _27025_, _27023_);
  and (_27028_, _03816_, _03552_);
  or (_27029_, _27028_, _03398_);
  or (_27030_, _27029_, _27027_);
  and (_27031_, _04005_, _03398_);
  nor (_27032_, _27031_, _10564_);
  nand (_27033_, _27032_, _27030_);
  and (_27034_, _26874_, _10564_);
  nor (_27035_, _27034_, _06309_);
  nand (_27036_, _27035_, _27033_);
  nor (_27038_, _06138_, _03552_);
  nor (_27039_, _27038_, _03903_);
  nand (_27040_, _27039_, _27036_);
  and (_27041_, _10154_, _03903_);
  nor (_27042_, _27041_, _08492_);
  and (_27043_, _27042_, _27040_);
  or (_27044_, _27043_, _26864_);
  nand (_27045_, _27044_, _10581_);
  nor (_27046_, _10581_, _03571_);
  nor (_27047_, _27046_, _03815_);
  nand (_27049_, _27047_, _27045_);
  and (_27050_, _03815_, _03552_);
  nor (_27051_, _27050_, _03401_);
  nand (_27052_, _27051_, _27049_);
  and (_27053_, _04005_, _03401_);
  nor (_27054_, _27053_, _10620_);
  nand (_27055_, _27054_, _27052_);
  nor (_27056_, _26874_, _08826_);
  and (_27057_, _08826_, _03938_);
  nor (_27058_, _27057_, _10621_);
  not (_27060_, _27058_);
  nor (_27061_, _27060_, _27056_);
  nor (_27062_, _27061_, _10625_);
  and (_27063_, _27062_, _27055_);
  or (_27064_, _27063_, _26863_);
  nand (_27065_, _27064_, _10079_);
  nor (_27066_, _10079_, _03552_);
  nor (_27067_, _27066_, _03897_);
  and (_27068_, _27067_, _27065_);
  and (_27069_, _10154_, _03897_);
  or (_27071_, _27069_, _04018_);
  nor (_27072_, _27071_, _27068_);
  and (_27073_, _04018_, _03938_);
  or (_27074_, _27073_, _27072_);
  nand (_27075_, _27074_, _25850_);
  and (_27076_, _04005_, _03405_);
  nor (_27077_, _27076_, _10643_);
  nand (_27078_, _27077_, _27075_);
  nor (_27079_, _26874_, _10627_);
  nor (_27080_, _08826_, _03552_);
  nor (_27082_, _27080_, _10644_);
  not (_27083_, _27082_);
  nor (_27084_, _27083_, _27079_);
  nor (_27085_, _27084_, _10656_);
  and (_27086_, _27085_, _27078_);
  or (_27087_, _27086_, _26862_);
  nand (_27088_, _27087_, _10658_);
  nor (_27089_, _10658_, _03552_);
  nor (_27090_, _27089_, _03908_);
  and (_27091_, _27090_, _27088_);
  and (_27093_, _10154_, _03908_);
  or (_27094_, _27093_, _04027_);
  nor (_27095_, _27094_, _27091_);
  and (_27096_, _04027_, _03938_);
  or (_27097_, _27096_, _27095_);
  nand (_27098_, _27097_, _25847_);
  and (_27099_, _04005_, _03388_);
  nor (_27100_, _27099_, _10074_);
  nand (_27101_, _27100_, _27098_);
  nor (_27102_, _26874_, \oc8051_golden_model_1.PSW [7]);
  nor (_27104_, _03552_, _08297_);
  nor (_27105_, _27104_, _10075_);
  not (_27106_, _27105_);
  nor (_27107_, _27106_, _27102_);
  nor (_27108_, _27107_, _10670_);
  and (_27109_, _27108_, _27101_);
  or (_27110_, _27109_, _26860_);
  nand (_27111_, _27110_, _08581_);
  nor (_27112_, _08581_, _03552_);
  nor (_27113_, _27112_, _03914_);
  and (_27115_, _27113_, _27111_);
  and (_27116_, _10154_, _03914_);
  or (_27117_, _27116_, _04011_);
  nor (_27118_, _27117_, _27115_);
  and (_27119_, _04011_, _03938_);
  or (_27120_, _27119_, _27118_);
  nand (_27121_, _27120_, _26042_);
  and (_27122_, _04005_, _03393_);
  nor (_27123_, _27122_, _10063_);
  nand (_27124_, _27123_, _27121_);
  nor (_27126_, _26874_, _08297_);
  nor (_27127_, _03552_, \oc8051_golden_model_1.PSW [7]);
  nor (_27128_, _27127_, _10064_);
  not (_27129_, _27128_);
  nor (_27130_, _27129_, _27126_);
  nor (_27131_, _27130_, _10688_);
  and (_27132_, _27131_, _27124_);
  or (_27133_, _27132_, _26859_);
  nand (_27134_, _27133_, _08628_);
  nor (_27135_, _08628_, _03552_);
  nor (_27137_, _27135_, _08657_);
  nand (_27138_, _27137_, _27134_);
  and (_27139_, _08657_, _03559_);
  nor (_27140_, _27139_, _04034_);
  and (_27141_, _27140_, _27138_);
  or (_27142_, _27141_, _26858_);
  nand (_27143_, _27142_, _03384_);
  and (_27144_, _04005_, _03383_);
  nor (_27145_, _27144_, _03913_);
  nand (_27146_, _27145_, _27143_);
  and (_27147_, _26952_, _10906_);
  nor (_27148_, _10154_, _10906_);
  or (_27149_, _27148_, _04097_);
  nor (_27150_, _27149_, _27147_);
  nor (_27151_, _27150_, _10712_);
  and (_27152_, _27151_, _27146_);
  or (_27153_, _27152_, _26857_);
  nand (_27154_, _27153_, _10056_);
  nor (_27155_, _10056_, _03552_);
  nor (_27156_, _27155_, _08772_);
  and (_27159_, _27156_, _27154_);
  and (_27160_, _08772_, _03559_);
  or (_27161_, _27160_, _03777_);
  nor (_27162_, _27161_, _27159_);
  and (_27163_, _06779_, _03777_);
  or (_27164_, _27163_, _27162_);
  nand (_27165_, _27164_, _03411_);
  and (_27166_, _04005_, _03410_);
  nor (_27167_, _27166_, _03775_);
  nand (_27168_, _27167_, _27165_);
  nor (_27170_, _26904_, _10906_);
  and (_27171_, _10155_, _10906_);
  nor (_27172_, _27171_, _27170_);
  and (_27173_, _27172_, _03775_);
  nor (_27174_, _27173_, _10937_);
  nand (_27175_, _27174_, _27168_);
  nor (_27176_, _10936_, _03559_);
  nor (_27177_, _27176_, _03773_);
  and (_27178_, _27177_, _27175_);
  or (_27179_, _27178_, _26856_);
  nand (_27181_, _27179_, _10943_);
  nor (_27182_, _10943_, _03558_);
  nor (_27183_, _27182_, _05223_);
  nand (_27184_, _27183_, _27181_);
  and (_27185_, _05223_, _04005_);
  nor (_27186_, _27185_, _03374_);
  nand (_27187_, _27186_, _27184_);
  and (_27188_, _27172_, _03374_);
  nor (_27189_, _27188_, _10959_);
  nand (_27190_, _27189_, _27187_);
  nor (_27192_, _10958_, _03559_);
  nor (_27193_, _27192_, _03772_);
  and (_27194_, _27193_, _27190_);
  or (_27195_, _27194_, _26855_);
  nand (_27196_, _27195_, _10965_);
  nor (_27197_, _10965_, _03558_);
  nor (_27198_, _27197_, _25834_);
  nand (_27199_, _27198_, _27196_);
  and (_27200_, _25834_, _04005_);
  nor (_27201_, _27200_, _10042_);
  and (_27203_, _27201_, _27199_);
  or (_27204_, _27203_, _26854_);
  or (_27205_, _27204_, _43156_);
  or (_27206_, _43152_, \oc8051_golden_model_1.PC [3]);
  and (_27207_, _27206_, _41894_);
  and (_43512_, _27207_, _27205_);
  and (_27208_, _03103_, \oc8051_golden_model_1.PC [4]);
  nor (_27209_, _03103_, \oc8051_golden_model_1.PC [4]);
  nor (_27210_, _27209_, _27208_);
  and (_27211_, _27210_, _10042_);
  or (_27213_, _27210_, _10958_);
  nand (_27214_, _06442_, _03410_);
  nor (_27215_, _10150_, _10906_);
  and (_27216_, _10177_, _10174_);
  nor (_27217_, _27216_, _10178_);
  and (_27218_, _27217_, _10906_);
  or (_27219_, _27218_, _27215_);
  and (_27220_, _27219_, _03913_);
  nand (_27221_, _10318_, _03746_);
  nor (_27222_, _26231_, _10317_);
  not (_27224_, _10486_);
  and (_27225_, _10318_, _03759_);
  nor (_27226_, _27210_, _10421_);
  nor (_27227_, _27210_, _10417_);
  nor (_27228_, _27217_, _25901_);
  or (_27229_, _27228_, _04722_);
  and (_27230_, _10265_, _10150_);
  or (_27231_, _27230_, _27229_);
  and (_27232_, _06442_, _03768_);
  nor (_27233_, _05011_, \oc8051_golden_model_1.PC [4]);
  not (_27235_, _27210_);
  and (_27236_, _27235_, _05011_);
  or (_27237_, _27236_, _27233_);
  and (_27238_, _27237_, _04708_);
  and (_27239_, _10318_, _04707_);
  or (_27240_, _27239_, _04263_);
  or (_27241_, _27240_, _27238_);
  nand (_27242_, _27210_, _04263_);
  and (_27243_, _27242_, _03770_);
  and (_27244_, _27243_, _27241_);
  or (_27246_, _27244_, _26516_);
  or (_27247_, _27246_, _27232_);
  or (_27248_, _27235_, _10402_);
  and (_27249_, _27248_, _04266_);
  and (_27250_, _27249_, _27247_);
  and (_27251_, _10338_, _10335_);
  nor (_27252_, _27251_, _10339_);
  nand (_27253_, _27252_, _10383_);
  nand (_27254_, _10382_, _10317_);
  and (_27255_, _27254_, _27253_);
  and (_27257_, _27255_, _04267_);
  or (_27258_, _27257_, _27250_);
  and (_27259_, _27258_, _04717_);
  or (_27260_, _27259_, _03850_);
  and (_27261_, _27260_, _10412_);
  and (_27262_, _27261_, _27231_);
  or (_27263_, _27262_, _27227_);
  and (_27264_, _27263_, _03764_);
  and (_27265_, _10318_, _03763_);
  or (_27266_, _27265_, _05045_);
  or (_27268_, _27266_, _27264_);
  or (_27269_, _06442_, _03431_);
  and (_27270_, _27269_, _04733_);
  and (_27271_, _27270_, _27268_);
  and (_27272_, _10318_, _03848_);
  or (_27273_, _27272_, _27271_);
  and (_27274_, _27273_, _10421_);
  or (_27275_, _27274_, _27226_);
  and (_27276_, _27275_, _03855_);
  nand (_27277_, _10318_, _03854_);
  nand (_27279_, _27277_, _10431_);
  or (_27280_, _27279_, _27276_);
  or (_27281_, _27235_, _10431_);
  and (_27282_, _27281_, _03760_);
  and (_27283_, _27282_, _27280_);
  or (_27284_, _27283_, _27225_);
  and (_27285_, _27284_, _03434_);
  and (_27286_, _06442_, _10255_);
  or (_27287_, _27286_, _03758_);
  or (_27288_, _27287_, _27285_);
  and (_27290_, _10317_, _03758_);
  nor (_27291_, _27290_, _26572_);
  and (_27292_, _27291_, _27288_);
  and (_27293_, _10476_, _10150_);
  nor (_27294_, _27217_, _10476_);
  or (_27295_, _27294_, _27293_);
  or (_27296_, _27295_, _04306_);
  and (_27297_, _27296_, _10442_);
  or (_27298_, _27297_, _27292_);
  or (_27299_, _27295_, _26577_);
  and (_27301_, _27299_, _10444_);
  and (_27302_, _27301_, _27298_);
  nand (_27303_, _10249_, _10149_);
  not (_27304_, _27217_);
  or (_27305_, _27304_, _10249_);
  and (_27306_, _27305_, _03925_);
  and (_27307_, _27306_, _27303_);
  or (_27308_, _27307_, _03868_);
  or (_27309_, _27308_, _27302_);
  or (_27310_, _27304_, _10498_);
  nand (_27312_, _10498_, _10149_);
  and (_27313_, _27312_, _27310_);
  or (_27314_, _27313_, _03918_);
  and (_27315_, _27314_, _27309_);
  or (_27316_, _27315_, _27224_);
  nor (_27317_, _27217_, _10515_);
  and (_27318_, _10515_, _10150_);
  or (_27319_, _27318_, _11857_);
  or (_27320_, _27319_, _27317_);
  nand (_27321_, _27210_, _10485_);
  and (_27323_, _27321_, _03753_);
  and (_27324_, _27323_, _27320_);
  and (_27325_, _27324_, _27316_);
  and (_27326_, _10318_, _03752_);
  or (_27327_, _27326_, _05049_);
  or (_27328_, _27327_, _27325_);
  or (_27329_, _06442_, _03428_);
  and (_27330_, _27329_, _26231_);
  and (_27331_, _27330_, _27328_);
  or (_27332_, _27331_, _27222_);
  and (_27334_, _27332_, _10092_);
  nor (_27335_, _27210_, _10092_);
  or (_27336_, _27335_, _03879_);
  or (_27337_, _27336_, _27334_);
  nand (_27338_, _10317_, _03879_);
  and (_27339_, _27338_, _03441_);
  and (_27340_, _27339_, _27337_);
  and (_27341_, _06442_, _25949_);
  or (_27342_, _27341_, _03878_);
  or (_27343_, _27342_, _27340_);
  nand (_27345_, _10317_, _03878_);
  and (_27346_, _27345_, _27343_);
  nor (_27347_, _27346_, _15018_);
  nor (_27348_, _27235_, _10087_);
  or (_27349_, _27348_, _10086_);
  or (_27350_, _27349_, _27347_);
  or (_27351_, _10317_, _10085_);
  and (_27352_, _27351_, _03426_);
  and (_27353_, _27352_, _27350_);
  and (_27354_, _27210_, _03425_);
  or (_27356_, _27354_, _03746_);
  or (_27357_, _27356_, _27353_);
  and (_27358_, _27357_, _27221_);
  or (_27359_, _27358_, _03456_);
  nand (_27360_, _06442_, _03456_);
  and (_27361_, _27360_, _09861_);
  and (_27362_, _27361_, _27359_);
  nand (_27363_, _10149_, _03921_);
  nand (_27364_, _27363_, _07926_);
  or (_27365_, _27364_, _27362_);
  or (_27367_, _10317_, _07926_);
  and (_27368_, _27367_, _03820_);
  and (_27369_, _27368_, _27365_);
  nand (_27370_, _10149_, _03455_);
  nand (_27371_, _27370_, _10556_);
  or (_27372_, _27371_, _27369_);
  not (_27373_, _03816_);
  or (_27374_, _27210_, _10556_);
  and (_27375_, _27374_, _27373_);
  and (_27376_, _27375_, _27372_);
  nor (_27378_, _10317_, _03398_);
  nor (_27379_, _27378_, _10560_);
  or (_27380_, _27379_, _27376_);
  nand (_27381_, _06442_, _03398_);
  and (_27382_, _27381_, _10565_);
  and (_27383_, _27382_, _27380_);
  and (_27384_, _27252_, _10564_);
  or (_27385_, _27384_, _06309_);
  or (_27386_, _27385_, _27383_);
  or (_27387_, _10317_, _06138_);
  and (_27389_, _27387_, _04778_);
  and (_27390_, _27389_, _27386_);
  and (_27391_, _10149_, _03903_);
  or (_27392_, _27391_, _08492_);
  or (_27393_, _27392_, _27390_);
  nand (_27394_, _10318_, _08492_);
  and (_27395_, _27394_, _10581_);
  and (_27396_, _27395_, _27393_);
  nor (_27397_, _10597_, _10595_);
  nor (_27398_, _27397_, _10598_);
  and (_27400_, _27398_, _10580_);
  or (_27401_, _27400_, _03815_);
  or (_27402_, _27401_, _27396_);
  nand (_27403_, _10318_, _03815_);
  and (_27404_, _27403_, _27402_);
  or (_27405_, _27404_, _03401_);
  nand (_27406_, _06442_, _03401_);
  and (_27407_, _27406_, _10621_);
  and (_27408_, _27407_, _27405_);
  or (_27409_, _27252_, _08826_);
  nand (_27410_, _10318_, _08826_);
  and (_27411_, _27410_, _10620_);
  and (_27412_, _27411_, _27409_);
  or (_27413_, _27412_, _27408_);
  and (_27414_, _27413_, _10082_);
  nor (_27415_, _27235_, _10082_);
  or (_27416_, _27415_, _10080_);
  or (_27417_, _27416_, _27414_);
  or (_27418_, _10317_, _10079_);
  and (_27419_, _27418_, _04790_);
  and (_27422_, _27419_, _27417_);
  and (_27423_, _10149_, _03897_);
  or (_27424_, _27423_, _04018_);
  or (_27425_, _27424_, _27422_);
  nand (_27426_, _10318_, _04018_);
  and (_27427_, _27426_, _27425_);
  or (_27428_, _27427_, _03405_);
  nand (_27429_, _06442_, _03405_);
  and (_27430_, _27429_, _10644_);
  and (_27431_, _27430_, _27428_);
  or (_27433_, _27252_, _10627_);
  or (_27434_, _10317_, _08826_);
  and (_27435_, _27434_, _10643_);
  and (_27436_, _27435_, _27433_);
  or (_27437_, _27436_, _27431_);
  and (_27438_, _27437_, _10654_);
  nor (_27439_, _27235_, _10654_);
  or (_27440_, _27439_, _10659_);
  or (_27441_, _27440_, _27438_);
  or (_27442_, _10658_, _10317_);
  and (_27444_, _27442_, _03909_);
  and (_27445_, _27444_, _27441_);
  and (_27446_, _10149_, _03908_);
  or (_27447_, _27446_, _04027_);
  or (_27448_, _27447_, _27445_);
  nand (_27449_, _10318_, _04027_);
  and (_27450_, _27449_, _27448_);
  or (_27451_, _27450_, _03388_);
  nand (_27452_, _06442_, _03388_);
  and (_27453_, _27452_, _10075_);
  and (_27455_, _27453_, _27451_);
  or (_27456_, _27252_, \oc8051_golden_model_1.PSW [7]);
  or (_27457_, _10317_, _08297_);
  and (_27458_, _27457_, _10074_);
  and (_27459_, _27458_, _27456_);
  or (_27460_, _27459_, _27455_);
  and (_27461_, _27460_, _10072_);
  nor (_27462_, _27235_, _10072_);
  or (_27463_, _27462_, _08582_);
  or (_27464_, _27463_, _27461_);
  or (_27466_, _10317_, _08581_);
  and (_27467_, _27466_, _06567_);
  and (_27468_, _27467_, _27464_);
  and (_27469_, _10149_, _03914_);
  or (_27470_, _27469_, _04011_);
  or (_27471_, _27470_, _27468_);
  nand (_27472_, _10318_, _04011_);
  and (_27473_, _27472_, _27471_);
  or (_27474_, _27473_, _03393_);
  nand (_27475_, _06442_, _03393_);
  and (_27477_, _27475_, _10064_);
  and (_27478_, _27477_, _27474_);
  or (_27479_, _27252_, _08297_);
  or (_27480_, _10317_, \oc8051_golden_model_1.PSW [7]);
  and (_27481_, _27480_, _10063_);
  and (_27482_, _27481_, _27479_);
  or (_27483_, _27482_, _27478_);
  and (_27484_, _27483_, _10061_);
  nor (_27485_, _27235_, _10061_);
  or (_27486_, _27485_, _08629_);
  or (_27488_, _27486_, _27484_);
  or (_27489_, _10317_, _08628_);
  and (_27490_, _27489_, _08658_);
  and (_27491_, _27490_, _27488_);
  and (_27492_, _27210_, _08657_);
  or (_27493_, _27492_, _04034_);
  or (_27494_, _27493_, _27491_);
  or (_27495_, _06969_, _10704_);
  and (_27496_, _27495_, _27494_);
  or (_27497_, _27496_, _03383_);
  nand (_27499_, _06442_, _03383_);
  and (_27500_, _27499_, _04097_);
  and (_27501_, _27500_, _27497_);
  or (_27502_, _27501_, _27220_);
  and (_27503_, _27502_, _10059_);
  nor (_27504_, _27235_, _10059_);
  or (_27505_, _27504_, _10057_);
  or (_27506_, _27505_, _27503_);
  or (_27507_, _10317_, _10056_);
  and (_27508_, _27507_, _08773_);
  and (_27510_, _27508_, _27506_);
  and (_27511_, _27210_, _08772_);
  or (_27512_, _27511_, _03777_);
  or (_27513_, _27512_, _27510_);
  or (_27514_, _06969_, _03778_);
  and (_27515_, _27514_, _27513_);
  or (_27516_, _27515_, _03410_);
  and (_27517_, _27516_, _27214_);
  or (_27518_, _27517_, _03775_);
  or (_27519_, _27217_, _10906_);
  nand (_27521_, _10150_, _10906_);
  and (_27522_, _27521_, _27519_);
  or (_27523_, _27522_, _03776_);
  and (_27524_, _27523_, _10936_);
  and (_27525_, _27524_, _27518_);
  nor (_27526_, _27235_, _10936_);
  or (_27527_, _27526_, _03773_);
  or (_27528_, _27527_, _27525_);
  nand (_27529_, _10318_, _03773_);
  and (_27530_, _27529_, _10943_);
  and (_27532_, _27530_, _27528_);
  nor (_27533_, _27235_, _10943_);
  or (_27534_, _27533_, _05223_);
  or (_27535_, _27534_, _27532_);
  nand (_27536_, _06442_, _05223_);
  and (_27537_, _27536_, _03375_);
  and (_27538_, _27537_, _27535_);
  and (_27539_, _27522_, _03374_);
  or (_27540_, _27539_, _10959_);
  or (_27541_, _27540_, _27538_);
  and (_27543_, _27541_, _27213_);
  or (_27544_, _27543_, _03772_);
  nand (_27545_, _10318_, _03772_);
  and (_27546_, _27545_, _10965_);
  and (_27547_, _27546_, _27544_);
  nor (_27548_, _27235_, _10965_);
  or (_27549_, _27548_, _25834_);
  or (_27550_, _27549_, _27547_);
  nand (_27551_, _25834_, _06442_);
  and (_27552_, _27551_, _10976_);
  and (_27554_, _27552_, _27550_);
  or (_27555_, _27554_, _27211_);
  or (_27556_, _27555_, _43156_);
  or (_27557_, _43152_, \oc8051_golden_model_1.PC [4]);
  and (_27558_, _27557_, _41894_);
  and (_43513_, _27558_, _27556_);
  nor (_27559_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_27560_, _10312_, _03119_);
  nor (_27561_, _27560_, _27559_);
  and (_27562_, _27561_, _10042_);
  and (_27564_, _10312_, _03772_);
  and (_27565_, _10312_, _03773_);
  nor (_27566_, _27561_, _10059_);
  nor (_27567_, _27561_, _10061_);
  nor (_27568_, _27561_, _10072_);
  nor (_27569_, _27561_, _10654_);
  nor (_27570_, _27561_, _10082_);
  and (_27571_, _10144_, _03921_);
  nor (_27572_, _10312_, _10085_);
  nor (_27573_, _27561_, _10087_);
  nor (_27575_, _27561_, _10092_);
  nor (_27576_, _26231_, _10312_);
  nor (_27577_, _06411_, _03428_);
  and (_27578_, _27561_, _10485_);
  and (_27579_, _10515_, _10144_);
  or (_27580_, _10147_, _10146_);
  not (_27581_, _27580_);
  nor (_27582_, _27581_, _10179_);
  and (_27583_, _27581_, _10179_);
  nor (_27584_, _27583_, _27582_);
  nor (_27586_, _27584_, _10515_);
  or (_27587_, _27586_, _27579_);
  and (_27588_, _27587_, _03920_);
  and (_27589_, _25906_, _10144_);
  nor (_27590_, _27584_, _25906_);
  or (_27591_, _27590_, _27589_);
  and (_27592_, _27591_, _03850_);
  or (_27593_, _10315_, _10314_);
  and (_27594_, _27593_, _10340_);
  nor (_27595_, _27593_, _10340_);
  or (_27597_, _27595_, _27594_);
  nor (_27598_, _27597_, _10382_);
  and (_27599_, _25887_, _10312_);
  or (_27600_, _27599_, _27598_);
  and (_27601_, _27600_, _04267_);
  nand (_27602_, _06411_, _03768_);
  or (_27603_, _05011_, \oc8051_golden_model_1.PC [5]);
  not (_27604_, _27561_);
  nand (_27605_, _27604_, _05011_);
  and (_27606_, _27605_, _27603_);
  or (_27608_, _27606_, _04707_);
  nand (_27609_, _10313_, _04707_);
  and (_27610_, _27609_, _26504_);
  and (_27611_, _27610_, _27608_);
  and (_27612_, _27561_, _04263_);
  or (_27613_, _27612_, _25875_);
  or (_27614_, _27613_, _27611_);
  or (_27615_, _27561_, _10402_);
  and (_27616_, _27615_, _04266_);
  and (_27617_, _27616_, _27614_);
  and (_27619_, _27617_, _27602_);
  or (_27620_, _27619_, _04716_);
  or (_27621_, _27620_, _27601_);
  nand (_27622_, _27604_, _04716_);
  and (_27623_, _27622_, _04722_);
  and (_27624_, _27623_, _27621_);
  or (_27625_, _27624_, _10413_);
  or (_27626_, _27625_, _27592_);
  or (_27627_, _27561_, _10412_);
  and (_27628_, _27627_, _03764_);
  and (_27630_, _27628_, _27626_);
  and (_27631_, _10312_, _03763_);
  or (_27632_, _27631_, _05045_);
  or (_27633_, _27632_, _27630_);
  nand (_27634_, _06411_, _05045_);
  and (_27635_, _27634_, _04733_);
  and (_27636_, _27635_, _27633_);
  nand (_27637_, _10312_, _03848_);
  nand (_27638_, _27637_, _10421_);
  or (_27639_, _27638_, _27636_);
  or (_27641_, _27561_, _10421_);
  and (_27642_, _27641_, _03855_);
  and (_27643_, _27642_, _27639_);
  nand (_27644_, _10312_, _03854_);
  nand (_27645_, _27644_, _10431_);
  or (_27646_, _27645_, _27643_);
  or (_27647_, _27561_, _10431_);
  and (_27648_, _27647_, _03760_);
  and (_27649_, _27648_, _27646_);
  and (_27650_, _10312_, _03759_);
  or (_27652_, _27650_, _10255_);
  or (_27653_, _27652_, _27649_);
  nand (_27654_, _06411_, _10255_);
  and (_27655_, _27654_, _04845_);
  and (_27656_, _27655_, _27653_);
  nand (_27657_, _10476_, _10145_);
  not (_27658_, _27584_);
  or (_27659_, _27658_, _10476_);
  and (_27660_, _27659_, _27657_);
  and (_27661_, _27660_, _04306_);
  and (_27663_, _10312_, _03758_);
  or (_27664_, _27663_, _26572_);
  or (_27665_, _27664_, _27661_);
  or (_27666_, _27665_, _27656_);
  or (_27667_, _27660_, _10441_);
  and (_27668_, _27667_, _27666_);
  or (_27669_, _27668_, _03925_);
  or (_27670_, _27658_, _10249_);
  nand (_27671_, _10249_, _10145_);
  and (_27672_, _27671_, _27670_);
  or (_27674_, _27672_, _10444_);
  and (_27675_, _27674_, _27669_);
  and (_27676_, _27675_, _03918_);
  and (_27677_, _10498_, _10144_);
  nor (_27678_, _27584_, _10498_);
  or (_27679_, _27678_, _27677_);
  and (_27680_, _27679_, _03868_);
  or (_27681_, _27680_, _27676_);
  and (_27682_, _27681_, _11857_);
  nor (_27683_, _27682_, _27588_);
  nor (_27685_, _27683_, _10485_);
  or (_27686_, _27685_, _27578_);
  and (_27687_, _27686_, _03753_);
  and (_27688_, _10312_, _03752_);
  or (_27689_, _27688_, _27687_);
  and (_27690_, _27689_, _03428_);
  or (_27691_, _27690_, _26232_);
  nor (_27692_, _27691_, _27577_);
  nor (_27693_, _27692_, _27576_);
  nor (_27694_, _27693_, _10093_);
  or (_27695_, _27694_, _03879_);
  nor (_27696_, _27695_, _27575_);
  and (_27697_, _10312_, _03879_);
  nor (_27698_, _27697_, _27696_);
  nor (_27699_, _27698_, _25949_);
  nor (_27700_, _06411_, _03441_);
  or (_27701_, _27700_, _27699_);
  and (_27702_, _27701_, _11730_);
  and (_27703_, _10312_, _03878_);
  nor (_27704_, _27703_, _15018_);
  not (_27707_, _27704_);
  nor (_27708_, _27707_, _27702_);
  nor (_27709_, _27708_, _27573_);
  nor (_27710_, _27709_, _10086_);
  or (_27711_, _27710_, _03425_);
  nor (_27712_, _27711_, _27572_);
  and (_27713_, _27561_, _03425_);
  or (_27714_, _27713_, _03746_);
  or (_27715_, _27714_, _27712_);
  nand (_27716_, _10313_, _03746_);
  and (_27718_, _27716_, _27715_);
  and (_27719_, _27718_, _06141_);
  nor (_27720_, _06411_, _06141_);
  or (_27721_, _27720_, _27719_);
  and (_27722_, _27721_, _09861_);
  or (_27723_, _27722_, _07927_);
  or (_27724_, _27723_, _27571_);
  nor (_27725_, _10312_, _07926_);
  nor (_27726_, _27725_, _03455_);
  nand (_27727_, _27726_, _27724_);
  and (_27729_, _10144_, _03455_);
  nor (_27730_, _27729_, _10558_);
  nand (_27731_, _27730_, _27727_);
  nor (_27732_, _27561_, _10556_);
  nor (_27733_, _27732_, _03816_);
  and (_27734_, _27733_, _27731_);
  and (_27735_, _10312_, _03816_);
  or (_27736_, _27735_, _03398_);
  or (_27737_, _27736_, _27734_);
  and (_27738_, _06411_, _03398_);
  nor (_27740_, _27738_, _10564_);
  nand (_27741_, _27740_, _27737_);
  nor (_27742_, _27597_, _10565_);
  nor (_27743_, _27742_, _06309_);
  nand (_27744_, _27743_, _27741_);
  nor (_27745_, _10312_, _06138_);
  nor (_27746_, _27745_, _03903_);
  nand (_27747_, _27746_, _27744_);
  and (_27748_, _10144_, _03903_);
  nor (_27749_, _27748_, _08492_);
  nand (_27751_, _27749_, _27747_);
  and (_27752_, _10313_, _08492_);
  nor (_27753_, _27752_, _10580_);
  nand (_27754_, _27753_, _27751_);
  or (_27755_, _10592_, _10591_);
  and (_27756_, _27755_, _10599_);
  nor (_27757_, _27755_, _10599_);
  or (_27758_, _27757_, _27756_);
  nor (_27759_, _27758_, _10581_);
  nor (_27760_, _27759_, _03815_);
  and (_27762_, _27760_, _27754_);
  and (_27763_, _10313_, _03815_);
  or (_27764_, _27763_, _27762_);
  nand (_27765_, _27764_, _11641_);
  and (_27766_, _06411_, _03401_);
  nor (_27767_, _27766_, _10620_);
  nand (_27768_, _27767_, _27765_);
  and (_27769_, _10312_, _08826_);
  nor (_27770_, _27597_, _08826_);
  or (_27771_, _27770_, _27769_);
  and (_27773_, _27771_, _10620_);
  nor (_27774_, _27773_, _10625_);
  and (_27775_, _27774_, _27768_);
  or (_27776_, _27775_, _27570_);
  nand (_27777_, _27776_, _10079_);
  nor (_27778_, _10312_, _10079_);
  nor (_27779_, _27778_, _03897_);
  and (_27780_, _27779_, _27777_);
  and (_27781_, _10144_, _03897_);
  or (_27782_, _27781_, _04018_);
  nor (_27784_, _27782_, _27780_);
  and (_27785_, _10313_, _04018_);
  or (_27786_, _27785_, _27784_);
  nand (_27787_, _27786_, _25850_);
  and (_27788_, _06411_, _03405_);
  nor (_27789_, _27788_, _10643_);
  nand (_27790_, _27789_, _27787_);
  and (_27791_, _27597_, _08826_);
  nor (_27792_, _10312_, _08826_);
  nor (_27793_, _27792_, _10644_);
  not (_27795_, _27793_);
  nor (_27796_, _27795_, _27791_);
  nor (_27797_, _27796_, _10656_);
  and (_27798_, _27797_, _27790_);
  or (_27799_, _27798_, _27569_);
  nand (_27800_, _27799_, _10658_);
  nor (_27801_, _10658_, _10312_);
  nor (_27802_, _27801_, _03908_);
  and (_27803_, _27802_, _27800_);
  and (_27804_, _10144_, _03908_);
  or (_27806_, _27804_, _04027_);
  nor (_27807_, _27806_, _27803_);
  and (_27808_, _10313_, _04027_);
  or (_27809_, _27808_, _27807_);
  nand (_27810_, _27809_, _25847_);
  and (_27811_, _06411_, _03388_);
  nor (_27812_, _27811_, _10074_);
  nand (_27813_, _27812_, _27810_);
  and (_27814_, _27597_, _08297_);
  nor (_27815_, _10312_, _08297_);
  nor (_27817_, _27815_, _10075_);
  not (_27818_, _27817_);
  nor (_27819_, _27818_, _27814_);
  nor (_27820_, _27819_, _10670_);
  and (_27821_, _27820_, _27813_);
  or (_27822_, _27821_, _27568_);
  nand (_27823_, _27822_, _08581_);
  nor (_27824_, _10312_, _08581_);
  nor (_27825_, _27824_, _03914_);
  and (_27826_, _27825_, _27823_);
  and (_27828_, _10144_, _03914_);
  or (_27829_, _27828_, _04011_);
  nor (_27830_, _27829_, _27826_);
  and (_27831_, _10313_, _04011_);
  or (_27832_, _27831_, _27830_);
  nand (_27833_, _27832_, _26042_);
  and (_27834_, _06411_, _03393_);
  nor (_27835_, _27834_, _10063_);
  nand (_27836_, _27835_, _27833_);
  and (_27837_, _27597_, \oc8051_golden_model_1.PSW [7]);
  nor (_27839_, _10312_, \oc8051_golden_model_1.PSW [7]);
  nor (_27840_, _27839_, _10064_);
  not (_27841_, _27840_);
  nor (_27842_, _27841_, _27837_);
  nor (_27843_, _27842_, _10688_);
  and (_27844_, _27843_, _27836_);
  or (_27845_, _27844_, _27567_);
  nand (_27846_, _27845_, _08628_);
  nor (_27847_, _10312_, _08628_);
  nor (_27848_, _27847_, _08657_);
  and (_27850_, _27848_, _27846_);
  and (_27851_, _27561_, _08657_);
  or (_27852_, _27851_, _04034_);
  nor (_27853_, _27852_, _27850_);
  and (_27854_, _06873_, _04034_);
  or (_27855_, _27854_, _27853_);
  nand (_27856_, _27855_, _03384_);
  and (_27857_, _06411_, _03383_);
  nor (_27858_, _27857_, _03913_);
  nand (_27859_, _27858_, _27856_);
  and (_27861_, _27584_, _10906_);
  nor (_27862_, _10144_, _10906_);
  or (_27863_, _27862_, _04097_);
  or (_27864_, _27863_, _27861_);
  and (_27865_, _27864_, _10059_);
  and (_27866_, _27865_, _27859_);
  or (_27867_, _27866_, _27566_);
  nand (_27868_, _27867_, _10056_);
  nor (_27869_, _10312_, _10056_);
  nor (_27870_, _27869_, _08772_);
  and (_27872_, _27870_, _27868_);
  and (_27873_, _27561_, _08772_);
  or (_27874_, _27873_, _03777_);
  nor (_27875_, _27874_, _27872_);
  and (_27876_, _06873_, _03777_);
  or (_27877_, _27876_, _27875_);
  nand (_27878_, _27877_, _03411_);
  and (_27879_, _06411_, _03410_);
  nor (_27880_, _27879_, _03775_);
  nand (_27881_, _27880_, _27878_);
  and (_27883_, _10145_, _10906_);
  nor (_27884_, _27658_, _10906_);
  nor (_27885_, _27884_, _27883_);
  and (_27886_, _27885_, _03775_);
  nor (_27887_, _27886_, _10937_);
  nand (_27888_, _27887_, _27881_);
  nor (_27889_, _27561_, _10936_);
  nor (_27890_, _27889_, _03773_);
  and (_27891_, _27890_, _27888_);
  or (_27892_, _27891_, _27565_);
  nand (_27894_, _27892_, _10943_);
  nor (_27895_, _27604_, _10943_);
  nor (_27896_, _27895_, _05223_);
  nand (_27897_, _27896_, _27894_);
  and (_27898_, _06411_, _05223_);
  nor (_27899_, _27898_, _03374_);
  nand (_27900_, _27899_, _27897_);
  and (_27901_, _27885_, _03374_);
  nor (_27902_, _27901_, _10959_);
  nand (_27903_, _27902_, _27900_);
  nor (_27905_, _27561_, _10958_);
  nor (_27906_, _27905_, _03772_);
  and (_27907_, _27906_, _27903_);
  or (_27908_, _27907_, _27564_);
  nand (_27909_, _27908_, _10965_);
  nor (_27910_, _27604_, _10965_);
  nor (_27911_, _27910_, _25834_);
  nand (_27912_, _27911_, _27909_);
  and (_27913_, _25834_, _06411_);
  nor (_27914_, _27913_, _10042_);
  and (_27916_, _27914_, _27912_);
  or (_27917_, _27916_, _27562_);
  or (_27918_, _27917_, _43156_);
  or (_27919_, _43152_, \oc8051_golden_model_1.PC [5]);
  and (_27920_, _27919_, _41894_);
  and (_43514_, _27920_, _27918_);
  and (_27921_, _06252_, _03103_);
  nor (_27922_, _27921_, \oc8051_golden_model_1.PC [6]);
  nor (_27923_, _27922_, _10043_);
  and (_27924_, _27923_, _10042_);
  nand (_27926_, _06379_, _05223_);
  or (_27927_, _27923_, _08773_);
  nand (_27928_, _10138_, _03914_);
  nand (_27929_, _10138_, _03908_);
  nand (_27930_, _10138_, _03897_);
  or (_27931_, _10305_, _06138_);
  nand (_27932_, _10306_, _03816_);
  or (_27933_, _27923_, _10092_);
  nand (_27934_, _10306_, _03759_);
  or (_27935_, _27923_, _10421_);
  or (_27937_, _27923_, _10417_);
  nor (_27938_, _10182_, _10141_);
  nor (_27939_, _27938_, _10183_);
  or (_27940_, _27939_, _10265_);
  nand (_27941_, _10265_, _10138_);
  and (_27942_, _27941_, _03850_);
  and (_27943_, _27942_, _27940_);
  nand (_27944_, _06379_, _03768_);
  or (_27945_, _05011_, \oc8051_golden_model_1.PC [6]);
  or (_27946_, _27923_, _05012_);
  and (_27948_, _27946_, _27945_);
  or (_27949_, _27948_, _04707_);
  nand (_27950_, _10306_, _04707_);
  and (_27951_, _27950_, _26504_);
  and (_27952_, _27951_, _27949_);
  and (_27953_, _27923_, _04263_);
  or (_27954_, _27953_, _03768_);
  or (_27955_, _27954_, _27952_);
  and (_27956_, _27955_, _10402_);
  and (_27957_, _27956_, _27944_);
  and (_27959_, _27923_, _26516_);
  or (_27960_, _27959_, _04267_);
  or (_27961_, _27960_, _27957_);
  nor (_27962_, _10343_, _10309_);
  nor (_27963_, _27962_, _10344_);
  and (_27964_, _27963_, _10383_);
  and (_27965_, _10382_, _10305_);
  or (_27966_, _27965_, _27964_);
  or (_27967_, _27966_, _04266_);
  and (_27968_, _27967_, _27961_);
  or (_27970_, _27968_, _04716_);
  and (_27971_, _27970_, _04722_);
  or (_27972_, _27971_, _10413_);
  or (_27973_, _27972_, _27943_);
  and (_27974_, _27973_, _27937_);
  or (_27975_, _27974_, _03763_);
  nand (_27976_, _10306_, _03763_);
  and (_27977_, _27976_, _03431_);
  and (_27978_, _27977_, _27975_);
  nor (_27979_, _06379_, _03431_);
  or (_27981_, _27979_, _03848_);
  or (_27982_, _27981_, _27978_);
  nand (_27983_, _10306_, _03848_);
  and (_27984_, _27983_, _27982_);
  or (_27985_, _27984_, _26168_);
  and (_27986_, _27985_, _27935_);
  or (_27987_, _27986_, _03854_);
  nand (_27988_, _10306_, _03854_);
  and (_27989_, _27988_, _10431_);
  and (_27990_, _27989_, _27987_);
  and (_27992_, _27923_, _10434_);
  or (_27993_, _27992_, _03759_);
  or (_27994_, _27993_, _27990_);
  and (_27995_, _27994_, _27934_);
  or (_27996_, _27995_, _10255_);
  nand (_27997_, _06379_, _10255_);
  and (_27998_, _27997_, _04845_);
  and (_27999_, _27998_, _27996_);
  nand (_28000_, _10305_, _03758_);
  nand (_28001_, _28000_, _10441_);
  or (_28003_, _28001_, _27999_);
  not (_28004_, _10476_);
  and (_28005_, _27939_, _28004_);
  and (_28006_, _10476_, _10137_);
  or (_28007_, _28006_, _10441_);
  or (_28008_, _28007_, _28005_);
  and (_28009_, _28008_, _28003_);
  or (_28010_, _28009_, _03925_);
  or (_28011_, _27939_, _10249_);
  nand (_28012_, _10249_, _10138_);
  and (_28014_, _28012_, _28011_);
  or (_28015_, _28014_, _10444_);
  and (_28016_, _28015_, _28010_);
  or (_28017_, _28016_, _03868_);
  and (_28018_, _27939_, _10500_);
  and (_28019_, _10498_, _10137_);
  or (_28020_, _28019_, _03918_);
  or (_28021_, _28020_, _28018_);
  and (_28022_, _28021_, _10486_);
  and (_28023_, _28022_, _28017_);
  or (_28025_, _27939_, _10515_);
  nand (_28026_, _10515_, _10138_);
  and (_28027_, _28026_, _03920_);
  and (_28028_, _28027_, _28025_);
  and (_28029_, _27923_, _10485_);
  or (_28030_, _28029_, _03752_);
  or (_28031_, _28030_, _28028_);
  or (_28032_, _28031_, _28023_);
  nand (_28033_, _10306_, _03752_);
  and (_28034_, _28033_, _28032_);
  or (_28036_, _28034_, _05049_);
  nand (_28037_, _06379_, _05049_);
  and (_28038_, _28037_, _26231_);
  and (_28039_, _28038_, _28036_);
  nor (_28040_, _26231_, _10306_);
  or (_28041_, _28040_, _10093_);
  or (_28042_, _28041_, _28039_);
  and (_28043_, _28042_, _27933_);
  or (_28044_, _28043_, _03879_);
  nand (_28045_, _10306_, _03879_);
  and (_28047_, _28045_, _03441_);
  and (_28048_, _28047_, _28044_);
  nor (_28049_, _06379_, _03441_);
  or (_28050_, _28049_, _28048_);
  and (_28051_, _28050_, _11730_);
  nand (_28052_, _10305_, _03878_);
  nand (_28053_, _28052_, _10087_);
  or (_28054_, _28053_, _28051_);
  or (_28055_, _27923_, _10087_);
  and (_28056_, _28055_, _10085_);
  and (_28058_, _28056_, _28054_);
  nor (_28059_, _10306_, _10085_);
  or (_28060_, _28059_, _28058_);
  and (_28061_, _28060_, _03426_);
  and (_28062_, _27923_, _03425_);
  or (_28063_, _28062_, _03746_);
  or (_28064_, _28063_, _28061_);
  nand (_28065_, _10306_, _03746_);
  and (_28066_, _28065_, _06141_);
  and (_28067_, _28066_, _28064_);
  nor (_28069_, _06379_, _06141_);
  or (_28070_, _28069_, _03921_);
  or (_28071_, _28070_, _28067_);
  nand (_28072_, _10138_, _03921_);
  and (_28073_, _28072_, _07926_);
  and (_28074_, _28073_, _28071_);
  nor (_28075_, _10306_, _07926_);
  or (_28076_, _28075_, _03455_);
  or (_28077_, _28076_, _28074_);
  nand (_28078_, _10138_, _03455_);
  and (_28080_, _28078_, _10556_);
  and (_28081_, _28080_, _28077_);
  and (_28082_, _27923_, _10558_);
  or (_28083_, _28082_, _03816_);
  or (_28084_, _28083_, _28081_);
  and (_28085_, _28084_, _27932_);
  or (_28086_, _28085_, _03398_);
  nand (_28087_, _06379_, _03398_);
  and (_28088_, _28087_, _10565_);
  and (_28089_, _28088_, _28086_);
  and (_28091_, _27963_, _10564_);
  or (_28092_, _28091_, _06309_);
  or (_28093_, _28092_, _28089_);
  and (_28094_, _28093_, _27931_);
  or (_28095_, _28094_, _03903_);
  nand (_28096_, _10138_, _03903_);
  and (_28097_, _28096_, _08493_);
  and (_28098_, _28097_, _28095_);
  and (_28099_, _10305_, _08492_);
  or (_28100_, _28099_, _10580_);
  or (_28102_, _28100_, _28098_);
  nor (_28103_, _10602_, _10590_);
  nor (_28104_, _28103_, _10603_);
  or (_28105_, _28104_, _10581_);
  and (_28106_, _28105_, _04391_);
  and (_28107_, _28106_, _28102_);
  and (_28108_, _10305_, _03815_);
  or (_28109_, _28108_, _03401_);
  or (_28110_, _28109_, _28107_);
  nand (_28111_, _06379_, _03401_);
  and (_28113_, _28111_, _10621_);
  and (_28114_, _28113_, _28110_);
  or (_28115_, _27963_, _08826_);
  or (_28116_, _10305_, _10627_);
  and (_28117_, _28116_, _10620_);
  and (_28118_, _28117_, _28115_);
  or (_28119_, _28118_, _10625_);
  or (_28120_, _28119_, _28114_);
  or (_28121_, _27923_, _10082_);
  and (_28122_, _28121_, _10079_);
  and (_28124_, _28122_, _28120_);
  nor (_28125_, _10306_, _10079_);
  or (_28126_, _28125_, _03897_);
  or (_28127_, _28126_, _28124_);
  and (_28128_, _28127_, _27930_);
  or (_28129_, _28128_, _04018_);
  nand (_28130_, _10306_, _04018_);
  and (_28131_, _28130_, _25850_);
  and (_28132_, _28131_, _28129_);
  nor (_28133_, _06379_, _25850_);
  or (_28134_, _28133_, _28132_);
  and (_28135_, _28134_, _10644_);
  or (_28136_, _27963_, _10627_);
  or (_28137_, _10305_, _08826_);
  and (_28138_, _28137_, _10643_);
  and (_28139_, _28138_, _28136_);
  or (_28140_, _28139_, _10656_);
  or (_28141_, _28140_, _28135_);
  or (_28142_, _27923_, _10654_);
  and (_28143_, _28142_, _10658_);
  and (_28146_, _28143_, _28141_);
  nor (_28147_, _10658_, _10306_);
  or (_28148_, _28147_, _03908_);
  or (_28149_, _28148_, _28146_);
  and (_28150_, _28149_, _27929_);
  or (_28151_, _28150_, _04027_);
  nand (_28152_, _10306_, _04027_);
  and (_28153_, _28152_, _25847_);
  and (_28154_, _28153_, _28151_);
  nor (_28155_, _06379_, _25847_);
  or (_28157_, _28155_, _28154_);
  and (_28158_, _28157_, _10075_);
  or (_28159_, _27963_, \oc8051_golden_model_1.PSW [7]);
  or (_28160_, _10305_, _08297_);
  and (_28161_, _28160_, _10074_);
  and (_28162_, _28161_, _28159_);
  or (_28163_, _28162_, _10670_);
  or (_28164_, _28163_, _28158_);
  or (_28165_, _27923_, _10072_);
  and (_28166_, _28165_, _08581_);
  and (_28168_, _28166_, _28164_);
  nor (_28169_, _10306_, _08581_);
  or (_28170_, _28169_, _03914_);
  or (_28171_, _28170_, _28168_);
  and (_28172_, _28171_, _27928_);
  or (_28173_, _28172_, _04011_);
  nand (_28174_, _10306_, _04011_);
  and (_28175_, _28174_, _26042_);
  and (_28176_, _28175_, _28173_);
  nor (_28177_, _06379_, _26042_);
  or (_28179_, _28177_, _28176_);
  and (_28180_, _28179_, _10064_);
  or (_28181_, _27963_, _08297_);
  or (_28182_, _10305_, \oc8051_golden_model_1.PSW [7]);
  and (_28183_, _28182_, _10063_);
  and (_28184_, _28183_, _28181_);
  or (_28185_, _28184_, _10688_);
  or (_28186_, _28185_, _28180_);
  or (_28187_, _27923_, _10061_);
  and (_28188_, _28187_, _08628_);
  and (_28190_, _28188_, _28186_);
  nor (_28191_, _10306_, _08628_);
  or (_28192_, _28191_, _08657_);
  or (_28193_, _28192_, _28190_);
  or (_28194_, _27923_, _08658_);
  and (_28195_, _28194_, _10704_);
  and (_28196_, _28195_, _28193_);
  and (_28197_, _06641_, _04034_);
  or (_28198_, _28197_, _03383_);
  or (_28199_, _28198_, _28196_);
  nand (_28201_, _06379_, _03383_);
  and (_28202_, _28201_, _04097_);
  and (_28203_, _28202_, _28199_);
  or (_28204_, _27939_, _10907_);
  or (_28205_, _10137_, _10906_);
  and (_28206_, _28205_, _03913_);
  and (_28207_, _28206_, _28204_);
  or (_28208_, _28207_, _10712_);
  or (_28209_, _28208_, _28203_);
  or (_28210_, _27923_, _10059_);
  and (_28212_, _28210_, _10056_);
  and (_28213_, _28212_, _28209_);
  nor (_28214_, _10306_, _10056_);
  or (_28215_, _28214_, _08772_);
  or (_28216_, _28215_, _28213_);
  and (_28217_, _28216_, _27927_);
  or (_28218_, _28217_, _03777_);
  or (_28219_, _06641_, _03778_);
  and (_28220_, _28219_, _03411_);
  and (_28221_, _28220_, _28218_);
  nor (_28223_, _06379_, _03411_);
  or (_28224_, _28223_, _03775_);
  or (_28225_, _28224_, _28221_);
  or (_28226_, _27939_, _10906_);
  nand (_28227_, _10138_, _10906_);
  and (_28228_, _28227_, _28226_);
  or (_28229_, _28228_, _03776_);
  and (_28230_, _28229_, _28225_);
  or (_28231_, _28230_, _10937_);
  or (_28232_, _27923_, _10936_);
  and (_28234_, _28232_, _28231_);
  or (_28235_, _28234_, _03773_);
  nand (_28236_, _10306_, _03773_);
  and (_28237_, _28236_, _10943_);
  and (_28238_, _28237_, _28235_);
  and (_28239_, _27923_, _26446_);
  or (_28240_, _28239_, _05223_);
  or (_28241_, _28240_, _28238_);
  and (_28242_, _28241_, _27926_);
  or (_28243_, _28242_, _03374_);
  or (_28245_, _28228_, _03375_);
  and (_28246_, _28245_, _10958_);
  and (_28247_, _28246_, _28243_);
  and (_28248_, _27923_, _10959_);
  or (_28249_, _28248_, _03772_);
  or (_28250_, _28249_, _28247_);
  nand (_28251_, _10306_, _03772_);
  and (_28252_, _28251_, _10965_);
  and (_28253_, _28252_, _28250_);
  not (_28254_, _10965_);
  and (_28256_, _27923_, _28254_);
  or (_28257_, _28256_, _25834_);
  or (_28258_, _28257_, _28253_);
  nand (_28259_, _25834_, _06379_);
  and (_28260_, _28259_, _10976_);
  and (_28261_, _28260_, _28258_);
  or (_28262_, _28261_, _27924_);
  or (_28263_, _28262_, _43156_);
  or (_28264_, _43152_, \oc8051_golden_model_1.PC [6]);
  and (_28265_, _28264_, _41894_);
  and (_43515_, _28265_, _28263_);
  nor (_28267_, _10043_, \oc8051_golden_model_1.PC [7]);
  nor (_28268_, _28267_, _10044_);
  and (_28269_, _28268_, _10042_);
  and (_28270_, _06257_, _03772_);
  and (_28271_, _06257_, _03773_);
  nor (_28272_, _28268_, _10059_);
  nor (_28273_, _28268_, _10061_);
  nor (_28274_, _28268_, _10072_);
  nor (_28275_, _28268_, _10654_);
  nor (_28277_, _28268_, _10082_);
  and (_28278_, _06258_, _03746_);
  nor (_28279_, _28268_, _10087_);
  nor (_28280_, _26231_, _06257_);
  and (_28281_, _06257_, _03758_);
  or (_28282_, _10301_, _10302_);
  and (_28283_, _28282_, _10345_);
  nor (_28284_, _28282_, _10345_);
  nor (_28285_, _28284_, _28283_);
  and (_28286_, _28285_, _10383_);
  and (_28288_, _25887_, _06257_);
  nor (_28289_, _28288_, _28286_);
  or (_28290_, _28289_, _04266_);
  and (_28291_, _06342_, _03768_);
  nor (_28292_, _05011_, \oc8051_golden_model_1.PC [7]);
  not (_28293_, _28268_);
  and (_28294_, _28293_, _05011_);
  nor (_28295_, _28294_, _28292_);
  and (_28296_, _28295_, _04708_);
  and (_28297_, _06257_, _04707_);
  or (_28299_, _28297_, _28296_);
  and (_28300_, _28299_, _26504_);
  and (_28301_, _28268_, _04263_);
  or (_28302_, _28301_, _25875_);
  nor (_28303_, _28302_, _28300_);
  nor (_28304_, _28268_, _10402_);
  or (_28305_, _28304_, _04267_);
  or (_28306_, _28305_, _28303_);
  or (_28307_, _28306_, _28291_);
  and (_28308_, _28307_, _04717_);
  and (_28310_, _28308_, _28290_);
  and (_28311_, _28293_, _04716_);
  nor (_28312_, _28311_, _28310_);
  and (_28313_, _28312_, _04722_);
  and (_28314_, _25906_, _06935_);
  or (_28315_, _10133_, _10134_);
  and (_28316_, _28315_, _10184_);
  nor (_28317_, _28315_, _10184_);
  or (_28318_, _28317_, _28316_);
  nor (_28319_, _28318_, _25906_);
  nor (_28320_, _28319_, _28314_);
  nor (_28321_, _28320_, _04722_);
  or (_28322_, _28321_, _10413_);
  nor (_28323_, _28322_, _28313_);
  nor (_28324_, _28268_, _10412_);
  nor (_28325_, _28324_, _03763_);
  not (_28326_, _28325_);
  nor (_28327_, _28326_, _28323_);
  and (_28328_, _06257_, _03763_);
  or (_28329_, _28328_, _28327_);
  and (_28332_, _28329_, _03431_);
  nor (_28333_, _06342_, _03431_);
  or (_28334_, _28333_, _28332_);
  and (_28335_, _28334_, _04733_);
  and (_28336_, _06257_, _03848_);
  nor (_28337_, _28336_, _26168_);
  not (_28338_, _28337_);
  nor (_28339_, _28338_, _28335_);
  nor (_28340_, _28268_, _10421_);
  nor (_28341_, _28340_, _03854_);
  not (_28343_, _28341_);
  nor (_28344_, _28343_, _28339_);
  and (_28345_, _06257_, _03854_);
  nor (_28346_, _28345_, _10434_);
  not (_28347_, _28346_);
  nor (_28348_, _28347_, _28344_);
  nor (_28349_, _28268_, _10431_);
  nor (_28350_, _28349_, _03759_);
  not (_28351_, _28350_);
  nor (_28352_, _28351_, _28348_);
  and (_28354_, _06257_, _03759_);
  or (_28355_, _28354_, _28352_);
  and (_28356_, _28355_, _03434_);
  nor (_28357_, _06342_, _03434_);
  or (_28358_, _28357_, _28356_);
  and (_28359_, _28358_, _04845_);
  or (_28360_, _28359_, _10442_);
  nor (_28361_, _28360_, _28281_);
  and (_28362_, _10476_, _06935_);
  nor (_28363_, _28318_, _10476_);
  or (_28365_, _28363_, _28362_);
  nor (_28366_, _28365_, _10441_);
  or (_28367_, _28366_, _28361_);
  nand (_28368_, _28367_, _10444_);
  and (_28369_, _10249_, _06935_);
  nor (_28370_, _28318_, _10249_);
  or (_28371_, _28370_, _10444_);
  nor (_28372_, _28371_, _28369_);
  nor (_28373_, _28372_, _03868_);
  nand (_28374_, _28373_, _28368_);
  and (_28376_, _28318_, _10500_);
  and (_28377_, _10498_, _06936_);
  or (_28378_, _28377_, _03918_);
  or (_28379_, _28378_, _28376_);
  nand (_28380_, _28379_, _28374_);
  nand (_28381_, _28380_, _10486_);
  and (_28382_, _10515_, _06935_);
  nor (_28383_, _28318_, _10515_);
  or (_28384_, _28383_, _28382_);
  and (_28385_, _28384_, _03920_);
  and (_28387_, _28268_, _10485_);
  nor (_28388_, _28387_, _28385_);
  and (_28389_, _28388_, _03753_);
  nand (_28390_, _28389_, _28381_);
  and (_28391_, _06258_, _03752_);
  nor (_28392_, _28391_, _05049_);
  nand (_28393_, _28392_, _28390_);
  nor (_28394_, _06342_, _03428_);
  nor (_28395_, _28394_, _26232_);
  and (_28396_, _28395_, _28393_);
  or (_28398_, _28396_, _28280_);
  nand (_28399_, _28398_, _10092_);
  nor (_28400_, _28268_, _10092_);
  nor (_28401_, _28400_, _03879_);
  nand (_28402_, _28401_, _28399_);
  and (_28403_, _06257_, _03879_);
  nor (_28404_, _28403_, _25949_);
  nand (_28405_, _28404_, _28402_);
  and (_28406_, _06342_, _25949_);
  nor (_28407_, _28406_, _03878_);
  nand (_28409_, _28407_, _28405_);
  and (_28410_, _06257_, _03878_);
  nor (_28411_, _28410_, _15018_);
  and (_28412_, _28411_, _28409_);
  or (_28413_, _28412_, _28279_);
  nand (_28414_, _28413_, _10085_);
  nor (_28415_, _10085_, _06257_);
  nor (_28416_, _28415_, _03425_);
  nand (_28417_, _28416_, _28414_);
  and (_28418_, _28268_, _03425_);
  nor (_28420_, _28418_, _03746_);
  and (_28421_, _28420_, _28417_);
  or (_28422_, _28421_, _28278_);
  nand (_28423_, _28422_, _06141_);
  and (_28424_, _06342_, _03456_);
  nor (_28425_, _28424_, _03921_);
  nand (_28426_, _28425_, _28423_);
  and (_28427_, _06935_, _03921_);
  nor (_28428_, _28427_, _07927_);
  nand (_28429_, _28428_, _28426_);
  nor (_28431_, _07926_, _06257_);
  nor (_28432_, _28431_, _03455_);
  nand (_28433_, _28432_, _28429_);
  and (_28434_, _06935_, _03455_);
  nor (_28435_, _28434_, _10558_);
  nand (_28436_, _28435_, _28433_);
  nor (_28437_, _28268_, _10556_);
  nor (_28438_, _28437_, _03816_);
  nand (_28439_, _28438_, _28436_);
  nor (_28440_, _06257_, _03398_);
  or (_28442_, _28440_, _10560_);
  nand (_28443_, _28442_, _28439_);
  and (_28444_, _06342_, _03398_);
  nor (_28445_, _28444_, _10564_);
  nand (_28446_, _28445_, _28443_);
  and (_28447_, _28285_, _10564_);
  nor (_28448_, _28447_, _06309_);
  nand (_28449_, _28448_, _28446_);
  nor (_28450_, _06257_, _06138_);
  nor (_28451_, _28450_, _03903_);
  nand (_28453_, _28451_, _28449_);
  and (_28454_, _06935_, _03903_);
  nor (_28455_, _28454_, _08492_);
  nand (_28456_, _28455_, _28453_);
  and (_28457_, _08492_, _06258_);
  nor (_28458_, _28457_, _10580_);
  nand (_28459_, _28458_, _28456_);
  or (_28460_, _10587_, _10586_);
  nor (_28461_, _28460_, _10604_);
  and (_28462_, _28460_, _10604_);
  nor (_28464_, _28462_, _28461_);
  and (_28465_, _28464_, _10580_);
  nor (_28466_, _28465_, _03815_);
  and (_28467_, _28466_, _28459_);
  and (_28468_, _06258_, _03815_);
  or (_28469_, _28468_, _28467_);
  nand (_28470_, _28469_, _11641_);
  and (_28471_, _06342_, _03401_);
  nor (_28472_, _28471_, _10620_);
  nand (_28473_, _28472_, _28470_);
  and (_28475_, _08826_, _06257_);
  and (_28476_, _28285_, _10627_);
  or (_28477_, _28476_, _28475_);
  and (_28478_, _28477_, _10620_);
  nor (_28479_, _28478_, _10625_);
  and (_28480_, _28479_, _28473_);
  or (_28481_, _28480_, _28277_);
  nand (_28482_, _28481_, _10079_);
  nor (_28483_, _10079_, _06257_);
  nor (_28484_, _28483_, _03897_);
  and (_28486_, _28484_, _28482_);
  and (_28487_, _06935_, _03897_);
  or (_28488_, _28487_, _04018_);
  nor (_28489_, _28488_, _28486_);
  and (_28490_, _06258_, _04018_);
  or (_28491_, _28490_, _28489_);
  nand (_28492_, _28491_, _25850_);
  and (_28493_, _06342_, _03405_);
  nor (_28494_, _28493_, _10643_);
  nand (_28495_, _28494_, _28492_);
  nor (_28497_, _28285_, _10627_);
  nor (_28498_, _08826_, _06257_);
  nor (_28499_, _28498_, _10644_);
  not (_28500_, _28499_);
  nor (_28501_, _28500_, _28497_);
  nor (_28502_, _28501_, _10656_);
  and (_28503_, _28502_, _28495_);
  or (_28504_, _28503_, _28275_);
  nand (_28505_, _28504_, _10658_);
  nor (_28506_, _10658_, _06257_);
  nor (_28508_, _28506_, _03908_);
  and (_28509_, _28508_, _28505_);
  and (_28510_, _06935_, _03908_);
  or (_28511_, _28510_, _04027_);
  nor (_28512_, _28511_, _28509_);
  and (_28513_, _06258_, _04027_);
  or (_28514_, _28513_, _28512_);
  nand (_28515_, _28514_, _25847_);
  and (_28516_, _06342_, _03388_);
  nor (_28517_, _28516_, _10074_);
  nand (_28519_, _28517_, _28515_);
  nor (_28520_, _28285_, \oc8051_golden_model_1.PSW [7]);
  nor (_28521_, _06257_, _08297_);
  nor (_28522_, _28521_, _10075_);
  not (_28523_, _28522_);
  nor (_28524_, _28523_, _28520_);
  nor (_28525_, _28524_, _10670_);
  and (_28526_, _28525_, _28519_);
  or (_28527_, _28526_, _28274_);
  nand (_28528_, _28527_, _08581_);
  nor (_28530_, _08581_, _06257_);
  nor (_28531_, _28530_, _03914_);
  and (_28532_, _28531_, _28528_);
  and (_28533_, _06935_, _03914_);
  or (_28534_, _28533_, _04011_);
  nor (_28535_, _28534_, _28532_);
  and (_28536_, _06258_, _04011_);
  or (_28537_, _28536_, _28535_);
  nand (_28538_, _28537_, _26042_);
  and (_28539_, _06342_, _03393_);
  nor (_28541_, _28539_, _10063_);
  nand (_28542_, _28541_, _28538_);
  nor (_28543_, _28285_, _08297_);
  nor (_28544_, _06257_, \oc8051_golden_model_1.PSW [7]);
  nor (_28545_, _28544_, _10064_);
  not (_28546_, _28545_);
  nor (_28547_, _28546_, _28543_);
  nor (_28548_, _28547_, _10688_);
  and (_28549_, _28548_, _28542_);
  or (_28550_, _28549_, _28273_);
  nand (_28552_, _28550_, _08628_);
  nor (_28553_, _08628_, _06257_);
  nor (_28554_, _28553_, _08657_);
  nand (_28555_, _28554_, _28552_);
  and (_28556_, _28268_, _08657_);
  nor (_28557_, _28556_, _04034_);
  and (_28558_, _28557_, _28555_);
  nor (_28559_, _06248_, _10704_);
  or (_28560_, _28559_, _28558_);
  nand (_28561_, _28560_, _03384_);
  and (_28563_, _06342_, _03383_);
  nor (_28564_, _28563_, _03913_);
  nand (_28565_, _28564_, _28561_);
  and (_28566_, _28318_, _10906_);
  nor (_28567_, _06935_, _10906_);
  or (_28568_, _28567_, _04097_);
  or (_28569_, _28568_, _28566_);
  and (_28570_, _28569_, _10059_);
  and (_28571_, _28570_, _28565_);
  or (_28572_, _28571_, _28272_);
  nand (_28574_, _28572_, _10056_);
  nor (_28575_, _10056_, _06257_);
  nor (_28576_, _28575_, _08772_);
  and (_28577_, _28576_, _28574_);
  and (_28578_, _28268_, _08772_);
  or (_28579_, _28578_, _03777_);
  nor (_28580_, _28579_, _28577_);
  nor (_28581_, _06248_, _03778_);
  or (_28582_, _28581_, _28580_);
  nand (_28583_, _28582_, _03411_);
  and (_28585_, _06342_, _03410_);
  nor (_28586_, _28585_, _03775_);
  nand (_28587_, _28586_, _28583_);
  and (_28588_, _06935_, _10906_);
  nor (_28589_, _28318_, _10906_);
  or (_28590_, _28589_, _28588_);
  and (_28591_, _28590_, _03775_);
  nor (_28592_, _28591_, _10937_);
  nand (_28593_, _28592_, _28587_);
  nor (_28594_, _28268_, _10936_);
  nor (_28596_, _28594_, _03773_);
  and (_28597_, _28596_, _28593_);
  or (_28598_, _28597_, _28271_);
  nand (_28599_, _28598_, _10943_);
  nor (_28600_, _28293_, _10943_);
  nor (_28601_, _28600_, _05223_);
  nand (_28602_, _28601_, _28599_);
  and (_28603_, _06342_, _05223_);
  nor (_28604_, _28603_, _03374_);
  nand (_28605_, _28604_, _28602_);
  and (_28607_, _28590_, _03374_);
  nor (_28608_, _28607_, _10959_);
  nand (_28609_, _28608_, _28605_);
  nor (_28610_, _28268_, _10958_);
  nor (_28611_, _28610_, _03772_);
  and (_28612_, _28611_, _28609_);
  or (_28613_, _28612_, _28270_);
  nand (_28614_, _28613_, _10965_);
  nor (_28615_, _28293_, _10965_);
  nor (_28616_, _28615_, _25834_);
  nand (_28618_, _28616_, _28614_);
  and (_28619_, _25834_, _06342_);
  nor (_28620_, _28619_, _10042_);
  and (_28621_, _28620_, _28618_);
  or (_28622_, _28621_, _28269_);
  or (_28623_, _28622_, _43156_);
  or (_28624_, _43152_, \oc8051_golden_model_1.PC [7]);
  and (_28625_, _28624_, _41894_);
  and (_43516_, _28625_, _28623_);
  nor (_28626_, _03715_, _10969_);
  nor (_28628_, _03715_, _03900_);
  nor (_28629_, _10044_, \oc8051_golden_model_1.PC [8]);
  nor (_28630_, _28629_, _10045_);
  not (_28631_, _28630_);
  and (_28632_, _28631_, _08772_);
  or (_28633_, _28632_, _03777_);
  and (_28634_, _10189_, _03914_);
  nor (_28635_, _28630_, _10072_);
  nor (_28636_, _10074_, _03388_);
  not (_28637_, _28636_);
  nor (_28639_, _28630_, _10082_);
  nor (_28640_, _10349_, _06138_);
  and (_28641_, _10349_, _03816_);
  nor (_28642_, _28630_, _10556_);
  and (_28643_, _10188_, _03455_);
  and (_28644_, _10249_, _10188_);
  nor (_28645_, _10192_, _10186_);
  nor (_28646_, _28645_, _10193_);
  not (_28647_, _28646_);
  nor (_28648_, _28647_, _10249_);
  or (_28650_, _28648_, _10444_);
  or (_28651_, _28650_, _28644_);
  and (_28652_, _10349_, _03759_);
  and (_28653_, _25901_, _10188_);
  nor (_28654_, _28647_, _25901_);
  or (_28655_, _28654_, _04722_);
  or (_28656_, _28655_, _28653_);
  nand (_28657_, _28631_, _04716_);
  nor (_28658_, _10352_, _10347_);
  nor (_28659_, _28658_, _10353_);
  and (_28661_, _28659_, _10383_);
  and (_28662_, _10382_, _10349_);
  or (_28663_, _28662_, _28661_);
  and (_28664_, _28663_, _04267_);
  or (_28665_, _28630_, _25870_);
  not (_28666_, _10349_);
  nand (_28667_, _28666_, _04230_);
  or (_28668_, _04707_, \oc8051_golden_model_1.PC [8]);
  or (_28669_, _28668_, _05011_);
  and (_28670_, _28669_, _28667_);
  or (_28672_, _28670_, _04263_);
  and (_28673_, _28672_, _28665_);
  or (_28674_, _28673_, _25875_);
  or (_28675_, _28630_, _10402_);
  and (_28676_, _28675_, _04266_);
  and (_28677_, _28676_, _28674_);
  or (_28678_, _28677_, _04716_);
  or (_28679_, _28678_, _28664_);
  and (_28680_, _28679_, _28657_);
  or (_28681_, _28680_, _03850_);
  and (_28683_, _28681_, _10412_);
  and (_28684_, _28683_, _28656_);
  nor (_28685_, _28631_, _10412_);
  or (_28686_, _28685_, _03763_);
  or (_28687_, _28686_, _28684_);
  nor (_28688_, _03848_, _05045_);
  nand (_28689_, _28666_, _03763_);
  and (_28690_, _28689_, _28688_);
  and (_28691_, _28690_, _28687_);
  nand (_28692_, _10349_, _03848_);
  nand (_28694_, _28692_, _10421_);
  or (_28695_, _28694_, _28691_);
  or (_28696_, _28630_, _10421_);
  and (_28697_, _28696_, _03855_);
  and (_28698_, _28697_, _28695_);
  nand (_28699_, _10349_, _03854_);
  nand (_28700_, _28699_, _10431_);
  or (_28701_, _28700_, _28698_);
  or (_28702_, _28630_, _10431_);
  and (_28703_, _28702_, _03760_);
  and (_28705_, _28703_, _28701_);
  or (_28706_, _28705_, _28652_);
  and (_28707_, _28706_, _10256_);
  nand (_28708_, _10476_, _10189_);
  or (_28709_, _28646_, _10476_);
  and (_28710_, _28709_, _28708_);
  and (_28711_, _28710_, _04306_);
  and (_28712_, _10349_, _03758_);
  or (_28713_, _28712_, _26572_);
  or (_28714_, _28713_, _28711_);
  or (_28716_, _28714_, _28707_);
  or (_28717_, _28710_, _10441_);
  and (_28718_, _28717_, _28716_);
  or (_28719_, _28718_, _03925_);
  and (_28720_, _28719_, _28651_);
  or (_28721_, _28720_, _03868_);
  and (_28722_, _10498_, _10188_);
  nor (_28723_, _28647_, _10498_);
  or (_28724_, _28723_, _03918_);
  or (_28725_, _28724_, _28722_);
  and (_28727_, _28725_, _10486_);
  and (_28728_, _28727_, _28721_);
  and (_28729_, _28630_, _10485_);
  or (_28730_, _28646_, _10515_);
  nand (_28731_, _10515_, _10189_);
  and (_28732_, _28731_, _03920_);
  and (_28733_, _28732_, _28730_);
  or (_28734_, _28733_, _28729_);
  or (_28735_, _28734_, _28728_);
  and (_28736_, _28735_, _03753_);
  and (_28738_, _10349_, _03752_);
  or (_28739_, _28738_, _05049_);
  or (_28740_, _28739_, _28736_);
  and (_28741_, _28740_, _26231_);
  nor (_28742_, _26231_, _28666_);
  or (_28743_, _28742_, _10093_);
  or (_28744_, _28743_, _28741_);
  or (_28745_, _28630_, _10092_);
  and (_28746_, _28745_, _11731_);
  and (_28747_, _28746_, _28744_);
  and (_28749_, _10349_, _03879_);
  or (_28750_, _28749_, _25949_);
  or (_28751_, _28750_, _28747_);
  and (_28752_, _28751_, _11730_);
  nand (_28753_, _10349_, _03878_);
  nand (_28754_, _28753_, _10087_);
  or (_28755_, _28754_, _28752_);
  or (_28756_, _28630_, _10087_);
  and (_28757_, _28756_, _10085_);
  and (_28758_, _28757_, _28755_);
  nor (_28760_, _28666_, _10085_);
  or (_28761_, _28760_, _03425_);
  or (_28762_, _28761_, _28758_);
  nand (_28763_, _28631_, _03425_);
  and (_28764_, _28763_, _28762_);
  or (_28765_, _28764_, _03746_);
  nand (_28766_, _28666_, _03746_);
  nor (_28767_, _03921_, _03456_);
  and (_28768_, _28767_, _28766_);
  and (_28769_, _28768_, _28765_);
  and (_28771_, _10188_, _03921_);
  or (_28772_, _28771_, _07927_);
  nor (_28773_, _28772_, _28769_);
  nor (_28774_, _10349_, _07926_);
  nor (_28775_, _28774_, _03455_);
  not (_28776_, _28775_);
  nor (_28777_, _28776_, _28773_);
  or (_28778_, _28777_, _10558_);
  nor (_28779_, _28778_, _28643_);
  or (_28780_, _28779_, _03816_);
  nor (_28782_, _28780_, _28642_);
  nor (_28783_, _28782_, _28641_);
  nor (_28784_, _28783_, _25975_);
  and (_28785_, _28659_, _10564_);
  nor (_28786_, _28785_, _06309_);
  not (_28787_, _28786_);
  nor (_28788_, _28787_, _28784_);
  nor (_28789_, _28788_, _28640_);
  and (_28790_, _28789_, _04778_);
  and (_28791_, _10188_, _03903_);
  or (_28793_, _28791_, _28790_);
  and (_28794_, _28793_, _08493_);
  and (_28795_, _10349_, _08492_);
  nor (_28796_, _28795_, _28794_);
  nor (_28797_, _28796_, _10580_);
  and (_28798_, _10606_, _10585_);
  nor (_28799_, _28798_, _10607_);
  and (_28800_, _28799_, _10580_);
  or (_28801_, _28800_, _28797_);
  and (_28802_, _28801_, _04391_);
  and (_28804_, _10349_, _03815_);
  or (_28805_, _28804_, _03401_);
  nor (_28806_, _28805_, _28802_);
  nor (_28807_, _28806_, _10620_);
  and (_28808_, _10349_, _08826_);
  and (_28809_, _28659_, _10627_);
  or (_28810_, _28809_, _28808_);
  and (_28811_, _28810_, _10620_);
  nor (_28812_, _28811_, _10625_);
  not (_28813_, _28812_);
  nor (_28815_, _28813_, _28807_);
  or (_28816_, _28815_, _10080_);
  nor (_28817_, _28816_, _28639_);
  nor (_28818_, _28666_, _10079_);
  nor (_28819_, _28818_, _03897_);
  not (_28820_, _28819_);
  nor (_28821_, _28820_, _28817_);
  and (_28822_, _10189_, _03897_);
  nor (_28823_, _28822_, _04018_);
  not (_28824_, _28823_);
  nor (_28826_, _28824_, _28821_);
  and (_28827_, _10349_, _04018_);
  or (_28828_, _28827_, _03405_);
  nor (_28829_, _28828_, _28826_);
  nor (_28830_, _28829_, _10643_);
  nor (_28831_, _28659_, _10627_);
  nor (_28832_, _10349_, _08826_);
  nor (_28833_, _28832_, _10644_);
  not (_28834_, _28833_);
  nor (_28835_, _28834_, _28831_);
  nor (_28837_, _28835_, _10656_);
  not (_28838_, _28837_);
  nor (_28839_, _28838_, _28830_);
  nor (_28840_, _28630_, _10654_);
  nor (_28841_, _28840_, _28839_);
  nor (_28842_, _28841_, _10659_);
  nor (_28843_, _10658_, _10349_);
  nor (_28844_, _28843_, _28842_);
  and (_28845_, _28844_, _03909_);
  and (_28846_, _10188_, _03908_);
  or (_28848_, _28846_, _28845_);
  and (_28849_, _28848_, _04785_);
  and (_28850_, _10349_, _04027_);
  nor (_28851_, _28850_, _28849_);
  nor (_28852_, _28851_, _28637_);
  nor (_28853_, _28659_, \oc8051_golden_model_1.PSW [7]);
  nor (_28854_, _10349_, _08297_);
  nor (_28855_, _28854_, _10075_);
  not (_28856_, _28855_);
  nor (_28857_, _28856_, _28853_);
  nor (_28858_, _28857_, _10670_);
  not (_28859_, _28858_);
  nor (_28860_, _28859_, _28852_);
  or (_28861_, _28860_, _08582_);
  or (_28862_, _28861_, _28635_);
  nor (_28863_, _28666_, _08581_);
  nor (_28864_, _28863_, _03914_);
  and (_28865_, _28864_, _28862_);
  or (_28866_, _28865_, _28634_);
  nand (_28867_, _28866_, _06572_);
  and (_28870_, _28666_, _04011_);
  nor (_28871_, _28870_, _26033_);
  nand (_28872_, _28871_, _28867_);
  nor (_28873_, _28659_, _08297_);
  nor (_28874_, _10349_, \oc8051_golden_model_1.PSW [7]);
  nor (_28875_, _28874_, _10064_);
  not (_28876_, _28875_);
  nor (_28877_, _28876_, _28873_);
  nor (_28878_, _28877_, _10688_);
  nand (_28879_, _28878_, _28872_);
  nor (_28881_, _28630_, _10061_);
  nor (_28882_, _28881_, _08629_);
  and (_28883_, _28882_, _28879_);
  nor (_28884_, _28666_, _08628_);
  or (_28885_, _28884_, _08657_);
  or (_28886_, _28885_, _28883_);
  and (_28887_, _28631_, _08657_);
  nor (_28888_, _28887_, _04034_);
  nand (_28889_, _28888_, _28886_);
  and (_28890_, _04700_, _04034_);
  nor (_28892_, _28890_, _03383_);
  nand (_28893_, _28892_, _28889_);
  nand (_28894_, _28893_, _04097_);
  nor (_28895_, _10188_, _10906_);
  and (_28896_, _28647_, _10906_);
  or (_28897_, _28896_, _04097_);
  or (_28898_, _28897_, _28895_);
  and (_28899_, _28898_, _10059_);
  nand (_28900_, _28899_, _28894_);
  nor (_28901_, _28630_, _10059_);
  nor (_28903_, _28901_, _10057_);
  nand (_28904_, _28903_, _28900_);
  nor (_28905_, _28666_, _10056_);
  nor (_28906_, _28905_, _08772_);
  and (_28907_, _28906_, _28904_);
  or (_28908_, _28907_, _28633_);
  and (_28909_, _04700_, _03777_);
  nor (_28910_, _28909_, _03410_);
  nand (_28911_, _28910_, _28908_);
  nand (_28912_, _28911_, _03776_);
  and (_28914_, _10189_, _10906_);
  nor (_28915_, _28646_, _10906_);
  nor (_28916_, _28915_, _28914_);
  and (_28917_, _28916_, _03775_);
  nor (_28918_, _28917_, _10937_);
  nand (_28919_, _28918_, _28912_);
  nor (_28920_, _28630_, _10936_);
  nor (_28921_, _28920_, _03773_);
  nand (_28922_, _28921_, _28919_);
  and (_28923_, _10349_, _03773_);
  nor (_28925_, _28923_, _26446_);
  nand (_28926_, _28925_, _28922_);
  nor (_28927_, _28630_, _10943_);
  nor (_28928_, _28927_, _03899_);
  and (_28929_, _28928_, _28926_);
  or (_28930_, _28929_, _28628_);
  nor (_28931_, _03414_, _03374_);
  nand (_28932_, _28931_, _28930_);
  and (_28933_, _28916_, _03374_);
  nor (_28934_, _28933_, _10959_);
  nand (_28936_, _28934_, _28932_);
  nor (_28937_, _28630_, _10958_);
  nor (_28938_, _28937_, _03772_);
  nand (_28939_, _28938_, _28936_);
  and (_28940_, _10349_, _03772_);
  nor (_28941_, _28940_, _28254_);
  nand (_28942_, _28941_, _28939_);
  nor (_28943_, _28630_, _10965_);
  nor (_28944_, _28943_, _03901_);
  and (_28945_, _28944_, _28942_);
  or (_28947_, _28945_, _28626_);
  nor (_28948_, _10042_, _03413_);
  and (_28949_, _28948_, _28947_);
  and (_28950_, _28630_, _10042_);
  or (_28951_, _28950_, _28949_);
  or (_28952_, _28951_, _43156_);
  or (_28953_, _43152_, \oc8051_golden_model_1.PC [8]);
  and (_28954_, _28953_, _41894_);
  and (_43517_, _28954_, _28952_);
  nor (_28955_, _04563_, _10969_);
  nor (_28957_, _04563_, _03900_);
  nor (_28958_, _10045_, \oc8051_golden_model_1.PC [9]);
  nor (_28959_, _28958_, _10046_);
  nor (_28960_, _28959_, _10059_);
  nor (_28961_, _28959_, _10061_);
  and (_28962_, _10128_, _03914_);
  nor (_28963_, _28959_, _10072_);
  and (_28964_, _10128_, _03908_);
  nor (_28965_, _28959_, _10654_);
  and (_28966_, _10128_, _03897_);
  nor (_28968_, _28959_, _10082_);
  and (_28969_, _10297_, _03816_);
  nor (_28970_, _28959_, _10556_);
  nor (_28971_, _10297_, _10085_);
  nor (_28972_, _03878_, _25949_);
  not (_28973_, _28972_);
  nor (_28974_, _28959_, _10092_);
  nor (_28975_, _10193_, _10190_);
  and (_28976_, _28975_, _10132_);
  nor (_28977_, _28975_, _10132_);
  nor (_28979_, _28977_, _28976_);
  nor (_28980_, _28979_, _25901_);
  and (_28981_, _25901_, _10128_);
  or (_28982_, _28981_, _04722_);
  or (_28983_, _28982_, _28980_);
  nor (_28984_, _10353_, _10350_);
  and (_28985_, _28984_, _10300_);
  nor (_28986_, _28984_, _10300_);
  nor (_28987_, _28986_, _28985_);
  nor (_28988_, _28987_, _10382_);
  and (_28990_, _25887_, _10297_);
  or (_28991_, _28990_, _28988_);
  or (_28992_, _28991_, _04266_);
  and (_28993_, _10402_, _05012_);
  or (_28994_, _28993_, _28959_);
  not (_28995_, _10297_);
  nand (_28996_, _28995_, _04707_);
  and (_28997_, _28996_, _26504_);
  or (_28998_, _04707_, \oc8051_golden_model_1.PC [9]);
  or (_28999_, _28998_, _05011_);
  and (_29001_, _28999_, _28997_);
  or (_29002_, _29001_, _25875_);
  and (_29003_, _29002_, _28994_);
  nand (_29004_, _28959_, _04263_);
  nand (_29005_, _29004_, _04266_);
  or (_29006_, _29005_, _29003_);
  and (_29007_, _29006_, _04717_);
  and (_29008_, _29007_, _28992_);
  and (_29009_, _28959_, _04716_);
  or (_29010_, _29009_, _03850_);
  or (_29012_, _29010_, _29008_);
  and (_29013_, _29012_, _28983_);
  or (_29014_, _29013_, _10413_);
  or (_29015_, _28959_, _10412_);
  and (_29016_, _29015_, _03764_);
  and (_29017_, _29016_, _29014_);
  and (_29018_, _10297_, _03763_);
  or (_29019_, _29018_, _05045_);
  or (_29020_, _29019_, _29017_);
  and (_29021_, _29020_, _04733_);
  nand (_29023_, _10297_, _03848_);
  nand (_29024_, _29023_, _10421_);
  or (_29025_, _29024_, _29021_);
  or (_29026_, _28959_, _10421_);
  and (_29027_, _29026_, _03855_);
  and (_29028_, _29027_, _29025_);
  nand (_29029_, _10297_, _03854_);
  nand (_29030_, _29029_, _10431_);
  or (_29031_, _29030_, _29028_);
  or (_29032_, _28959_, _10431_);
  and (_29034_, _29032_, _03760_);
  and (_29035_, _29034_, _29031_);
  and (_29036_, _10297_, _03759_);
  or (_29037_, _29036_, _10255_);
  or (_29038_, _29037_, _29035_);
  and (_29039_, _29038_, _04845_);
  nand (_29040_, _10297_, _03758_);
  nand (_29041_, _29040_, _10441_);
  or (_29042_, _29041_, _29039_);
  nor (_29043_, _28979_, _10476_);
  and (_29045_, _10476_, _10128_);
  or (_29046_, _29045_, _10441_);
  or (_29047_, _29046_, _29043_);
  and (_29048_, _29047_, _29042_);
  or (_29049_, _29048_, _03925_);
  nand (_29050_, _10249_, _10129_);
  not (_29051_, _28979_);
  or (_29052_, _29051_, _10249_);
  and (_29053_, _29052_, _29050_);
  or (_29054_, _29053_, _10444_);
  and (_29056_, _29054_, _29049_);
  or (_29057_, _29056_, _03868_);
  and (_29058_, _10498_, _10128_);
  nor (_29059_, _28979_, _10498_);
  or (_29060_, _29059_, _03918_);
  or (_29061_, _29060_, _29058_);
  and (_29062_, _29061_, _10486_);
  and (_29063_, _29062_, _29057_);
  and (_29064_, _10515_, _10128_);
  nor (_29065_, _28979_, _10515_);
  or (_29067_, _29065_, _29064_);
  and (_29068_, _29067_, _03920_);
  and (_29069_, _28959_, _10485_);
  nor (_29070_, _29069_, _29068_);
  and (_29071_, _29070_, _03753_);
  not (_29072_, _29071_);
  nor (_29073_, _29072_, _29063_);
  and (_29074_, _28995_, _03752_);
  nor (_29075_, _29074_, _05049_);
  nand (_29076_, _29075_, _26231_);
  nor (_29078_, _29076_, _29073_);
  nor (_29079_, _26231_, _28995_);
  nor (_29080_, _29079_, _10093_);
  not (_29081_, _29080_);
  nor (_29082_, _29081_, _29078_);
  or (_29083_, _29082_, _03879_);
  nor (_29084_, _29083_, _28974_);
  and (_29085_, _10297_, _03879_);
  nor (_29086_, _29085_, _29084_);
  nor (_29087_, _29086_, _28973_);
  and (_29089_, _10297_, _03878_);
  nor (_29090_, _29089_, _15018_);
  not (_29091_, _29090_);
  nor (_29092_, _29091_, _29087_);
  nor (_29093_, _28959_, _10087_);
  nor (_29094_, _29093_, _29092_);
  nor (_29095_, _29094_, _10086_);
  or (_29096_, _29095_, _03425_);
  nor (_29097_, _29096_, _28971_);
  and (_29098_, _28959_, _03425_);
  or (_29100_, _29098_, _29097_);
  and (_29101_, _29100_, _03747_);
  and (_29102_, _10297_, _03746_);
  or (_29103_, _29102_, _29101_);
  and (_29104_, _29103_, _06141_);
  and (_29105_, _29104_, _09861_);
  and (_29106_, _10128_, _03921_);
  nor (_29107_, _29106_, _07927_);
  not (_29108_, _29107_);
  nor (_29109_, _29108_, _29105_);
  nor (_29111_, _10297_, _07926_);
  nor (_29112_, _29111_, _03455_);
  not (_29113_, _29112_);
  nor (_29114_, _29113_, _29109_);
  and (_29115_, _10128_, _03455_);
  nor (_29116_, _29115_, _10558_);
  not (_29117_, _29116_);
  nor (_29118_, _29117_, _29114_);
  or (_29119_, _29118_, _03816_);
  nor (_29120_, _29119_, _28970_);
  nor (_29122_, _29120_, _28969_);
  nor (_29123_, _29122_, _25975_);
  nor (_29124_, _28987_, _10565_);
  nor (_29125_, _29124_, _06309_);
  not (_29126_, _29125_);
  nor (_29127_, _29126_, _29123_);
  nor (_29128_, _10297_, _06138_);
  nor (_29129_, _29128_, _03903_);
  not (_29130_, _29129_);
  nor (_29131_, _29130_, _29127_);
  and (_29133_, _10128_, _03903_);
  or (_29134_, _29133_, _29131_);
  and (_29135_, _29134_, _08493_);
  and (_29136_, _10297_, _08492_);
  or (_29137_, _29136_, _29135_);
  and (_29138_, _29137_, _10581_);
  nor (_29139_, _10607_, \oc8051_golden_model_1.DPH [1]);
  not (_29140_, _29139_);
  nor (_29141_, _10608_, _10581_);
  and (_29142_, _29141_, _29140_);
  nor (_29144_, _29142_, _29138_);
  nor (_29145_, _29144_, _03815_);
  and (_29146_, _10297_, _03815_);
  or (_29147_, _29146_, _03401_);
  nor (_29148_, _29147_, _29145_);
  nor (_29149_, _29148_, _10620_);
  and (_29150_, _10297_, _08826_);
  nor (_29151_, _28987_, _08826_);
  or (_29152_, _29151_, _29150_);
  and (_29153_, _29152_, _10620_);
  nor (_29155_, _29153_, _10625_);
  not (_29156_, _29155_);
  nor (_29157_, _29156_, _29149_);
  nor (_29158_, _29157_, _28968_);
  nor (_29159_, _29158_, _10080_);
  nor (_29160_, _10297_, _10079_);
  nor (_29161_, _29160_, _03897_);
  not (_29162_, _29161_);
  nor (_29163_, _29162_, _29159_);
  nor (_29164_, _29163_, _28966_);
  nor (_29166_, _29164_, _04018_);
  and (_29167_, _10297_, _04018_);
  nor (_29168_, _29167_, _29166_);
  and (_29169_, _29168_, _25850_);
  or (_29170_, _29169_, _10643_);
  and (_29171_, _28987_, _08826_);
  nor (_29172_, _10297_, _08826_);
  nor (_29173_, _29172_, _10644_);
  not (_29174_, _29173_);
  nor (_29175_, _29174_, _29171_);
  nor (_29177_, _29175_, _10656_);
  and (_29178_, _29177_, _29170_);
  or (_29179_, _29178_, _28965_);
  and (_29180_, _29179_, _10658_);
  nor (_29181_, _10658_, _10297_);
  nor (_29182_, _29181_, _03908_);
  not (_29183_, _29182_);
  nor (_29184_, _29183_, _29180_);
  or (_29185_, _29184_, _28964_);
  nand (_29186_, _29185_, _04785_);
  and (_29188_, _10297_, _04027_);
  nor (_29189_, _29188_, _03388_);
  nand (_29190_, _29189_, _29186_);
  nand (_29191_, _29190_, _10075_);
  and (_29192_, _28987_, _08297_);
  nor (_29193_, _10297_, _08297_);
  nor (_29194_, _29193_, _10075_);
  not (_29195_, _29194_);
  nor (_29196_, _29195_, _29192_);
  nor (_29197_, _29196_, _10670_);
  and (_29199_, _29197_, _29191_);
  or (_29200_, _29199_, _28963_);
  nand (_29201_, _29200_, _08581_);
  nor (_29202_, _10297_, _08581_);
  nor (_29203_, _29202_, _03914_);
  and (_29204_, _29203_, _29201_);
  or (_29205_, _29204_, _28962_);
  nand (_29206_, _29205_, _06572_);
  and (_29207_, _10297_, _04011_);
  nor (_29208_, _29207_, _03393_);
  nand (_29210_, _29208_, _29206_);
  nand (_29211_, _29210_, _10064_);
  and (_29212_, _28987_, \oc8051_golden_model_1.PSW [7]);
  nor (_29213_, _10297_, \oc8051_golden_model_1.PSW [7]);
  nor (_29214_, _29213_, _10064_);
  not (_29215_, _29214_);
  nor (_29216_, _29215_, _29212_);
  nor (_29217_, _29216_, _10688_);
  and (_29218_, _29217_, _29211_);
  or (_29219_, _29218_, _28961_);
  nand (_29221_, _29219_, _08628_);
  nor (_29222_, _10297_, _08628_);
  nor (_29223_, _29222_, _08657_);
  nand (_29224_, _29223_, _29221_);
  and (_29225_, _28959_, _08657_);
  nor (_29226_, _29225_, _04034_);
  nand (_29227_, _29226_, _29224_);
  nor (_29228_, _03913_, _03383_);
  not (_29229_, _29228_);
  nor (_29230_, _04900_, _10704_);
  nor (_29232_, _29230_, _29229_);
  nand (_29233_, _29232_, _29227_);
  nor (_29234_, _10128_, _10906_);
  and (_29235_, _28979_, _10906_);
  or (_29236_, _29235_, _04097_);
  or (_29237_, _29236_, _29234_);
  and (_29238_, _29237_, _10059_);
  and (_29239_, _29238_, _29233_);
  or (_29240_, _29239_, _28960_);
  nand (_29241_, _29240_, _10056_);
  nor (_29243_, _10297_, _10056_);
  nor (_29244_, _29243_, _08772_);
  nand (_29245_, _29244_, _29241_);
  and (_29246_, _28959_, _08772_);
  nor (_29247_, _29246_, _03777_);
  nand (_29248_, _29247_, _29245_);
  nor (_29249_, _03775_, _03410_);
  not (_29250_, _29249_);
  nor (_29251_, _04900_, _03778_);
  nor (_29252_, _29251_, _29250_);
  nand (_29254_, _29252_, _29248_);
  and (_29255_, _10129_, _10906_);
  nor (_29256_, _29051_, _10906_);
  nor (_29257_, _29256_, _29255_);
  and (_29258_, _29257_, _03775_);
  nor (_29259_, _29258_, _10937_);
  nand (_29260_, _29259_, _29254_);
  nor (_29261_, _28959_, _10936_);
  nor (_29262_, _29261_, _03773_);
  nand (_29263_, _29262_, _29260_);
  and (_29265_, _10297_, _03773_);
  nor (_29266_, _29265_, _26446_);
  nand (_29267_, _29266_, _29263_);
  nor (_29268_, _28959_, _10943_);
  nor (_29269_, _29268_, _03899_);
  and (_29270_, _29269_, _29267_);
  or (_29271_, _29270_, _28957_);
  nand (_29272_, _29271_, _28931_);
  and (_29273_, _29257_, _03374_);
  nor (_29274_, _29273_, _10959_);
  nand (_29276_, _29274_, _29272_);
  nor (_29277_, _28959_, _10958_);
  nor (_29278_, _29277_, _03772_);
  nand (_29279_, _29278_, _29276_);
  and (_29280_, _10297_, _03772_);
  nor (_29281_, _29280_, _28254_);
  nand (_29282_, _29281_, _29279_);
  nor (_29283_, _28959_, _10965_);
  nor (_29284_, _29283_, _03901_);
  and (_29285_, _29284_, _29282_);
  or (_29286_, _29285_, _28955_);
  and (_29287_, _29286_, _28948_);
  and (_29288_, _28959_, _10042_);
  or (_29289_, _29288_, _29287_);
  or (_29290_, _29289_, _43156_);
  or (_29291_, _43152_, \oc8051_golden_model_1.PC [9]);
  and (_29292_, _29291_, _41894_);
  and (_43518_, _29292_, _29290_);
  nor (_29293_, _10046_, \oc8051_golden_model_1.PC [10]);
  nor (_29294_, _29293_, _10047_);
  or (_29296_, _29294_, _10936_);
  or (_29297_, _29294_, _08773_);
  or (_29298_, _29294_, _08658_);
  nand (_29299_, _10115_, _03914_);
  nand (_29300_, _10115_, _03908_);
  nand (_29301_, _10115_, _03897_);
  nor (_29302_, _10620_, _03401_);
  and (_29303_, _29294_, _10558_);
  and (_29304_, _29294_, _15018_);
  nand (_29305_, _10249_, _10115_);
  nor (_29307_, _10197_, _10194_);
  not (_29308_, _29307_);
  and (_29309_, _29308_, _10125_);
  nor (_29310_, _29308_, _10125_);
  nor (_29311_, _29310_, _29309_);
  or (_29312_, _29311_, _10249_);
  and (_29313_, _29312_, _03925_);
  and (_29314_, _29313_, _29305_);
  or (_29315_, _29294_, _10421_);
  and (_29316_, _25870_, _10402_);
  or (_29318_, _29316_, _29294_);
  not (_29319_, _10291_);
  nand (_29320_, _29319_, _04230_);
  or (_29321_, _04707_, \oc8051_golden_model_1.PC [10]);
  or (_29322_, _29321_, _05011_);
  and (_29323_, _29322_, _29320_);
  or (_29324_, _29323_, _04263_);
  and (_29325_, _29324_, _29318_);
  and (_29326_, _29294_, _26516_);
  nand (_29327_, _04266_, _03770_);
  or (_29329_, _29327_, _29326_);
  or (_29330_, _29329_, _29325_);
  nor (_29331_, _10357_, _10354_);
  not (_29332_, _29331_);
  and (_29333_, _29332_, _10294_);
  nor (_29334_, _29332_, _10294_);
  nor (_29335_, _29334_, _29333_);
  and (_29336_, _29335_, _10383_);
  and (_29337_, _10382_, _10291_);
  or (_29338_, _29337_, _29336_);
  or (_29340_, _29338_, _04266_);
  and (_29341_, _29340_, _29330_);
  or (_29342_, _29341_, _04716_);
  or (_29343_, _29294_, _04717_);
  and (_29344_, _29343_, _04722_);
  and (_29345_, _29344_, _29342_);
  or (_29346_, _29311_, _10265_);
  nand (_29347_, _25901_, _10115_);
  and (_29348_, _29347_, _29346_);
  and (_29349_, _29348_, _03850_);
  or (_29351_, _29349_, _29345_);
  or (_29352_, _29351_, _10413_);
  or (_29353_, _29294_, _10412_);
  and (_29354_, _29353_, _03764_);
  and (_29355_, _29354_, _29352_);
  or (_29356_, _29355_, _05045_);
  and (_29357_, _29356_, _04733_);
  or (_29358_, _29319_, _03856_);
  nand (_29359_, _29358_, _10421_);
  or (_29360_, _29359_, _29357_);
  and (_29362_, _29360_, _29315_);
  or (_29363_, _29362_, _03854_);
  nand (_29364_, _29319_, _03854_);
  and (_29365_, _29364_, _10431_);
  and (_29366_, _29365_, _29363_);
  and (_29367_, _29294_, _10434_);
  or (_29368_, _29367_, _29366_);
  and (_29369_, _29368_, _03760_);
  and (_29370_, _10291_, _03759_);
  or (_29371_, _29370_, _10255_);
  or (_29373_, _29371_, _29369_);
  and (_29374_, _29373_, _04845_);
  nand (_29375_, _10476_, _10115_);
  or (_29376_, _29311_, _10476_);
  and (_29377_, _29376_, _29375_);
  and (_29378_, _29377_, _04306_);
  and (_29379_, _10291_, _03758_);
  or (_29380_, _29379_, _26572_);
  or (_29381_, _29380_, _29378_);
  or (_29382_, _29381_, _29374_);
  or (_29384_, _29377_, _10441_);
  and (_29385_, _29384_, _10444_);
  and (_29386_, _29385_, _29382_);
  or (_29387_, _29386_, _29314_);
  and (_29388_, _29387_, _03918_);
  and (_29389_, _29311_, _10500_);
  and (_29390_, _10498_, _10114_);
  or (_29391_, _29390_, _29389_);
  and (_29392_, _29391_, _03868_);
  or (_29393_, _29392_, _29388_);
  and (_29395_, _29393_, _10486_);
  and (_29396_, _29294_, _10485_);
  or (_29397_, _29311_, _10515_);
  nand (_29398_, _10515_, _10115_);
  and (_29399_, _29398_, _03920_);
  and (_29400_, _29399_, _29397_);
  or (_29401_, _29400_, _29396_);
  or (_29402_, _29401_, _29395_);
  and (_29403_, _26231_, _03753_);
  and (_29404_, _29403_, _29402_);
  nor (_29405_, _29403_, _29319_);
  nand (_29406_, _10092_, _03428_);
  or (_29407_, _29406_, _29405_);
  or (_29408_, _29407_, _29404_);
  or (_29409_, _29294_, _10092_);
  and (_29410_, _29409_, _11731_);
  and (_29411_, _29410_, _29408_);
  nand (_29412_, _10291_, _03879_);
  nand (_29413_, _29412_, _28972_);
  or (_29414_, _29413_, _29411_);
  nand (_29417_, _29319_, _03878_);
  and (_29418_, _29417_, _10087_);
  and (_29419_, _29418_, _29414_);
  or (_29420_, _29419_, _29304_);
  and (_29421_, _29420_, _10085_);
  nor (_29422_, _29319_, _10085_);
  or (_29423_, _29422_, _03425_);
  or (_29424_, _29423_, _29421_);
  or (_29425_, _29294_, _03426_);
  and (_29426_, _29425_, _03747_);
  and (_29428_, _29426_, _29424_);
  nand (_29429_, _10291_, _03746_);
  nand (_29430_, _29429_, _28767_);
  or (_29431_, _29430_, _29428_);
  nand (_29432_, _10115_, _03921_);
  and (_29433_, _29432_, _07926_);
  and (_29434_, _29433_, _29431_);
  nor (_29435_, _29319_, _07926_);
  or (_29436_, _29435_, _03455_);
  or (_29437_, _29436_, _29434_);
  nand (_29439_, _10115_, _03455_);
  and (_29440_, _29439_, _10556_);
  and (_29441_, _29440_, _29437_);
  or (_29442_, _29441_, _29303_);
  and (_29443_, _29442_, _27373_);
  nand (_29444_, _10291_, _03816_);
  nand (_29445_, _29444_, _25974_);
  or (_29446_, _29445_, _29443_);
  or (_29447_, _29335_, _10565_);
  and (_29448_, _29447_, _06138_);
  and (_29450_, _29448_, _29446_);
  nor (_29451_, _29319_, _06138_);
  or (_29452_, _29451_, _03903_);
  or (_29453_, _29452_, _29450_);
  nand (_29454_, _10115_, _03903_);
  and (_29455_, _29454_, _08493_);
  and (_29456_, _29455_, _29453_);
  and (_29457_, _10291_, _08492_);
  or (_29458_, _29457_, _10580_);
  or (_29459_, _29458_, _29456_);
  nor (_29461_, _10608_, \oc8051_golden_model_1.DPH [2]);
  nor (_29462_, _29461_, _10609_);
  or (_29463_, _29462_, _10581_);
  and (_29464_, _29463_, _04391_);
  and (_29465_, _29464_, _29459_);
  and (_29466_, _10291_, _03815_);
  or (_29467_, _29466_, _29465_);
  and (_29468_, _29467_, _29302_);
  or (_29469_, _29335_, _08826_);
  or (_29470_, _10291_, _10627_);
  and (_29472_, _29470_, _10620_);
  and (_29473_, _29472_, _29469_);
  or (_29474_, _29473_, _10625_);
  or (_29475_, _29474_, _29468_);
  or (_29476_, _29294_, _10082_);
  and (_29477_, _29476_, _10079_);
  and (_29478_, _29477_, _29475_);
  nor (_29479_, _29319_, _10079_);
  or (_29480_, _29479_, _03897_);
  or (_29481_, _29480_, _29478_);
  and (_29483_, _29481_, _29301_);
  or (_29484_, _29483_, _04018_);
  nand (_29485_, _29319_, _04018_);
  nor (_29486_, _10643_, _03405_);
  and (_29487_, _29486_, _29485_);
  and (_29488_, _29487_, _29484_);
  or (_29489_, _29335_, _10627_);
  or (_29490_, _10291_, _08826_);
  and (_29491_, _29490_, _10643_);
  and (_29492_, _29491_, _29489_);
  or (_29494_, _29492_, _10656_);
  or (_29495_, _29494_, _29488_);
  or (_29496_, _29294_, _10654_);
  and (_29497_, _29496_, _10658_);
  and (_29498_, _29497_, _29495_);
  nor (_29499_, _10658_, _29319_);
  or (_29500_, _29499_, _03908_);
  or (_29501_, _29500_, _29498_);
  and (_29502_, _29501_, _29300_);
  or (_29503_, _29502_, _04027_);
  nand (_29505_, _29319_, _04027_);
  and (_29506_, _29505_, _28636_);
  and (_29507_, _29506_, _29503_);
  or (_29508_, _29335_, \oc8051_golden_model_1.PSW [7]);
  or (_29509_, _10291_, _08297_);
  and (_29510_, _29509_, _10074_);
  and (_29511_, _29510_, _29508_);
  or (_29512_, _29511_, _10670_);
  or (_29513_, _29512_, _29507_);
  or (_29514_, _29294_, _10072_);
  and (_29516_, _29514_, _08581_);
  and (_29517_, _29516_, _29513_);
  nor (_29518_, _29319_, _08581_);
  or (_29519_, _29518_, _03914_);
  or (_29520_, _29519_, _29517_);
  and (_29521_, _29520_, _29299_);
  or (_29522_, _29521_, _04011_);
  nand (_29523_, _29319_, _04011_);
  and (_29524_, _29523_, _26032_);
  and (_29525_, _29524_, _29522_);
  or (_29527_, _29335_, _08297_);
  or (_29528_, _10291_, \oc8051_golden_model_1.PSW [7]);
  and (_29529_, _29528_, _10063_);
  and (_29530_, _29529_, _29527_);
  or (_29531_, _29530_, _10688_);
  or (_29532_, _29531_, _29525_);
  or (_29533_, _29294_, _10061_);
  and (_29534_, _29533_, _08628_);
  and (_29535_, _29534_, _29532_);
  nor (_29536_, _29319_, _08628_);
  or (_29538_, _29536_, _08657_);
  or (_29539_, _29538_, _29535_);
  and (_29540_, _29539_, _29298_);
  or (_29541_, _29540_, _04034_);
  or (_29542_, _05307_, _10704_);
  and (_29543_, _29542_, _29228_);
  and (_29544_, _29543_, _29541_);
  or (_29545_, _29311_, _10907_);
  or (_29546_, _10114_, _10906_);
  and (_29547_, _29546_, _03913_);
  and (_29549_, _29547_, _29545_);
  or (_29550_, _29549_, _10712_);
  or (_29551_, _29550_, _29544_);
  or (_29552_, _29294_, _10059_);
  and (_29553_, _29552_, _10056_);
  and (_29554_, _29553_, _29551_);
  nor (_29555_, _29319_, _10056_);
  or (_29556_, _29555_, _08772_);
  or (_29557_, _29556_, _29554_);
  and (_29558_, _29557_, _29297_);
  or (_29560_, _29558_, _03777_);
  or (_29561_, _05307_, _03778_);
  and (_29562_, _29561_, _29249_);
  and (_29563_, _29562_, _29560_);
  nand (_29564_, _10115_, _10906_);
  or (_29565_, _29311_, _10906_);
  and (_29566_, _29565_, _29564_);
  and (_29567_, _29566_, _03775_);
  or (_29568_, _29567_, _10937_);
  or (_29569_, _29568_, _29563_);
  and (_29571_, _29569_, _29296_);
  or (_29572_, _29571_, _03773_);
  nand (_29573_, _29319_, _03773_);
  and (_29574_, _29573_, _10943_);
  and (_29575_, _29574_, _29572_);
  and (_29576_, _29294_, _26446_);
  or (_29577_, _29576_, _03899_);
  or (_29578_, _29577_, _29575_);
  nand (_29579_, _04139_, _03899_);
  and (_29580_, _29579_, _28931_);
  and (_29582_, _29580_, _29578_);
  and (_29583_, _29566_, _03374_);
  or (_29584_, _29583_, _10959_);
  or (_29585_, _29584_, _29582_);
  or (_29586_, _29294_, _10958_);
  and (_29587_, _29586_, _29585_);
  or (_29588_, _29587_, _03772_);
  nand (_29589_, _29319_, _03772_);
  and (_29590_, _29589_, _10965_);
  and (_29591_, _29590_, _29588_);
  and (_29593_, _29294_, _28254_);
  or (_29594_, _29593_, _03901_);
  or (_29595_, _29594_, _29591_);
  nand (_29596_, _04139_, _03901_);
  and (_29597_, _29596_, _28948_);
  and (_29598_, _29597_, _29595_);
  and (_29599_, _29294_, _10042_);
  or (_29600_, _29599_, _29598_);
  or (_29601_, _29600_, _43156_);
  or (_29602_, _43152_, \oc8051_golden_model_1.PC [10]);
  and (_29604_, _29602_, _41894_);
  and (_43519_, _29604_, _29601_);
  nor (_29605_, _10047_, \oc8051_golden_model_1.PC [11]);
  nor (_29606_, _29605_, _10048_);
  not (_29607_, _29606_);
  and (_29608_, _29607_, _10042_);
  nor (_29609_, _29606_, _10059_);
  nor (_29610_, _29606_, _10061_);
  nor (_29611_, _10286_, _10065_);
  or (_29612_, _29611_, _10063_);
  nor (_29614_, _29606_, _10072_);
  nor (_29615_, _29606_, _10082_);
  nor (_29616_, _10560_, _10286_);
  and (_29617_, _10119_, _03455_);
  and (_29618_, _10286_, _03854_);
  nor (_29619_, _29607_, _10417_);
  and (_29620_, _25906_, _10119_);
  nor (_29621_, _29309_, _10116_);
  and (_29622_, _29621_, _10123_);
  nor (_29623_, _29621_, _10123_);
  nor (_29625_, _29623_, _29622_);
  nor (_29626_, _29625_, _25906_);
  or (_29627_, _29626_, _29620_);
  and (_29628_, _29627_, _03850_);
  nor (_29629_, _29333_, _10292_);
  and (_29630_, _29629_, _10289_);
  nor (_29631_, _29629_, _10289_);
  nor (_29632_, _29631_, _29630_);
  nor (_29633_, _29632_, _10382_);
  and (_29634_, _25887_, _10286_);
  or (_29636_, _29634_, _29633_);
  or (_29637_, _29636_, _04266_);
  or (_29638_, _29606_, _29316_);
  not (_29639_, _10286_);
  nand (_29640_, _29639_, _04230_);
  or (_29641_, _04707_, \oc8051_golden_model_1.PC [11]);
  or (_29642_, _29641_, _05011_);
  and (_29643_, _29642_, _29640_);
  or (_29644_, _29643_, _04263_);
  and (_29645_, _29644_, _03770_);
  and (_29647_, _29645_, _29638_);
  and (_29648_, _10286_, _03768_);
  nor (_29649_, _29607_, _10402_);
  or (_29650_, _29649_, _04267_);
  or (_29651_, _29650_, _29648_);
  or (_29652_, _29651_, _29647_);
  and (_29653_, _29652_, _26151_);
  and (_29654_, _29653_, _29637_);
  or (_29655_, _29654_, _29628_);
  and (_29656_, _29655_, _10412_);
  or (_29658_, _29656_, _29619_);
  and (_29659_, _29658_, _10416_);
  or (_29660_, _10416_, _29639_);
  nand (_29661_, _29660_, _10421_);
  or (_29662_, _29661_, _29659_);
  or (_29663_, _29606_, _10421_);
  and (_29664_, _29663_, _03855_);
  and (_29665_, _29664_, _29662_);
  or (_29666_, _29665_, _29618_);
  and (_29667_, _29666_, _10431_);
  or (_29668_, _29607_, _10431_);
  nand (_29669_, _29668_, _10257_);
  or (_29670_, _29669_, _29667_);
  or (_29671_, _10257_, _10286_);
  and (_29672_, _29671_, _10441_);
  and (_29673_, _29672_, _29670_);
  nand (_29674_, _10476_, _10120_);
  not (_29675_, _29625_);
  or (_29676_, _29675_, _10476_);
  and (_29677_, _29676_, _10442_);
  and (_29680_, _29677_, _29674_);
  or (_29681_, _29680_, _03925_);
  or (_29682_, _29681_, _29673_);
  and (_29683_, _10249_, _10119_);
  nor (_29684_, _29625_, _10249_);
  or (_29685_, _29684_, _29683_);
  or (_29686_, _29685_, _10444_);
  and (_29687_, _29686_, _29682_);
  nor (_29688_, _29687_, _03868_);
  and (_29689_, _10498_, _10119_);
  nor (_29691_, _29625_, _10498_);
  or (_29692_, _29691_, _03918_);
  nor (_29693_, _29692_, _29689_);
  or (_29694_, _29693_, _27224_);
  or (_29695_, _29694_, _29688_);
  not (_29696_, _10515_);
  and (_29697_, _29625_, _29696_);
  and (_29698_, _10515_, _10120_);
  or (_29699_, _29698_, _11857_);
  or (_29700_, _29699_, _29697_);
  nand (_29702_, _29606_, _10485_);
  and (_29703_, _29702_, _10523_);
  and (_29704_, _29703_, _29700_);
  and (_29705_, _29704_, _29695_);
  nor (_29706_, _10523_, _10286_);
  or (_29707_, _29706_, _10093_);
  or (_29708_, _29707_, _29705_);
  or (_29709_, _29607_, _10092_);
  and (_29710_, _29709_, _10531_);
  nand (_29711_, _29710_, _29708_);
  or (_29713_, _10531_, _10286_);
  and (_29714_, _29713_, _10087_);
  and (_29715_, _29714_, _29711_);
  nor (_29716_, _29607_, _10087_);
  nor (_29717_, _29716_, _10086_);
  not (_29718_, _29717_);
  nor (_29719_, _29718_, _29715_);
  nor (_29720_, _10286_, _10085_);
  nor (_29721_, _29720_, _03425_);
  not (_29722_, _29721_);
  nor (_29724_, _29722_, _29719_);
  and (_29725_, _29606_, _03425_);
  nor (_29726_, _29725_, _10543_);
  not (_29727_, _29726_);
  nor (_29728_, _29727_, _29724_);
  nor (_29729_, _10542_, _10286_);
  nor (_29730_, _29729_, _03921_);
  not (_29731_, _29730_);
  nor (_29732_, _29731_, _29728_);
  and (_29733_, _10119_, _03921_);
  nor (_29735_, _29733_, _07927_);
  not (_29736_, _29735_);
  nor (_29737_, _29736_, _29732_);
  nor (_29738_, _10286_, _07926_);
  nor (_29739_, _29738_, _03455_);
  not (_29740_, _29739_);
  nor (_29741_, _29740_, _29737_);
  nor (_29742_, _29741_, _29617_);
  nor (_29743_, _29742_, _10558_);
  nor (_29744_, _29607_, _10556_);
  nor (_29746_, _29744_, _10561_);
  not (_29747_, _29746_);
  nor (_29748_, _29747_, _29743_);
  or (_29749_, _29748_, _10564_);
  nor (_29750_, _29749_, _29616_);
  nor (_29751_, _29632_, _10565_);
  nor (_29752_, _29751_, _06309_);
  not (_29753_, _29752_);
  nor (_29754_, _29753_, _29750_);
  nor (_29755_, _29639_, _03903_);
  nor (_29757_, _29755_, _06139_);
  nor (_29758_, _29757_, _29754_);
  and (_29759_, _10119_, _03903_);
  or (_29760_, _29759_, _29758_);
  and (_29761_, _29760_, _08493_);
  and (_29762_, _10286_, _08492_);
  or (_29763_, _29762_, _29761_);
  and (_29764_, _29763_, _10581_);
  nor (_29765_, _10609_, \oc8051_golden_model_1.DPH [3]);
  or (_29766_, _29765_, _10581_);
  or (_29768_, _29766_, _10610_);
  and (_29769_, _29768_, _10583_);
  not (_29770_, _29769_);
  nor (_29771_, _29770_, _29764_);
  nor (_29772_, _10583_, _10286_);
  nor (_29773_, _29772_, _10620_);
  not (_29774_, _29773_);
  nor (_29775_, _29774_, _29771_);
  and (_29776_, _10286_, _08826_);
  nor (_29777_, _29632_, _08826_);
  or (_29779_, _29777_, _29776_);
  and (_29780_, _29779_, _10620_);
  nor (_29781_, _29780_, _10625_);
  not (_29782_, _29781_);
  nor (_29783_, _29782_, _29775_);
  nor (_29784_, _29783_, _29615_);
  nor (_29785_, _29784_, _10080_);
  nor (_29786_, _10286_, _10079_);
  nor (_29787_, _29786_, _03897_);
  not (_29788_, _29787_);
  nor (_29790_, _29788_, _29785_);
  not (_29791_, _10639_);
  and (_29792_, _10119_, _03897_);
  nor (_29793_, _29792_, _29791_);
  not (_29794_, _29793_);
  nor (_29795_, _29794_, _29790_);
  nor (_29796_, _10639_, _10286_);
  nor (_29797_, _29796_, _10643_);
  not (_29798_, _29797_);
  nor (_29799_, _29798_, _29795_);
  and (_29801_, _10286_, _10627_);
  nor (_29802_, _29632_, _10627_);
  or (_29803_, _29802_, _29801_);
  and (_29804_, _29803_, _10643_);
  nor (_29805_, _29804_, _29799_);
  nor (_29806_, _29805_, _10656_);
  nor (_29807_, _29607_, _10654_);
  nor (_29808_, _29807_, _10659_);
  not (_29809_, _29808_);
  or (_29810_, _29809_, _29806_);
  nor (_29812_, _10658_, _10286_);
  nor (_29813_, _29812_, _03908_);
  and (_29814_, _29813_, _29810_);
  not (_29815_, _10076_);
  and (_29816_, _10119_, _03908_);
  nor (_29817_, _29816_, _29815_);
  not (_29818_, _29817_);
  nor (_29819_, _29818_, _29814_);
  nor (_29820_, _10286_, _10076_);
  or (_29821_, _29820_, _10074_);
  or (_29823_, _29821_, _29819_);
  and (_29824_, _29632_, _08297_);
  nor (_29825_, _10286_, _08297_);
  nor (_29826_, _29825_, _10075_);
  not (_29827_, _29826_);
  nor (_29828_, _29827_, _29824_);
  nor (_29829_, _29828_, _10670_);
  and (_29830_, _29829_, _29823_);
  or (_29831_, _29830_, _29614_);
  nand (_29832_, _29831_, _08581_);
  nor (_29833_, _10286_, _08581_);
  nor (_29834_, _29833_, _03914_);
  nand (_29835_, _29834_, _29832_);
  not (_29836_, _10065_);
  and (_29837_, _10119_, _03914_);
  nor (_29838_, _29837_, _29836_);
  and (_29839_, _29838_, _29835_);
  or (_29840_, _29839_, _29612_);
  and (_29841_, _29632_, \oc8051_golden_model_1.PSW [7]);
  nor (_29842_, _10286_, \oc8051_golden_model_1.PSW [7]);
  nor (_29844_, _29842_, _10064_);
  not (_29845_, _29844_);
  nor (_29846_, _29845_, _29841_);
  nor (_29847_, _29846_, _10688_);
  and (_29848_, _29847_, _29840_);
  or (_29849_, _29848_, _29610_);
  nand (_29850_, _29849_, _08628_);
  nor (_29851_, _10286_, _08628_);
  nor (_29852_, _29851_, _08657_);
  and (_29853_, _29852_, _29850_);
  and (_29855_, _29606_, _08657_);
  or (_29856_, _29855_, _04034_);
  nor (_29857_, _29856_, _29853_);
  nor (_29858_, _05119_, _10704_);
  or (_29859_, _29858_, _29857_);
  nand (_29860_, _29859_, _03384_);
  and (_29861_, _29639_, _03383_);
  nor (_29862_, _29861_, _03913_);
  nand (_29863_, _29862_, _29860_);
  nor (_29864_, _10119_, _10906_);
  and (_29866_, _29625_, _10906_);
  or (_29867_, _29866_, _04097_);
  nor (_29868_, _29867_, _29864_);
  nor (_29869_, _29868_, _10712_);
  and (_29870_, _29869_, _29863_);
  or (_29871_, _29870_, _29609_);
  nand (_29872_, _29871_, _10056_);
  nor (_29873_, _10286_, _10056_);
  nor (_29874_, _29873_, _08772_);
  and (_29875_, _29874_, _29872_);
  and (_29877_, _29606_, _08772_);
  or (_29878_, _29877_, _03777_);
  nor (_29879_, _29878_, _29875_);
  nor (_29880_, _05119_, _03778_);
  or (_29881_, _29880_, _29879_);
  nand (_29882_, _29881_, _03411_);
  and (_29883_, _29639_, _03410_);
  nor (_29884_, _29883_, _03775_);
  nand (_29885_, _29884_, _29882_);
  nor (_29886_, _29675_, _10906_);
  and (_29888_, _10120_, _10906_);
  nor (_29889_, _29888_, _29886_);
  and (_29890_, _29889_, _03775_);
  nor (_29891_, _29890_, _10937_);
  nand (_29892_, _29891_, _29885_);
  nor (_29893_, _29606_, _10936_);
  nor (_29894_, _29893_, _03773_);
  nand (_29895_, _29894_, _29892_);
  and (_29896_, _10286_, _03773_);
  nor (_29897_, _29896_, _26446_);
  nand (_29899_, _29897_, _29895_);
  nor (_29900_, _29606_, _10943_);
  nor (_29901_, _29900_, _03899_);
  and (_29902_, _29901_, _29899_);
  nor (_29903_, _03900_, _03678_);
  or (_29904_, _29903_, _03414_);
  or (_29905_, _29904_, _29902_);
  and (_29906_, _29639_, _03414_);
  nor (_29907_, _29906_, _03374_);
  nand (_29908_, _29907_, _29905_);
  and (_29910_, _29889_, _03374_);
  nor (_29911_, _29910_, _10959_);
  nand (_29912_, _29911_, _29908_);
  nor (_29913_, _29606_, _10958_);
  nor (_29914_, _29913_, _03772_);
  nand (_29915_, _29914_, _29912_);
  and (_29916_, _10286_, _03772_);
  nor (_29917_, _29916_, _28254_);
  nand (_29918_, _29917_, _29915_);
  nor (_29919_, _29606_, _10965_);
  nor (_29921_, _29919_, _03901_);
  and (_29922_, _29921_, _29918_);
  nor (_29923_, _10969_, _03678_);
  or (_29924_, _29923_, _03413_);
  nor (_29925_, _29924_, _29922_);
  and (_29926_, _29639_, _03413_);
  or (_29927_, _29926_, _29925_);
  and (_29928_, _29927_, _10976_);
  nor (_29929_, _29928_, _29608_);
  or (_29930_, _29929_, _43156_);
  or (_29932_, _43152_, \oc8051_golden_model_1.PC [11]);
  and (_29933_, _29932_, _41894_);
  and (_43522_, _29933_, _29930_);
  nor (_29934_, _10048_, \oc8051_golden_model_1.PC [12]);
  nor (_29935_, _29934_, _10049_);
  not (_29936_, _29935_);
  and (_29937_, _29936_, _08772_);
  not (_29938_, _10283_);
  nor (_29939_, _29938_, _10065_);
  and (_29940_, _10111_, _03914_);
  nor (_29942_, _29935_, _10072_);
  nor (_29943_, _29938_, _10076_);
  and (_29944_, _10111_, _03908_);
  nor (_29945_, _29935_, _10654_);
  nor (_29946_, _10639_, _29938_);
  and (_29947_, _10111_, _03897_);
  nor (_29948_, _29935_, _10082_);
  nor (_29949_, _10583_, _29938_);
  nor (_29950_, _10610_, \oc8051_golden_model_1.DPH [4]);
  nor (_29951_, _29950_, _10611_);
  nor (_29953_, _29951_, _10581_);
  and (_29954_, _10364_, _10361_);
  nor (_29955_, _29954_, _10365_);
  and (_29956_, _29955_, _10564_);
  or (_29957_, _10523_, _10283_);
  or (_29958_, _29935_, _10421_);
  or (_29959_, _10416_, _10283_);
  and (_29960_, _10204_, _10201_);
  nor (_29961_, _29960_, _10205_);
  or (_29962_, _29961_, _10265_);
  nand (_29964_, _10265_, _10111_);
  and (_29965_, _29964_, _03850_);
  and (_29966_, _29965_, _29962_);
  and (_29967_, _29955_, _10383_);
  and (_29968_, _10382_, _10283_);
  or (_29969_, _29968_, _29967_);
  or (_29970_, _29969_, _04266_);
  nand (_29971_, _29938_, _03768_);
  and (_29972_, _29971_, _10402_);
  nand (_29973_, _29938_, _04230_);
  or (_29974_, _04707_, \oc8051_golden_model_1.PC [12]);
  or (_29975_, _29974_, _05011_);
  and (_29976_, _29975_, _29973_);
  or (_29977_, _29976_, _04263_);
  or (_29978_, _29935_, _25870_);
  and (_29979_, _29978_, _29977_);
  or (_29980_, _29979_, _03768_);
  and (_29981_, _29980_, _29972_);
  nor (_29982_, _29936_, _10402_);
  or (_29983_, _29982_, _04267_);
  or (_29986_, _29983_, _29981_);
  and (_29987_, _29986_, _26151_);
  and (_29988_, _29987_, _29970_);
  or (_29989_, _29988_, _29966_);
  and (_29990_, _29989_, _10412_);
  not (_29991_, _10416_);
  nor (_29992_, _29936_, _10417_);
  or (_29993_, _29992_, _29991_);
  or (_29994_, _29993_, _29990_);
  and (_29995_, _29994_, _29959_);
  or (_29997_, _29995_, _26168_);
  and (_29998_, _29997_, _29958_);
  or (_29999_, _29998_, _03854_);
  nand (_30000_, _29938_, _03854_);
  and (_30001_, _30000_, _10431_);
  and (_30002_, _30001_, _29999_);
  nor (_30003_, _29936_, _10431_);
  or (_30004_, _30003_, _30002_);
  and (_30005_, _30004_, _10257_);
  or (_30006_, _10257_, _29938_);
  nand (_30008_, _30006_, _10441_);
  or (_30009_, _30008_, _30005_);
  and (_30010_, _10476_, _10110_);
  not (_30011_, _29961_);
  nor (_30012_, _30011_, _10476_);
  or (_30013_, _30012_, _30010_);
  or (_30014_, _30013_, _10441_);
  and (_30015_, _30014_, _30009_);
  or (_30016_, _30015_, _03925_);
  and (_30017_, _10249_, _10110_);
  nor (_30019_, _30011_, _10249_);
  or (_30020_, _30019_, _30017_);
  or (_30021_, _30020_, _10444_);
  and (_30022_, _30021_, _03918_);
  and (_30023_, _30022_, _30016_);
  nor (_30024_, _30011_, _10498_);
  and (_30025_, _10498_, _10110_);
  or (_30026_, _30025_, _30024_);
  and (_30027_, _30026_, _03868_);
  or (_30028_, _30027_, _30023_);
  and (_30030_, _30028_, _10486_);
  or (_30031_, _29961_, _10515_);
  nand (_30032_, _10515_, _10111_);
  and (_30033_, _30032_, _03920_);
  and (_30034_, _30033_, _30031_);
  nand (_30035_, _29935_, _10485_);
  nand (_30036_, _30035_, _10523_);
  or (_30037_, _30036_, _30034_);
  or (_30038_, _30037_, _30030_);
  and (_30039_, _30038_, _29957_);
  or (_30041_, _30039_, _10093_);
  or (_30042_, _29935_, _10092_);
  and (_30043_, _30042_, _10531_);
  and (_30044_, _30043_, _30041_);
  or (_30045_, _10531_, _29938_);
  nand (_30046_, _30045_, _10087_);
  or (_30047_, _30046_, _30044_);
  or (_30048_, _29935_, _10087_);
  and (_30049_, _30048_, _10085_);
  and (_30050_, _30049_, _30047_);
  nor (_30052_, _29938_, _10085_);
  or (_30053_, _30052_, _03425_);
  or (_30054_, _30053_, _30050_);
  nand (_30055_, _29936_, _03425_);
  and (_30056_, _30055_, _10542_);
  and (_30057_, _30056_, _30054_);
  nor (_30058_, _10542_, _29938_);
  or (_30059_, _30058_, _03921_);
  or (_30060_, _30059_, _30057_);
  nand (_30061_, _10111_, _03921_);
  and (_30063_, _30061_, _07926_);
  and (_30064_, _30063_, _30060_);
  nor (_30065_, _29938_, _07926_);
  or (_30066_, _30065_, _03455_);
  or (_30067_, _30066_, _30064_);
  nand (_30068_, _10111_, _03455_);
  and (_30069_, _30068_, _10556_);
  and (_30070_, _30069_, _30067_);
  nor (_30071_, _29936_, _10556_);
  or (_30072_, _30071_, _10561_);
  or (_30074_, _30072_, _30070_);
  or (_30075_, _10560_, _10283_);
  and (_30076_, _30075_, _10565_);
  and (_30077_, _30076_, _30074_);
  or (_30078_, _30077_, _29956_);
  nor (_30079_, _30078_, _06309_);
  nor (_30080_, _10283_, _06138_);
  nor (_30081_, _30080_, _30079_);
  and (_30082_, _30081_, _04778_);
  and (_30083_, _10110_, _03903_);
  or (_30085_, _30083_, _30082_);
  and (_30086_, _30085_, _08493_);
  and (_30087_, _10283_, _08492_);
  or (_30088_, _30087_, _10580_);
  nor (_30089_, _30088_, _30086_);
  or (_30090_, _30089_, _10584_);
  nor (_30091_, _30090_, _29953_);
  nor (_30092_, _30091_, _29949_);
  nor (_30093_, _30092_, _10620_);
  and (_30094_, _10283_, _08826_);
  and (_30096_, _29955_, _10627_);
  or (_30097_, _30096_, _30094_);
  and (_30098_, _30097_, _10620_);
  nor (_30099_, _30098_, _10625_);
  not (_30100_, _30099_);
  nor (_30101_, _30100_, _30093_);
  or (_30102_, _30101_, _10080_);
  nor (_30103_, _30102_, _29948_);
  nor (_30104_, _29938_, _10079_);
  nor (_30105_, _30104_, _03897_);
  not (_30107_, _30105_);
  nor (_30108_, _30107_, _30103_);
  or (_30109_, _30108_, _29791_);
  nor (_30110_, _30109_, _29947_);
  nor (_30111_, _30110_, _29946_);
  nor (_30112_, _30111_, _10643_);
  nor (_30113_, _29955_, _10627_);
  nor (_30114_, _10283_, _08826_);
  nor (_30115_, _30114_, _10644_);
  not (_30116_, _30115_);
  nor (_30118_, _30116_, _30113_);
  nor (_30119_, _30118_, _10656_);
  not (_30120_, _30119_);
  nor (_30121_, _30120_, _30112_);
  or (_30122_, _30121_, _10659_);
  nor (_30123_, _30122_, _29945_);
  nor (_30124_, _10658_, _29938_);
  nor (_30125_, _30124_, _03908_);
  not (_30126_, _30125_);
  nor (_30127_, _30126_, _30123_);
  or (_30129_, _30127_, _29815_);
  nor (_30130_, _30129_, _29944_);
  nor (_30131_, _30130_, _29943_);
  nor (_30132_, _30131_, _10074_);
  nor (_30133_, _29955_, \oc8051_golden_model_1.PSW [7]);
  nor (_30134_, _10283_, _08297_);
  nor (_30135_, _30134_, _10075_);
  not (_30136_, _30135_);
  nor (_30137_, _30136_, _30133_);
  nor (_30138_, _30137_, _10670_);
  not (_30140_, _30138_);
  nor (_30141_, _30140_, _30132_);
  or (_30142_, _30141_, _08582_);
  nor (_30143_, _30142_, _29942_);
  nor (_30144_, _29938_, _08581_);
  nor (_30145_, _30144_, _03914_);
  not (_30146_, _30145_);
  nor (_30147_, _30146_, _30143_);
  or (_30148_, _30147_, _29836_);
  nor (_30149_, _30148_, _29940_);
  or (_30151_, _30149_, _29939_);
  nand (_30152_, _30151_, _10064_);
  nor (_30153_, _29955_, _08297_);
  nor (_30154_, _10283_, \oc8051_golden_model_1.PSW [7]);
  nor (_30155_, _30154_, _10064_);
  not (_30156_, _30155_);
  nor (_30157_, _30156_, _30153_);
  nor (_30158_, _30157_, _10688_);
  nand (_30159_, _30158_, _30152_);
  nor (_30160_, _29935_, _10061_);
  nor (_30162_, _30160_, _08629_);
  nand (_30163_, _30162_, _30159_);
  nor (_30164_, _29938_, _08628_);
  nor (_30165_, _30164_, _08657_);
  nand (_30166_, _30165_, _30163_);
  and (_30167_, _29936_, _08657_);
  nor (_30168_, _30167_, _04034_);
  and (_30169_, _30168_, _30166_);
  and (_30170_, _05950_, _04034_);
  or (_30171_, _30170_, _03383_);
  or (_30173_, _30171_, _30169_);
  and (_30174_, _29938_, _03383_);
  nor (_30175_, _30174_, _03913_);
  nand (_30176_, _30175_, _30173_);
  nor (_30177_, _10110_, _10906_);
  and (_30178_, _30011_, _10906_);
  or (_30179_, _30178_, _04097_);
  nor (_30180_, _30179_, _30177_);
  nor (_30181_, _30180_, _10712_);
  nand (_30182_, _30181_, _30176_);
  nor (_30184_, _29935_, _10059_);
  nor (_30185_, _30184_, _10057_);
  nand (_30186_, _30185_, _30182_);
  nor (_30187_, _29938_, _10056_);
  nor (_30188_, _30187_, _08772_);
  and (_30189_, _30188_, _30186_);
  or (_30190_, _30189_, _29937_);
  nand (_30191_, _30190_, _03778_);
  nor (_30192_, _05950_, _03778_);
  nor (_30193_, _30192_, _03410_);
  and (_30195_, _30193_, _30191_);
  and (_30196_, _10283_, _03410_);
  or (_30197_, _30196_, _03775_);
  nor (_30198_, _30197_, _30195_);
  nor (_30199_, _29961_, _10906_);
  and (_30200_, _10111_, _10906_);
  nor (_30201_, _30200_, _30199_);
  nor (_30202_, _30201_, _03776_);
  or (_30203_, _30202_, _30198_);
  and (_30204_, _30203_, _10936_);
  nor (_30206_, _29935_, _10936_);
  or (_30207_, _30206_, _30204_);
  nand (_30208_, _30207_, _03774_);
  and (_30209_, _29938_, _03773_);
  nor (_30210_, _30209_, _26446_);
  nand (_30211_, _30210_, _30208_);
  nor (_30212_, _29936_, _10943_);
  nor (_30213_, _30212_, _03899_);
  nand (_30214_, _30213_, _30211_);
  and (_30215_, _04526_, _03899_);
  nor (_30217_, _30215_, _03414_);
  and (_30218_, _30217_, _30214_);
  and (_30219_, _10283_, _03414_);
  or (_30220_, _30219_, _03374_);
  or (_30221_, _30220_, _30218_);
  nor (_30222_, _30201_, _03375_);
  nor (_30223_, _30222_, _10959_);
  nand (_30224_, _30223_, _30221_);
  nor (_30225_, _29936_, _10958_);
  nor (_30226_, _30225_, _03772_);
  nand (_30228_, _30226_, _30224_);
  and (_30229_, _29938_, _03772_);
  nor (_30230_, _30229_, _28254_);
  nand (_30231_, _30230_, _30228_);
  nor (_30232_, _29936_, _10965_);
  nor (_30233_, _30232_, _03901_);
  nand (_30234_, _30233_, _30231_);
  and (_30235_, _04526_, _03901_);
  nor (_30236_, _30235_, _03413_);
  and (_30237_, _30236_, _30234_);
  and (_30239_, _10283_, _03413_);
  or (_30240_, _30239_, _30237_);
  and (_30241_, _30240_, _10976_);
  and (_30242_, _29935_, _10042_);
  or (_30243_, _30242_, _30241_);
  or (_30244_, _30243_, _43156_);
  or (_30245_, _43152_, \oc8051_golden_model_1.PC [12]);
  and (_30246_, _30245_, _41894_);
  and (_43523_, _30246_, _30244_);
  nor (_30247_, _10049_, \oc8051_golden_model_1.PC [13]);
  nor (_30249_, _30247_, _10050_);
  nor (_30250_, _30249_, _10059_);
  nor (_30251_, _30249_, _10061_);
  nor (_30252_, _10279_, _10065_);
  or (_30253_, _30252_, _10063_);
  nor (_30254_, _30249_, _10072_);
  nor (_30255_, _10279_, _10076_);
  or (_30256_, _30255_, _10074_);
  nor (_30257_, _10639_, _10279_);
  and (_30258_, _10279_, _08826_);
  or (_30260_, _10281_, _10280_);
  not (_30261_, _30260_);
  nor (_30262_, _30261_, _10366_);
  and (_30263_, _30261_, _10366_);
  nor (_30264_, _30263_, _30262_);
  nor (_30265_, _30264_, _08826_);
  or (_30266_, _30265_, _30258_);
  and (_30267_, _30266_, _10620_);
  nor (_30268_, _10611_, \oc8051_golden_model_1.DPH [5]);
  or (_30269_, _30268_, _10612_);
  or (_30271_, _30269_, _10581_);
  nor (_30272_, _10279_, _06138_);
  and (_30273_, _10105_, _03455_);
  or (_30274_, _10108_, _10107_);
  not (_30275_, _30274_);
  nor (_30276_, _30275_, _10206_);
  and (_30277_, _30275_, _10206_);
  nor (_30278_, _30277_, _30276_);
  nor (_30279_, _30278_, _10249_);
  and (_30280_, _10249_, _10105_);
  nor (_30282_, _30280_, _30279_);
  or (_30283_, _30282_, _10444_);
  or (_30284_, _10257_, _10279_);
  and (_30285_, _10279_, _03854_);
  not (_30286_, _30278_);
  or (_30287_, _30286_, _10265_);
  and (_30288_, _30287_, _03850_);
  nand (_30289_, _10265_, _10106_);
  and (_30290_, _30289_, _30288_);
  nor (_30291_, _30264_, _10382_);
  and (_30293_, _10382_, _10279_);
  or (_30294_, _30293_, _30291_);
  and (_30295_, _30294_, _04267_);
  or (_30296_, _30249_, _29316_);
  not (_30297_, _10279_);
  nand (_30298_, _30297_, _04230_);
  or (_30299_, _03768_, \oc8051_golden_model_1.PC [13]);
  or (_30300_, _30299_, _04707_);
  or (_30301_, _30300_, _05011_);
  and (_30302_, _30301_, _30298_);
  or (_30303_, _30302_, _04263_);
  nand (_30304_, _30297_, _03768_);
  and (_30305_, _30304_, _30303_);
  or (_30306_, _30305_, _26516_);
  and (_30307_, _30306_, _04266_);
  and (_30308_, _30307_, _30296_);
  or (_30309_, _30308_, _04716_);
  or (_30310_, _30309_, _30295_);
  and (_30311_, _30310_, _04722_);
  or (_30312_, _30311_, _10413_);
  or (_30315_, _30312_, _30290_);
  or (_30316_, _30249_, _10417_);
  and (_30317_, _30316_, _10416_);
  and (_30318_, _30317_, _30315_);
  or (_30319_, _10416_, _30297_);
  nand (_30320_, _30319_, _10421_);
  or (_30321_, _30320_, _30318_);
  or (_30322_, _30249_, _10421_);
  and (_30323_, _30322_, _03855_);
  and (_30324_, _30323_, _30321_);
  or (_30326_, _30324_, _30285_);
  and (_30327_, _30326_, _10431_);
  not (_30328_, _30249_);
  or (_30329_, _30328_, _10431_);
  nand (_30330_, _30329_, _10257_);
  or (_30331_, _30330_, _30327_);
  and (_30332_, _30331_, _30284_);
  or (_30333_, _30332_, _10442_);
  and (_30334_, _10476_, _10105_);
  nor (_30335_, _30278_, _10476_);
  or (_30337_, _30335_, _30334_);
  or (_30338_, _30337_, _10441_);
  and (_30339_, _30338_, _10444_);
  nand (_30340_, _30339_, _30333_);
  and (_30341_, _30340_, _03918_);
  and (_30342_, _30341_, _30283_);
  and (_30343_, _10498_, _10105_);
  nor (_30344_, _30278_, _10498_);
  or (_30345_, _30344_, _03918_);
  nor (_30346_, _30345_, _30343_);
  or (_30348_, _30346_, _27224_);
  or (_30349_, _30348_, _30342_);
  and (_30350_, _30278_, _29696_);
  and (_30351_, _10515_, _10106_);
  or (_30352_, _30351_, _11857_);
  or (_30353_, _30352_, _30350_);
  nand (_30354_, _30249_, _10485_);
  and (_30355_, _30354_, _10523_);
  and (_30356_, _30355_, _30353_);
  and (_30357_, _30356_, _30349_);
  nor (_30359_, _10523_, _10279_);
  or (_30360_, _30359_, _10093_);
  or (_30361_, _30360_, _30357_);
  or (_30362_, _30328_, _10092_);
  and (_30363_, _30362_, _10531_);
  nand (_30364_, _30363_, _30361_);
  or (_30365_, _10531_, _10279_);
  and (_30366_, _30365_, _10087_);
  and (_30367_, _30366_, _30364_);
  nor (_30368_, _30328_, _10087_);
  nor (_30370_, _30368_, _10086_);
  not (_30371_, _30370_);
  nor (_30372_, _30371_, _30367_);
  nor (_30373_, _10279_, _10085_);
  nor (_30374_, _30373_, _03425_);
  not (_30375_, _30374_);
  nor (_30376_, _30375_, _30372_);
  and (_30377_, _30249_, _03425_);
  nor (_30378_, _30377_, _10543_);
  not (_30380_, _30378_);
  nor (_30383_, _30380_, _30376_);
  nor (_30385_, _10542_, _10279_);
  nor (_30387_, _30385_, _03921_);
  not (_30389_, _30387_);
  nor (_30391_, _30389_, _30383_);
  and (_30393_, _10105_, _03921_);
  nor (_30395_, _30393_, _07927_);
  not (_30397_, _30395_);
  nor (_30399_, _30397_, _30391_);
  nor (_30401_, _10279_, _07926_);
  nor (_30403_, _30401_, _03455_);
  not (_30404_, _30403_);
  nor (_30405_, _30404_, _30399_);
  nor (_30406_, _30405_, _30273_);
  nor (_30407_, _30406_, _10558_);
  nor (_30408_, _30328_, _10556_);
  nor (_30409_, _30408_, _10561_);
  not (_30410_, _30409_);
  nor (_30411_, _30410_, _30407_);
  nor (_30412_, _10560_, _10279_);
  nor (_30414_, _30412_, _10564_);
  not (_30415_, _30414_);
  nor (_30416_, _30415_, _30411_);
  nor (_30417_, _30264_, _10565_);
  nor (_30418_, _30417_, _06309_);
  not (_30419_, _30418_);
  nor (_30420_, _30419_, _30416_);
  nor (_30421_, _30420_, _30272_);
  and (_30422_, _30421_, _04778_);
  and (_30423_, _10105_, _03903_);
  or (_30425_, _30423_, _30422_);
  and (_30426_, _30425_, _08493_);
  and (_30427_, _10279_, _08492_);
  nor (_30428_, _30427_, _30426_);
  nor (_30429_, _30428_, _10580_);
  nor (_30430_, _30429_, _10584_);
  and (_30431_, _30430_, _30271_);
  nor (_30432_, _10583_, _10279_);
  nor (_30433_, _30432_, _10620_);
  not (_30434_, _30433_);
  nor (_30436_, _30434_, _30431_);
  nor (_30437_, _30436_, _30267_);
  nor (_30438_, _30437_, _10625_);
  nor (_30439_, _30328_, _10082_);
  nor (_30440_, _30439_, _10080_);
  not (_30441_, _30440_);
  nor (_30442_, _30441_, _30438_);
  nor (_30443_, _10279_, _10079_);
  nor (_30444_, _30443_, _03897_);
  not (_30445_, _30444_);
  nor (_30447_, _30445_, _30442_);
  and (_30448_, _10105_, _03897_);
  nor (_30449_, _30448_, _29791_);
  not (_30450_, _30449_);
  nor (_30451_, _30450_, _30447_);
  or (_30452_, _30451_, _10643_);
  nor (_30453_, _30452_, _30257_);
  and (_30454_, _30264_, _08826_);
  nor (_30455_, _10279_, _08826_);
  nor (_30456_, _30455_, _10644_);
  not (_30458_, _30456_);
  nor (_30459_, _30458_, _30454_);
  nor (_30460_, _30459_, _30453_);
  or (_30461_, _30460_, _10656_);
  or (_30462_, _30328_, _10654_);
  and (_30463_, _30462_, _10658_);
  and (_30464_, _30463_, _30461_);
  nor (_30465_, _10658_, _10279_);
  nor (_30466_, _30465_, _03908_);
  not (_30467_, _30466_);
  nor (_30469_, _30467_, _30464_);
  and (_30470_, _10105_, _03908_);
  nor (_30471_, _30470_, _29815_);
  not (_30472_, _30471_);
  nor (_30473_, _30472_, _30469_);
  or (_30474_, _30473_, _30256_);
  and (_30475_, _30264_, _08297_);
  nor (_30476_, _10279_, _08297_);
  nor (_30477_, _30476_, _10075_);
  not (_30478_, _30477_);
  nor (_30480_, _30478_, _30475_);
  nor (_30481_, _30480_, _10670_);
  and (_30482_, _30481_, _30474_);
  or (_30483_, _30482_, _30254_);
  nand (_30484_, _30483_, _08581_);
  nor (_30485_, _10279_, _08581_);
  nor (_30486_, _30485_, _03914_);
  nand (_30487_, _30486_, _30484_);
  and (_30488_, _10105_, _03914_);
  nor (_30489_, _30488_, _29836_);
  and (_30491_, _30489_, _30487_);
  or (_30492_, _30491_, _30253_);
  and (_30493_, _30264_, \oc8051_golden_model_1.PSW [7]);
  nor (_30494_, _10279_, \oc8051_golden_model_1.PSW [7]);
  nor (_30495_, _30494_, _10064_);
  not (_30496_, _30495_);
  nor (_30497_, _30496_, _30493_);
  nor (_30498_, _30497_, _10688_);
  and (_30499_, _30498_, _30492_);
  or (_30500_, _30499_, _30251_);
  nand (_30502_, _30500_, _08628_);
  nor (_30503_, _10279_, _08628_);
  nor (_30504_, _30503_, _08657_);
  and (_30505_, _30504_, _30502_);
  and (_30506_, _30249_, _08657_);
  or (_30507_, _30506_, _04034_);
  nor (_30508_, _30507_, _30505_);
  nor (_30509_, _05857_, _10704_);
  or (_30510_, _30509_, _30508_);
  nand (_30511_, _30510_, _03384_);
  and (_30513_, _30297_, _03383_);
  nor (_30514_, _30513_, _03913_);
  nand (_30515_, _30514_, _30511_);
  and (_30516_, _30278_, _10906_);
  nor (_30517_, _10105_, _10906_);
  or (_30518_, _30517_, _04097_);
  or (_30519_, _30518_, _30516_);
  and (_30520_, _30519_, _10059_);
  and (_30521_, _30520_, _30515_);
  or (_30522_, _30521_, _30250_);
  nand (_30524_, _30522_, _10056_);
  nor (_30525_, _10279_, _10056_);
  nor (_30526_, _30525_, _08772_);
  and (_30527_, _30526_, _30524_);
  and (_30528_, _30249_, _08772_);
  or (_30529_, _30528_, _03777_);
  nor (_30530_, _30529_, _30527_);
  nor (_30531_, _05857_, _03778_);
  or (_30532_, _30531_, _30530_);
  nand (_30533_, _30532_, _03411_);
  and (_30535_, _30297_, _03410_);
  nor (_30536_, _30535_, _03775_);
  nand (_30537_, _30536_, _30533_);
  and (_30538_, _10106_, _10906_);
  nor (_30539_, _30286_, _10906_);
  nor (_30540_, _30539_, _30538_);
  and (_30541_, _30540_, _03775_);
  nor (_30542_, _30541_, _10937_);
  nand (_30543_, _30542_, _30537_);
  nor (_30544_, _30249_, _10936_);
  nor (_30546_, _30544_, _03773_);
  nand (_30547_, _30546_, _30543_);
  and (_30548_, _10279_, _03773_);
  nor (_30549_, _30548_, _26446_);
  nand (_30550_, _30549_, _30547_);
  nor (_30551_, _30249_, _10943_);
  nor (_30552_, _30551_, _03899_);
  and (_30553_, _30552_, _30550_);
  nor (_30554_, _04093_, _03900_);
  or (_30555_, _30554_, _03414_);
  or (_30557_, _30555_, _30553_);
  and (_30558_, _30297_, _03414_);
  nor (_30559_, _30558_, _03374_);
  nand (_30560_, _30559_, _30557_);
  and (_30561_, _30540_, _03374_);
  nor (_30562_, _30561_, _10959_);
  nand (_30563_, _30562_, _30560_);
  nor (_30564_, _30249_, _10958_);
  nor (_30565_, _30564_, _03772_);
  nand (_30566_, _30565_, _30563_);
  and (_30568_, _10279_, _03772_);
  nor (_30569_, _30568_, _28254_);
  nand (_30570_, _30569_, _30566_);
  nor (_30571_, _30249_, _10965_);
  nor (_30572_, _30571_, _03901_);
  nand (_30573_, _30572_, _30570_);
  nor (_30574_, _04093_, _10969_);
  nor (_30575_, _30574_, _03413_);
  and (_30576_, _30575_, _30573_);
  and (_30577_, _30297_, _03413_);
  or (_30578_, _30577_, _30576_);
  and (_30579_, _30578_, _10976_);
  and (_30580_, _30328_, _10042_);
  nor (_30581_, _30580_, _30579_);
  or (_30582_, _30581_, _43156_);
  or (_30583_, _43152_, \oc8051_golden_model_1.PC [13]);
  and (_30584_, _30583_, _41894_);
  and (_43524_, _30584_, _30582_);
  nand (_30585_, _03901_, _03810_);
  or (_30586_, _10050_, \oc8051_golden_model_1.PC [14]);
  and (_30588_, _30586_, _10051_);
  or (_30589_, _30588_, _08773_);
  and (_30590_, _10274_, _29836_);
  and (_30591_, _10274_, _29815_);
  and (_30592_, _29791_, _10274_);
  and (_30593_, _10584_, _10274_);
  nor (_30594_, _10369_, _10277_);
  nor (_30595_, _30594_, _10370_);
  and (_30596_, _30595_, _10564_);
  or (_30597_, _10523_, _10274_);
  nor (_30599_, _10209_, _10103_);
  nor (_30600_, _30599_, _10210_);
  or (_30601_, _30600_, _10476_);
  nand (_30602_, _10476_, _10100_);
  and (_30603_, _30602_, _30601_);
  or (_30604_, _30603_, _10441_);
  or (_30605_, _30588_, _10421_);
  or (_30606_, _10416_, _10274_);
  or (_30607_, _30600_, _10265_);
  and (_30608_, _30607_, _03850_);
  nand (_30610_, _10265_, _10100_);
  and (_30611_, _30610_, _30608_);
  and (_30612_, _30595_, _10383_);
  and (_30613_, _10382_, _10274_);
  or (_30614_, _30613_, _30612_);
  or (_30615_, _30614_, _04266_);
  or (_30616_, _10274_, _03770_);
  and (_30617_, _30616_, _10402_);
  or (_30618_, _10274_, _10389_);
  or (_30619_, _04707_, \oc8051_golden_model_1.PC [14]);
  or (_30621_, _30619_, _05011_);
  and (_30622_, _30621_, _30618_);
  or (_30623_, _30622_, _04263_);
  or (_30624_, _30588_, _25870_);
  and (_30625_, _30624_, _30623_);
  or (_30626_, _30625_, _03768_);
  and (_30627_, _30626_, _30617_);
  and (_30628_, _30588_, _26516_);
  or (_30629_, _30628_, _04267_);
  or (_30630_, _30629_, _30627_);
  and (_30632_, _30630_, _26151_);
  and (_30633_, _30632_, _30615_);
  or (_30634_, _30633_, _30611_);
  and (_30635_, _30634_, _10412_);
  not (_30636_, _10417_);
  and (_30637_, _30588_, _30636_);
  or (_30638_, _30637_, _29991_);
  or (_30639_, _30638_, _30635_);
  and (_30640_, _30639_, _30606_);
  or (_30641_, _30640_, _26168_);
  and (_30643_, _30641_, _30605_);
  or (_30644_, _30643_, _03854_);
  or (_30645_, _10274_, _03855_);
  and (_30646_, _30645_, _10431_);
  and (_30647_, _30646_, _30644_);
  and (_30648_, _30588_, _10434_);
  or (_30649_, _30648_, _30647_);
  and (_30650_, _30649_, _10257_);
  and (_30651_, _10433_, _10274_);
  or (_30652_, _30651_, _10442_);
  or (_30654_, _30652_, _30650_);
  and (_30655_, _30654_, _30604_);
  or (_30656_, _30655_, _03925_);
  or (_30657_, _30600_, _10249_);
  nand (_30658_, _10249_, _10100_);
  and (_30659_, _30658_, _30657_);
  or (_30660_, _30659_, _10444_);
  and (_30661_, _30660_, _03918_);
  and (_30662_, _30661_, _30656_);
  and (_30663_, _10498_, _10099_);
  and (_30665_, _30600_, _10500_);
  or (_30666_, _30665_, _30663_);
  and (_30667_, _30666_, _03868_);
  or (_30668_, _30667_, _30662_);
  and (_30669_, _30668_, _10486_);
  or (_30670_, _30600_, _10515_);
  nand (_30671_, _10515_, _10100_);
  and (_30672_, _30671_, _03920_);
  and (_30673_, _30672_, _30670_);
  nand (_30674_, _30588_, _10485_);
  nand (_30676_, _30674_, _10523_);
  or (_30677_, _30676_, _30673_);
  or (_30678_, _30677_, _30669_);
  and (_30679_, _30678_, _30597_);
  or (_30680_, _30679_, _10093_);
  or (_30681_, _30588_, _10092_);
  and (_30682_, _30681_, _10531_);
  and (_30683_, _30682_, _30680_);
  not (_30684_, _10274_);
  or (_30685_, _10531_, _30684_);
  nand (_30687_, _30685_, _10087_);
  or (_30688_, _30687_, _30683_);
  or (_30689_, _30588_, _10087_);
  and (_30690_, _30689_, _10085_);
  and (_30691_, _30690_, _30688_);
  nor (_30692_, _30684_, _10085_);
  or (_30693_, _30692_, _03425_);
  or (_30694_, _30693_, _30691_);
  or (_30695_, _30588_, _03426_);
  and (_30696_, _30695_, _10542_);
  and (_30698_, _30696_, _30694_);
  nor (_30699_, _10542_, _30684_);
  or (_30700_, _30699_, _03921_);
  or (_30701_, _30700_, _30698_);
  or (_30702_, _10099_, _09861_);
  and (_30703_, _30702_, _07926_);
  and (_30704_, _30703_, _30701_);
  nor (_30705_, _30684_, _07926_);
  or (_30706_, _30705_, _03455_);
  or (_30707_, _30706_, _30704_);
  or (_30709_, _10099_, _03820_);
  and (_30710_, _30709_, _10556_);
  and (_30711_, _30710_, _30707_);
  and (_30712_, _30588_, _10558_);
  or (_30713_, _30712_, _10561_);
  or (_30714_, _30713_, _30711_);
  or (_30715_, _10560_, _10274_);
  and (_30716_, _30715_, _10565_);
  and (_30717_, _30716_, _30714_);
  or (_30718_, _30717_, _30596_);
  and (_30720_, _30718_, _06138_);
  nor (_30721_, _30684_, _06138_);
  or (_30722_, _30721_, _03903_);
  or (_30723_, _30722_, _30720_);
  or (_30724_, _10099_, _04778_);
  and (_30725_, _30724_, _08493_);
  and (_30726_, _30725_, _30723_);
  and (_30727_, _10274_, _08492_);
  or (_30728_, _30727_, _10580_);
  or (_30729_, _30728_, _30726_);
  nor (_30731_, _10612_, \oc8051_golden_model_1.DPH [6]);
  nor (_30732_, _30731_, _10613_);
  or (_30733_, _30732_, _10581_);
  and (_30734_, _30733_, _10583_);
  and (_30735_, _30734_, _30729_);
  or (_30736_, _30735_, _30593_);
  and (_30737_, _30736_, _10621_);
  or (_30738_, _30595_, _08826_);
  or (_30739_, _10274_, _10627_);
  and (_30740_, _30739_, _10620_);
  and (_30742_, _30740_, _30738_);
  or (_30743_, _30742_, _10625_);
  or (_30744_, _30743_, _30737_);
  or (_30745_, _30588_, _10082_);
  and (_30746_, _30745_, _10079_);
  and (_30747_, _30746_, _30744_);
  nor (_30748_, _30684_, _10079_);
  or (_30749_, _30748_, _03897_);
  or (_30750_, _30749_, _30747_);
  or (_30751_, _10099_, _04790_);
  and (_30753_, _30751_, _10639_);
  and (_30754_, _30753_, _30750_);
  or (_30755_, _30754_, _30592_);
  and (_30756_, _30755_, _10644_);
  or (_30757_, _30595_, _10627_);
  or (_30758_, _10274_, _08826_);
  and (_30759_, _30758_, _10643_);
  and (_30760_, _30759_, _30757_);
  or (_30761_, _30760_, _10656_);
  or (_30762_, _30761_, _30756_);
  or (_30764_, _30588_, _10654_);
  and (_30765_, _30764_, _10658_);
  and (_30766_, _30765_, _30762_);
  nor (_30767_, _10658_, _30684_);
  or (_30768_, _30767_, _03908_);
  or (_30769_, _30768_, _30766_);
  or (_30770_, _10099_, _03909_);
  and (_30771_, _30770_, _10076_);
  and (_30772_, _30771_, _30769_);
  or (_30773_, _30772_, _30591_);
  and (_30775_, _30773_, _10075_);
  or (_30776_, _30595_, \oc8051_golden_model_1.PSW [7]);
  or (_30777_, _10274_, _08297_);
  and (_30778_, _30777_, _10074_);
  and (_30779_, _30778_, _30776_);
  or (_30780_, _30779_, _10670_);
  or (_30781_, _30780_, _30775_);
  or (_30782_, _30588_, _10072_);
  and (_30783_, _30782_, _08581_);
  and (_30784_, _30783_, _30781_);
  nor (_30786_, _30684_, _08581_);
  or (_30787_, _30786_, _03914_);
  or (_30788_, _30787_, _30784_);
  or (_30789_, _10099_, _06567_);
  and (_30790_, _30789_, _10065_);
  and (_30791_, _30790_, _30788_);
  or (_30792_, _30791_, _30590_);
  and (_30793_, _30792_, _10064_);
  or (_30794_, _30595_, _08297_);
  or (_30795_, _10274_, \oc8051_golden_model_1.PSW [7]);
  and (_30796_, _30795_, _10063_);
  and (_30797_, _30796_, _30794_);
  or (_30798_, _30797_, _10688_);
  or (_30799_, _30798_, _30793_);
  or (_30800_, _30588_, _10061_);
  and (_30801_, _30800_, _08628_);
  and (_30802_, _30801_, _30799_);
  nor (_30803_, _30684_, _08628_);
  or (_30804_, _30803_, _08657_);
  or (_30805_, _30804_, _30802_);
  or (_30808_, _30588_, _08658_);
  and (_30809_, _30808_, _10704_);
  and (_30810_, _30809_, _30805_);
  and (_30811_, _06065_, _04034_);
  or (_30812_, _30811_, _03383_);
  or (_30813_, _30812_, _30810_);
  or (_30814_, _10274_, _03384_);
  and (_30815_, _30814_, _04097_);
  and (_30816_, _30815_, _30813_);
  or (_30817_, _10099_, _10906_);
  or (_30819_, _30600_, _10907_);
  and (_30820_, _30819_, _03913_);
  and (_30821_, _30820_, _30817_);
  or (_30822_, _30821_, _10712_);
  or (_30823_, _30822_, _30816_);
  or (_30824_, _30588_, _10059_);
  and (_30825_, _30824_, _10056_);
  and (_30826_, _30825_, _30823_);
  nor (_30827_, _30684_, _10056_);
  or (_30828_, _30827_, _08772_);
  or (_30830_, _30828_, _30826_);
  and (_30831_, _30830_, _30589_);
  or (_30832_, _30831_, _03777_);
  or (_30833_, _06065_, _03778_);
  and (_30834_, _30833_, _03411_);
  and (_30835_, _30834_, _30832_);
  and (_30836_, _10274_, _03410_);
  or (_30837_, _30836_, _03775_);
  or (_30838_, _30837_, _30835_);
  nand (_30839_, _10100_, _10906_);
  or (_30841_, _30600_, _10906_);
  and (_30842_, _30841_, _30839_);
  or (_30843_, _30842_, _03776_);
  and (_30844_, _30843_, _30838_);
  or (_30845_, _30844_, _10937_);
  or (_30846_, _30588_, _10936_);
  and (_30847_, _30846_, _30845_);
  or (_30848_, _30847_, _03773_);
  or (_30849_, _10274_, _03774_);
  and (_30850_, _30849_, _10943_);
  and (_30852_, _30850_, _30848_);
  and (_30853_, _30588_, _26446_);
  or (_30854_, _30853_, _03899_);
  or (_30855_, _30854_, _30852_);
  nand (_30856_, _03899_, _03810_);
  and (_30857_, _30856_, _10953_);
  and (_30858_, _30857_, _30855_);
  and (_30859_, _10274_, _03414_);
  or (_30860_, _30859_, _03374_);
  or (_30861_, _30860_, _30858_);
  or (_30863_, _30842_, _03375_);
  and (_30864_, _30863_, _10958_);
  and (_30865_, _30864_, _30861_);
  and (_30866_, _30588_, _10959_);
  or (_30867_, _30866_, _03772_);
  or (_30868_, _30867_, _30865_);
  or (_30869_, _10274_, _04060_);
  and (_30870_, _30869_, _10965_);
  and (_30871_, _30870_, _30868_);
  and (_30872_, _30588_, _28254_);
  or (_30874_, _30872_, _03901_);
  or (_30875_, _30874_, _30871_);
  and (_30876_, _30875_, _30585_);
  or (_30877_, _30876_, _03413_);
  or (_30878_, _10274_, _10977_);
  and (_30879_, _30878_, _10976_);
  and (_30880_, _30879_, _30877_);
  and (_30881_, _30588_, _10042_);
  or (_30882_, _30881_, _30880_);
  or (_30883_, _30882_, _43156_);
  or (_30885_, _43152_, \oc8051_golden_model_1.PC [14]);
  and (_30886_, _30885_, _41894_);
  and (_43525_, _30886_, _30883_);
  nor (_30887_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_30888_, _30887_, _05397_);
  not (_30889_, _05498_);
  and (_30890_, _30889_, \oc8051_golden_model_1.P2 [0]);
  nand (_30891_, _11126_, _03498_);
  or (_30892_, _11126_, _03498_);
  and (_30893_, _30892_, _30891_);
  and (_30895_, _30893_, _05498_);
  or (_30896_, _30895_, _30890_);
  and (_30897_, _30896_, _04018_);
  and (_30898_, _05498_, _06479_);
  or (_30899_, _30898_, _30890_);
  or (_30900_, _30899_, _04778_);
  and (_30901_, _11126_, _05498_);
  or (_30902_, _30901_, _30890_);
  or (_30903_, _30902_, _04722_);
  and (_30904_, _05498_, \oc8051_golden_model_1.ACC [0]);
  or (_30906_, _30904_, _30890_);
  and (_30907_, _30906_, _04707_);
  and (_30908_, _04708_, \oc8051_golden_model_1.P2 [0]);
  or (_30909_, _30908_, _03850_);
  or (_30910_, _30909_, _30907_);
  and (_30911_, _30910_, _03764_);
  and (_30912_, _30911_, _30903_);
  not (_30913_, _06106_);
  and (_30914_, _30913_, \oc8051_golden_model_1.P2 [0]);
  and (_30915_, _06112_, \oc8051_golden_model_1.P0 [0]);
  and (_30917_, _06106_, \oc8051_golden_model_1.P2 [0]);
  or (_30918_, _30917_, _30915_);
  and (_30919_, _06114_, \oc8051_golden_model_1.P1 [0]);
  and (_30920_, _06108_, \oc8051_golden_model_1.P3 [0]);
  or (_30921_, _30920_, _30919_);
  nor (_30922_, _30921_, _30918_);
  and (_30923_, _30922_, _10810_);
  nand (_30924_, _30923_, _10807_);
  or (_30925_, _30924_, _05715_);
  or (_30926_, _30925_, _05432_);
  and (_30928_, _30926_, _06106_);
  or (_30929_, _30928_, _30914_);
  and (_30930_, _30929_, _03763_);
  or (_30931_, _30930_, _30912_);
  and (_30932_, _30931_, _04733_);
  and (_30933_, _05498_, _04700_);
  or (_30934_, _30933_, _30890_);
  and (_30935_, _30934_, _03848_);
  or (_30936_, _30935_, _03854_);
  or (_30937_, _30936_, _30932_);
  or (_30939_, _30906_, _03855_);
  and (_30940_, _30939_, _03760_);
  and (_30941_, _30940_, _30937_);
  and (_30942_, _30890_, _03759_);
  or (_30943_, _30942_, _03752_);
  or (_30944_, _30943_, _30941_);
  or (_30945_, _30902_, _03753_);
  and (_30946_, _30945_, _03747_);
  and (_30947_, _30946_, _30944_);
  or (_30948_, _30914_, _14237_);
  and (_30950_, _30948_, _03746_);
  and (_30951_, _30950_, _30929_);
  or (_30952_, _30951_, _07927_);
  or (_30953_, _30952_, _30947_);
  and (_30954_, _06962_, _05498_);
  or (_30955_, _30890_, _03738_);
  or (_30956_, _30955_, _30954_);
  or (_30957_, _30934_, _07925_);
  and (_30958_, _30957_, _03820_);
  and (_30959_, _30958_, _30956_);
  and (_30961_, _30959_, _30953_);
  and (_30962_, _06505_, \oc8051_golden_model_1.P1 [0]);
  and (_30963_, _06507_, \oc8051_golden_model_1.P3 [0]);
  or (_30964_, _30963_, _30962_);
  nor (_30965_, _30964_, _12125_);
  nand (_30966_, _30965_, _12124_);
  or (_30967_, _30966_, _12117_);
  and (_30968_, _06501_, \oc8051_golden_model_1.P0 [0]);
  and (_30969_, _06515_, \oc8051_golden_model_1.P2 [0]);
  or (_30970_, _30969_, _12136_);
  nor (_30972_, _30970_, _30968_);
  nand (_30973_, _30972_, _12135_);
  nor (_30974_, _30973_, _30967_);
  nand (_30975_, _30974_, _12161_);
  or (_30976_, _30975_, _12116_);
  and (_30977_, _30976_, _05498_);
  or (_30978_, _30977_, _30890_);
  and (_30979_, _30978_, _03455_);
  or (_30980_, _30979_, _03903_);
  or (_30981_, _30980_, _30961_);
  and (_30983_, _30981_, _30900_);
  or (_30984_, _30983_, _03897_);
  nand (_30985_, _11126_, _04382_);
  nor (_30986_, _11126_, _04382_);
  not (_30987_, _30986_);
  and (_30988_, _30987_, _30985_);
  and (_30989_, _30988_, _05498_);
  or (_30990_, _30890_, _04790_);
  or (_30991_, _30990_, _30989_);
  and (_30992_, _30991_, _04792_);
  and (_30994_, _30992_, _30984_);
  or (_30995_, _30994_, _30897_);
  and (_30996_, _30995_, _03909_);
  nand (_30997_, _30899_, _03908_);
  nor (_30998_, _30997_, _30901_);
  or (_30999_, _30998_, _30996_);
  and (_31000_, _30999_, _04785_);
  not (_31001_, _11126_);
  or (_31002_, _30890_, _31001_);
  and (_31003_, _30906_, _04027_);
  and (_31005_, _31003_, _31002_);
  or (_31006_, _31005_, _03914_);
  or (_31007_, _31006_, _31000_);
  and (_31008_, _30985_, _05498_);
  or (_31009_, _30890_, _06567_);
  or (_31010_, _31009_, _31008_);
  and (_31011_, _31010_, _06572_);
  and (_31012_, _31011_, _31007_);
  and (_31013_, _30891_, _05498_);
  or (_31014_, _31013_, _30890_);
  and (_31016_, _31014_, _04011_);
  or (_31017_, _31016_, _03773_);
  or (_31018_, _31017_, _31012_);
  or (_31019_, _30902_, _03774_);
  and (_31020_, _31019_, _03375_);
  and (_31021_, _31020_, _31018_);
  and (_31022_, _30890_, _03374_);
  or (_31023_, _31022_, _03772_);
  or (_31024_, _31023_, _31021_);
  or (_31025_, _30902_, _04060_);
  and (_31026_, _31025_, _43152_);
  and (_31027_, _31026_, _31024_);
  or (_43528_, _31027_, _30888_);
  and (_31028_, _11115_, _04595_);
  nor (_31029_, _11115_, _04595_);
  nor (_31030_, _31029_, _31028_);
  or (_31031_, _31030_, _30889_);
  or (_31032_, _05498_, \oc8051_golden_model_1.P2 [1]);
  and (_31033_, _31032_, _03897_);
  and (_31034_, _31033_, _31031_);
  nor (_31037_, _11241_, _11127_);
  and (_31038_, _31037_, _05498_);
  not (_31039_, _31038_);
  and (_31040_, _31039_, _31032_);
  or (_31041_, _31040_, _04722_);
  nand (_31042_, _05498_, _03474_);
  and (_31043_, _31042_, _31032_);
  and (_31044_, _31043_, _04707_);
  and (_31045_, _04708_, \oc8051_golden_model_1.P2 [1]);
  or (_31046_, _31045_, _03850_);
  or (_31048_, _31046_, _31044_);
  and (_31049_, _31048_, _03764_);
  and (_31050_, _31049_, _31041_);
  and (_31051_, _06112_, \oc8051_golden_model_1.P0 [1]);
  and (_31052_, _06106_, \oc8051_golden_model_1.P2 [1]);
  nor (_31053_, _31052_, _31051_);
  and (_31054_, _06114_, \oc8051_golden_model_1.P1 [1]);
  and (_31055_, _06108_, \oc8051_golden_model_1.P3 [1]);
  nor (_31056_, _31055_, _31054_);
  and (_31057_, _31056_, _31053_);
  and (_31059_, _31057_, _10755_);
  and (_31060_, _31059_, _10752_);
  and (_31061_, _31060_, _10742_);
  nand (_31062_, _31061_, _10741_);
  and (_31063_, _31062_, _06106_);
  and (_31064_, _30913_, \oc8051_golden_model_1.P2 [1]);
  or (_31065_, _31064_, _31063_);
  and (_31066_, _31065_, _03763_);
  or (_31067_, _31066_, _03848_);
  or (_31068_, _31067_, _31050_);
  and (_31070_, _30889_, \oc8051_golden_model_1.P2 [1]);
  and (_31071_, _05498_, _04900_);
  or (_31072_, _31071_, _31070_);
  or (_31073_, _31072_, _04733_);
  and (_31074_, _31073_, _31068_);
  or (_31075_, _31074_, _03854_);
  or (_31076_, _31043_, _03855_);
  and (_31077_, _31076_, _03760_);
  and (_31078_, _31077_, _31075_);
  nor (_31079_, _31061_, _10740_);
  and (_31081_, _31079_, _06106_);
  or (_31082_, _31081_, _31064_);
  and (_31083_, _31082_, _03759_);
  or (_31084_, _31083_, _31078_);
  nor (_31085_, _03752_, _03746_);
  and (_31086_, _31085_, _31084_);
  or (_31087_, _31061_, _10741_);
  and (_31088_, _31063_, _03747_);
  and (_31089_, _31088_, _31087_);
  or (_31090_, _31089_, _31064_);
  and (_31092_, _31090_, _03752_);
  or (_31093_, _31079_, _12292_);
  and (_31094_, _31093_, _06106_);
  or (_31095_, _31094_, _31064_);
  and (_31096_, _31095_, _03746_);
  or (_31097_, _31096_, _07927_);
  or (_31098_, _31097_, _31092_);
  or (_31099_, _31098_, _31086_);
  and (_31100_, _06961_, _05498_);
  or (_31101_, _31070_, _03738_);
  or (_31103_, _31101_, _31100_);
  or (_31104_, _31072_, _07925_);
  and (_31105_, _31104_, _03820_);
  and (_31106_, _31105_, _31103_);
  and (_31107_, _31106_, _31099_);
  and (_31108_, _06505_, \oc8051_golden_model_1.P1 [1]);
  and (_31109_, _06507_, \oc8051_golden_model_1.P3 [1]);
  or (_31110_, _31109_, _31108_);
  or (_31111_, _31110_, _12329_);
  and (_31112_, _06501_, \oc8051_golden_model_1.P0 [1]);
  and (_31114_, _06515_, \oc8051_golden_model_1.P2 [1]);
  or (_31115_, _31114_, _31112_);
  nor (_31116_, _31115_, _31111_);
  and (_31117_, _31116_, _12347_);
  and (_31118_, _31117_, _12328_);
  nand (_31119_, _31118_, _12321_);
  or (_31120_, _31119_, _12305_);
  and (_31121_, _31120_, _05498_);
  or (_31122_, _31121_, _31070_);
  and (_31123_, _31122_, _03455_);
  or (_31125_, _31123_, _31107_);
  and (_31126_, _31125_, _04778_);
  nand (_31127_, _05498_, _04595_);
  and (_31128_, _31032_, _03903_);
  and (_31129_, _31128_, _31127_);
  or (_31130_, _31129_, _31126_);
  and (_31131_, _31130_, _04790_);
  or (_31132_, _31131_, _31034_);
  and (_31133_, _31132_, _04792_);
  nand (_31134_, _11115_, _03474_);
  or (_31136_, _11115_, _03474_);
  and (_31137_, _31136_, _31134_);
  or (_31138_, _31137_, _30889_);
  and (_31139_, _31032_, _04018_);
  and (_31140_, _31139_, _31138_);
  or (_31141_, _31140_, _31133_);
  and (_31142_, _31141_, _03909_);
  or (_31143_, _31029_, _30889_);
  and (_31144_, _31032_, _03908_);
  and (_31145_, _31144_, _31143_);
  or (_31147_, _31145_, _31142_);
  and (_31148_, _31147_, _04785_);
  not (_31149_, _11115_);
  or (_31150_, _31070_, _31149_);
  and (_31151_, _31043_, _04027_);
  and (_31152_, _31151_, _31150_);
  or (_31153_, _31152_, _31148_);
  and (_31154_, _31153_, _04012_);
  or (_31155_, _31127_, _31149_);
  and (_31156_, _31032_, _03914_);
  and (_31158_, _31156_, _31155_);
  or (_31159_, _31134_, _30889_);
  and (_31160_, _31032_, _04011_);
  and (_31161_, _31160_, _31159_);
  or (_31162_, _31161_, _03773_);
  or (_31163_, _31162_, _31158_);
  or (_31164_, _31163_, _31154_);
  or (_31165_, _31040_, _03774_);
  and (_31166_, _31165_, _03375_);
  and (_31167_, _31166_, _31164_);
  and (_31169_, _31082_, _03374_);
  or (_31170_, _31169_, _03772_);
  or (_31171_, _31170_, _31167_);
  or (_31172_, _31070_, _04060_);
  or (_31173_, _31172_, _31038_);
  and (_31174_, _31173_, _43152_);
  and (_31175_, _31174_, _31171_);
  nor (_31176_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_31177_, _31176_, _05397_);
  or (_43529_, _31177_, _31175_);
  and (_31179_, _30889_, \oc8051_golden_model_1.P2 [2]);
  nand (_31180_, _11103_, _07190_);
  or (_31181_, _11103_, _07190_);
  and (_31182_, _31181_, _31180_);
  and (_31183_, _31182_, _05498_);
  or (_31184_, _31183_, _31179_);
  and (_31185_, _31184_, _04018_);
  and (_31186_, _05498_, _06495_);
  or (_31187_, _31186_, _31179_);
  or (_31188_, _31187_, _04778_);
  and (_31190_, _05498_, _05307_);
  or (_31191_, _31190_, _31179_);
  or (_31192_, _31191_, _04733_);
  nor (_31193_, _11127_, _11103_);
  or (_31194_, _31193_, _11128_);
  and (_31195_, _31194_, _05498_);
  or (_31196_, _31195_, _31179_);
  or (_31197_, _31196_, _04722_);
  and (_31198_, _05498_, \oc8051_golden_model_1.ACC [2]);
  or (_31199_, _31198_, _31179_);
  and (_31201_, _31199_, _04707_);
  and (_31202_, _04708_, \oc8051_golden_model_1.P2 [2]);
  or (_31203_, _31202_, _03850_);
  or (_31204_, _31203_, _31201_);
  and (_31205_, _31204_, _03764_);
  and (_31206_, _31205_, _31197_);
  and (_31207_, _30913_, \oc8051_golden_model_1.P2 [2]);
  and (_31208_, _06112_, \oc8051_golden_model_1.P0 [2]);
  and (_31209_, _06106_, \oc8051_golden_model_1.P2 [2]);
  nor (_31210_, _31209_, _31208_);
  and (_31212_, _06114_, \oc8051_golden_model_1.P1 [2]);
  and (_31213_, _06108_, \oc8051_golden_model_1.P3 [2]);
  nor (_31214_, _31213_, _31212_);
  and (_31215_, _31214_, _31210_);
  and (_31216_, _31215_, _10726_);
  and (_31217_, _31216_, _10723_);
  and (_31218_, _31217_, _10713_);
  nand (_31219_, _31218_, _10738_);
  and (_31220_, _31219_, _06106_);
  or (_31221_, _31220_, _31207_);
  and (_31223_, _31221_, _03763_);
  or (_31224_, _31223_, _03848_);
  or (_31225_, _31224_, _31206_);
  and (_31226_, _31225_, _31192_);
  or (_31227_, _31226_, _03854_);
  or (_31228_, _31199_, _03855_);
  and (_31229_, _31228_, _03760_);
  and (_31230_, _31229_, _31227_);
  nor (_31231_, _31218_, _10737_);
  and (_31232_, _31231_, _06106_);
  or (_31234_, _31232_, _31207_);
  and (_31235_, _31234_, _03759_);
  or (_31236_, _31235_, _03752_);
  or (_31237_, _31236_, _31230_);
  or (_31238_, _31218_, _10738_);
  and (_31239_, _31220_, _31238_);
  or (_31240_, _31207_, _03753_);
  or (_31241_, _31240_, _31239_);
  and (_31242_, _31241_, _03747_);
  and (_31243_, _31242_, _31237_);
  or (_31245_, _31231_, _12513_);
  and (_31246_, _31245_, _06106_);
  or (_31247_, _31246_, _31207_);
  and (_31248_, _31247_, _03746_);
  or (_31249_, _31248_, _07927_);
  or (_31250_, _31249_, _31243_);
  and (_31251_, _06965_, _05498_);
  or (_31252_, _31179_, _03738_);
  or (_31253_, _31252_, _31251_);
  or (_31254_, _31191_, _07925_);
  and (_31256_, _31254_, _03820_);
  and (_31257_, _31256_, _31253_);
  and (_31258_, _31257_, _31250_);
  and (_31259_, _06501_, \oc8051_golden_model_1.P0 [2]);
  and (_31260_, _06515_, \oc8051_golden_model_1.P2 [2]);
  or (_31261_, _31260_, _12532_);
  or (_31262_, _31261_, _31259_);
  and (_31263_, _06505_, \oc8051_golden_model_1.P1 [2]);
  and (_31264_, _06507_, \oc8051_golden_model_1.P3 [2]);
  or (_31265_, _31264_, _31263_);
  nor (_31267_, _31265_, _12533_);
  nand (_31268_, _31267_, _12541_);
  nor (_31269_, _31268_, _31262_);
  and (_31270_, _31269_, _12529_);
  nand (_31271_, _31270_, _12569_);
  or (_31272_, _31271_, _12526_);
  and (_31273_, _31272_, _05498_);
  or (_31274_, _31273_, _31179_);
  and (_31275_, _31274_, _03455_);
  or (_31276_, _31275_, _03903_);
  or (_31278_, _31276_, _31258_);
  and (_31279_, _31278_, _31188_);
  or (_31280_, _31279_, _03897_);
  nand (_31281_, _11103_, _04180_);
  or (_31282_, _11103_, _04180_);
  and (_31283_, _31282_, _31281_);
  and (_31284_, _31283_, _05498_);
  or (_31285_, _31179_, _04790_);
  or (_31286_, _31285_, _31284_);
  and (_31287_, _31286_, _04792_);
  and (_31289_, _31287_, _31280_);
  or (_31290_, _31289_, _31185_);
  and (_31291_, _31290_, _03909_);
  or (_31292_, _31179_, _11240_);
  and (_31293_, _31187_, _03908_);
  and (_31294_, _31293_, _31292_);
  or (_31295_, _31294_, _31291_);
  and (_31296_, _31295_, _04785_);
  and (_31297_, _31199_, _04027_);
  and (_31298_, _31297_, _31292_);
  or (_31300_, _31298_, _03914_);
  or (_31301_, _31300_, _31296_);
  and (_31302_, _31281_, _05498_);
  or (_31303_, _31179_, _06567_);
  or (_31304_, _31303_, _31302_);
  and (_31305_, _31304_, _06572_);
  and (_31306_, _31305_, _31301_);
  and (_31307_, _31180_, _05498_);
  or (_31308_, _31307_, _31179_);
  and (_31309_, _31308_, _04011_);
  or (_31311_, _31309_, _03773_);
  or (_31312_, _31311_, _31306_);
  or (_31313_, _31196_, _03774_);
  and (_31314_, _31313_, _03375_);
  and (_31315_, _31314_, _31312_);
  and (_31316_, _31234_, _03374_);
  or (_31317_, _31316_, _03772_);
  or (_31318_, _31317_, _31315_);
  nor (_31319_, _11241_, _11240_);
  nor (_31320_, _31319_, _11242_);
  and (_31321_, _31320_, _05498_);
  or (_31322_, _31179_, _04060_);
  or (_31323_, _31322_, _31321_);
  and (_31324_, _31323_, _43152_);
  and (_31325_, _31324_, _31318_);
  nor (_31326_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_31327_, _31326_, _05397_);
  or (_43530_, _31327_, _31325_);
  and (_31328_, _30889_, \oc8051_golden_model_1.P2 [3]);
  nand (_31329_, _11087_, _07184_);
  or (_31331_, _11087_, _07184_);
  and (_31332_, _31331_, _31329_);
  and (_31333_, _31332_, _05498_);
  or (_31334_, _31333_, _31328_);
  and (_31335_, _31334_, _04018_);
  and (_31336_, _05498_, _06345_);
  or (_31337_, _31336_, _31328_);
  or (_31338_, _31337_, _04778_);
  nor (_31339_, _11128_, _11087_);
  or (_31340_, _31339_, _11129_);
  and (_31342_, _31340_, _05498_);
  or (_31343_, _31342_, _31328_);
  or (_31344_, _31343_, _04722_);
  and (_31345_, _05498_, \oc8051_golden_model_1.ACC [3]);
  or (_31346_, _31345_, _31328_);
  and (_31347_, _31346_, _04707_);
  and (_31348_, _04708_, \oc8051_golden_model_1.P2 [3]);
  or (_31349_, _31348_, _03850_);
  or (_31350_, _31349_, _31347_);
  and (_31351_, _31350_, _03764_);
  and (_31353_, _31351_, _31344_);
  and (_31354_, _30913_, \oc8051_golden_model_1.P2 [3]);
  and (_31355_, _06112_, \oc8051_golden_model_1.P0 [3]);
  and (_31356_, _06106_, \oc8051_golden_model_1.P2 [3]);
  nor (_31357_, _31356_, _31355_);
  and (_31358_, _06114_, \oc8051_golden_model_1.P1 [3]);
  and (_31359_, _06108_, \oc8051_golden_model_1.P3 [3]);
  nor (_31360_, _31359_, _31358_);
  and (_31361_, _31360_, _31357_);
  and (_31362_, _31361_, _10863_);
  and (_31364_, _31362_, _10860_);
  and (_31365_, _31364_, _10850_);
  nand (_31366_, _31365_, _10875_);
  and (_31367_, _31366_, _06106_);
  or (_31368_, _31367_, _31354_);
  and (_31369_, _31368_, _03763_);
  or (_31370_, _31369_, _03848_);
  or (_31371_, _31370_, _31353_);
  and (_31372_, _05498_, _05119_);
  or (_31373_, _31372_, _31328_);
  or (_31375_, _31373_, _04733_);
  and (_31376_, _31375_, _31371_);
  or (_31377_, _31376_, _03854_);
  or (_31378_, _31346_, _03855_);
  and (_31379_, _31378_, _03760_);
  and (_31380_, _31379_, _31377_);
  nor (_31381_, _31365_, _10874_);
  and (_31382_, _31381_, _06106_);
  or (_31383_, _31382_, _31354_);
  and (_31384_, _31383_, _03759_);
  or (_31386_, _31384_, _03752_);
  or (_31387_, _31386_, _31380_);
  or (_31388_, _31365_, _10875_);
  or (_31389_, _31354_, _31388_);
  and (_31390_, _31389_, _31368_);
  or (_31391_, _31390_, _03753_);
  and (_31392_, _31391_, _03747_);
  and (_31393_, _31392_, _31387_);
  or (_31394_, _31381_, _12666_);
  and (_31395_, _31394_, _06106_);
  or (_31397_, _31395_, _31354_);
  and (_31398_, _31397_, _03746_);
  or (_31399_, _31398_, _07927_);
  or (_31400_, _31399_, _31393_);
  and (_31401_, _06964_, _05498_);
  or (_31402_, _31328_, _03738_);
  or (_31403_, _31402_, _31401_);
  or (_31404_, _31373_, _07925_);
  and (_31405_, _31404_, _03820_);
  and (_31406_, _31405_, _31403_);
  and (_31408_, _31406_, _31400_);
  and (_31409_, _06501_, \oc8051_golden_model_1.P0 [3]);
  and (_31410_, _06515_, \oc8051_golden_model_1.P2 [3]);
  or (_31411_, _31410_, _31409_);
  and (_31412_, _06505_, \oc8051_golden_model_1.P1 [3]);
  and (_31413_, _06507_, \oc8051_golden_model_1.P3 [3]);
  or (_31414_, _31413_, _31412_);
  or (_31415_, _31414_, _12758_);
  nor (_31416_, _31415_, _31411_);
  and (_31417_, _31416_, _12770_);
  and (_31419_, _31417_, _12751_);
  nand (_31420_, _31419_, _12744_);
  or (_31421_, _31420_, _12729_);
  and (_31422_, _31421_, _05498_);
  or (_31423_, _31422_, _31328_);
  and (_31424_, _31423_, _03455_);
  or (_31425_, _31424_, _03903_);
  or (_31426_, _31425_, _31408_);
  and (_31427_, _31426_, _31338_);
  or (_31428_, _31427_, _03897_);
  nand (_31430_, _11087_, _04005_);
  or (_31431_, _11087_, _04005_);
  and (_31432_, _31431_, _31430_);
  and (_31433_, _31432_, _05498_);
  or (_31434_, _31328_, _04790_);
  or (_31435_, _31434_, _31433_);
  and (_31436_, _31435_, _04792_);
  and (_31437_, _31436_, _31428_);
  or (_31438_, _31437_, _31335_);
  and (_31439_, _31438_, _03909_);
  or (_31441_, _31328_, _11239_);
  and (_31442_, _31337_, _03908_);
  and (_31443_, _31442_, _31441_);
  or (_31444_, _31443_, _31439_);
  and (_31445_, _31444_, _04785_);
  and (_31446_, _31346_, _04027_);
  and (_31447_, _31446_, _31441_);
  or (_31448_, _31447_, _03914_);
  or (_31449_, _31448_, _31445_);
  and (_31450_, _31430_, _05498_);
  or (_31452_, _31328_, _06567_);
  or (_31453_, _31452_, _31450_);
  and (_31454_, _31453_, _06572_);
  and (_31455_, _31454_, _31449_);
  and (_31456_, _31329_, _05498_);
  or (_31457_, _31456_, _31328_);
  and (_31458_, _31457_, _04011_);
  or (_31459_, _31458_, _03773_);
  or (_31460_, _31459_, _31455_);
  or (_31461_, _31343_, _03774_);
  and (_31463_, _31461_, _03375_);
  and (_31464_, _31463_, _31460_);
  and (_31465_, _31383_, _03374_);
  or (_31466_, _31465_, _03772_);
  or (_31467_, _31466_, _31464_);
  nor (_31468_, _11242_, _11239_);
  nor (_31469_, _31468_, _11243_);
  and (_31470_, _31469_, _05498_);
  or (_31471_, _31328_, _04060_);
  or (_31472_, _31471_, _31470_);
  and (_31474_, _31472_, _43152_);
  and (_31475_, _31474_, _31467_);
  nor (_31476_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_31477_, _31476_, _05397_);
  or (_43531_, _31477_, _31475_);
  nor (_31478_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_31479_, _31478_, _05397_);
  and (_31480_, _30889_, \oc8051_golden_model_1.P2 [4]);
  nand (_31481_, _11076_, _07090_);
  or (_31482_, _11076_, _07090_);
  and (_31484_, _31482_, _31481_);
  and (_31485_, _31484_, _05498_);
  or (_31486_, _31485_, _31480_);
  and (_31487_, _31486_, _04018_);
  and (_31488_, _06456_, _05498_);
  or (_31489_, _31488_, _31480_);
  or (_31490_, _31489_, _04778_);
  nor (_31491_, _11129_, _11076_);
  or (_31492_, _31491_, _11130_);
  and (_31493_, _31492_, _05498_);
  or (_31495_, _31493_, _31480_);
  or (_31496_, _31495_, _04722_);
  and (_31497_, _05498_, \oc8051_golden_model_1.ACC [4]);
  or (_31498_, _31497_, _31480_);
  and (_31499_, _31498_, _04707_);
  and (_31500_, _04708_, \oc8051_golden_model_1.P2 [4]);
  or (_31501_, _31500_, _03850_);
  or (_31502_, _31501_, _31499_);
  and (_31503_, _31502_, _03764_);
  and (_31504_, _31503_, _31496_);
  and (_31506_, _30913_, \oc8051_golden_model_1.P2 [4]);
  and (_31507_, _06108_, \oc8051_golden_model_1.P3 [4]);
  nor (_31508_, _31507_, _10776_);
  and (_31509_, _31508_, _10783_);
  and (_31510_, _06114_, \oc8051_golden_model_1.P1 [4]);
  not (_31511_, _31510_);
  and (_31512_, _06112_, \oc8051_golden_model_1.P0 [4]);
  and (_31513_, _06106_, \oc8051_golden_model_1.P2 [4]);
  nor (_31514_, _31513_, _31512_);
  and (_31515_, _31514_, _31511_);
  and (_31517_, _31515_, _10775_);
  and (_31518_, _31517_, _31509_);
  and (_31519_, _31518_, _10768_);
  nand (_31520_, _31519_, _10792_);
  and (_31521_, _31520_, _06106_);
  or (_31522_, _31521_, _31506_);
  and (_31523_, _31522_, _03763_);
  or (_31524_, _31523_, _03848_);
  or (_31525_, _31524_, _31504_);
  and (_31526_, _05950_, _05498_);
  or (_31528_, _31526_, _31480_);
  or (_31529_, _31528_, _04733_);
  and (_31530_, _31529_, _31525_);
  or (_31531_, _31530_, _03854_);
  or (_31532_, _31498_, _03855_);
  and (_31533_, _31532_, _03760_);
  and (_31534_, _31533_, _31531_);
  nor (_31535_, _31519_, _10791_);
  and (_31536_, _31535_, _06106_);
  or (_31537_, _31536_, _31506_);
  and (_31539_, _31537_, _03759_);
  or (_31540_, _31539_, _03752_);
  or (_31541_, _31540_, _31534_);
  or (_31542_, _31519_, _10792_);
  or (_31543_, _31506_, _31542_);
  and (_31544_, _31543_, _31522_);
  or (_31545_, _31544_, _03753_);
  and (_31546_, _31545_, _03747_);
  and (_31547_, _31546_, _31541_);
  or (_31548_, _31535_, _12871_);
  and (_31550_, _31548_, _06106_);
  or (_31551_, _31550_, _31506_);
  and (_31552_, _31551_, _03746_);
  or (_31553_, _31552_, _07927_);
  or (_31554_, _31553_, _31547_);
  and (_31555_, _06969_, _05498_);
  or (_31556_, _31480_, _03738_);
  or (_31557_, _31556_, _31555_);
  or (_31558_, _31528_, _07925_);
  and (_31559_, _31558_, _03820_);
  and (_31561_, _31559_, _31557_);
  and (_31562_, _31561_, _31554_);
  and (_31563_, _06501_, \oc8051_golden_model_1.P0 [4]);
  and (_31564_, _06515_, \oc8051_golden_model_1.P2 [4]);
  or (_31565_, _31564_, _12947_);
  nor (_31566_, _31565_, _31563_);
  and (_31567_, _31566_, _12944_);
  nand (_31568_, _31567_, _12937_);
  and (_31569_, _06505_, \oc8051_golden_model_1.P1 [4]);
  and (_31570_, _06507_, \oc8051_golden_model_1.P3 [4]);
  or (_31572_, _31570_, _31569_);
  or (_31573_, _31572_, _12948_);
  nor (_31574_, _31573_, _12960_);
  and (_31575_, _31574_, _12977_);
  nand (_31576_, _31575_, _12959_);
  or (_31577_, _31576_, _31568_);
  or (_31578_, _31577_, _12934_);
  and (_31579_, _31578_, _05498_);
  or (_31580_, _31579_, _31480_);
  and (_31581_, _31580_, _03455_);
  or (_31583_, _31581_, _03903_);
  or (_31584_, _31583_, _31562_);
  and (_31585_, _31584_, _31490_);
  or (_31586_, _31585_, _03897_);
  nand (_31587_, _11076_, _06442_);
  or (_31588_, _11076_, _06442_);
  and (_31589_, _31588_, _31587_);
  and (_31590_, _31589_, _05498_);
  or (_31591_, _31590_, _31480_);
  or (_31592_, _31591_, _04790_);
  and (_31594_, _31592_, _04792_);
  and (_31595_, _31594_, _31586_);
  or (_31596_, _31595_, _31487_);
  and (_31597_, _31596_, _03909_);
  or (_31598_, _31480_, _11238_);
  and (_31599_, _31489_, _03908_);
  and (_31600_, _31599_, _31598_);
  or (_31601_, _31600_, _31597_);
  and (_31602_, _31601_, _04785_);
  and (_31603_, _31498_, _04027_);
  and (_31604_, _31603_, _31598_);
  or (_31605_, _31604_, _03914_);
  or (_31606_, _31605_, _31602_);
  and (_31607_, _31587_, _05498_);
  or (_31608_, _31480_, _06567_);
  or (_31609_, _31608_, _31607_);
  and (_31610_, _31609_, _06572_);
  and (_31611_, _31610_, _31606_);
  and (_31612_, _31481_, _05498_);
  or (_31613_, _31612_, _31480_);
  and (_31616_, _31613_, _04011_);
  or (_31617_, _31616_, _03773_);
  or (_31618_, _31617_, _31611_);
  or (_31619_, _31495_, _03774_);
  and (_31620_, _31619_, _03375_);
  and (_31621_, _31620_, _31618_);
  and (_31622_, _31537_, _03374_);
  or (_31623_, _31622_, _03772_);
  or (_31624_, _31623_, _31621_);
  nor (_31625_, _11243_, _11238_);
  nor (_31627_, _31625_, _11244_);
  and (_31628_, _31627_, _05498_);
  or (_31629_, _31480_, _04060_);
  or (_31630_, _31629_, _31628_);
  and (_31631_, _31630_, _43152_);
  and (_31632_, _31631_, _31624_);
  or (_43532_, _31632_, _31479_);
  and (_31633_, _30889_, \oc8051_golden_model_1.P2 [5]);
  nand (_31634_, _11060_, _07084_);
  or (_31635_, _11060_, _07084_);
  and (_31637_, _31635_, _31634_);
  and (_31638_, _31637_, _05498_);
  or (_31639_, _31638_, _31633_);
  and (_31640_, _31639_, _04018_);
  and (_31641_, _06447_, _05498_);
  or (_31642_, _31641_, _31633_);
  or (_31643_, _31642_, _04778_);
  nor (_31644_, _11130_, _11060_);
  or (_31645_, _31644_, _11131_);
  and (_31646_, _31645_, _05498_);
  or (_31648_, _31646_, _31633_);
  or (_31649_, _31648_, _04722_);
  and (_31650_, _05498_, \oc8051_golden_model_1.ACC [5]);
  or (_31651_, _31650_, _31633_);
  and (_31652_, _31651_, _04707_);
  and (_31653_, _04708_, \oc8051_golden_model_1.P2 [5]);
  or (_31654_, _31653_, _03850_);
  or (_31655_, _31654_, _31652_);
  and (_31656_, _31655_, _03764_);
  and (_31657_, _31656_, _31649_);
  and (_31659_, _30913_, \oc8051_golden_model_1.P2 [5]);
  and (_31660_, _06112_, \oc8051_golden_model_1.P0 [5]);
  and (_31661_, _06106_, \oc8051_golden_model_1.P2 [5]);
  nor (_31662_, _31661_, _31660_);
  and (_31663_, _06114_, \oc8051_golden_model_1.P1 [5]);
  and (_31664_, _06108_, \oc8051_golden_model_1.P3 [5]);
  nor (_31665_, _31664_, _31663_);
  and (_31666_, _31665_, _31662_);
  and (_31667_, _31666_, _10890_);
  and (_31668_, _31667_, _10887_);
  and (_31670_, _31668_, _10877_);
  nand (_31671_, _31670_, _10902_);
  and (_31672_, _31671_, _06106_);
  or (_31673_, _31672_, _31659_);
  and (_31674_, _31673_, _03763_);
  or (_31675_, _31674_, _03848_);
  or (_31676_, _31675_, _31657_);
  and (_31677_, _05857_, _05498_);
  or (_31678_, _31677_, _31633_);
  or (_31679_, _31678_, _04733_);
  and (_31681_, _31679_, _31676_);
  or (_31682_, _31681_, _03854_);
  or (_31683_, _31651_, _03855_);
  and (_31684_, _31683_, _03760_);
  and (_31685_, _31684_, _31682_);
  nor (_31686_, _31670_, _10901_);
  and (_31687_, _31686_, _06106_);
  or (_31688_, _31687_, _31659_);
  and (_31689_, _31688_, _03759_);
  or (_31690_, _31689_, _03752_);
  or (_31692_, _31690_, _31685_);
  or (_31693_, _31670_, _10902_);
  or (_31694_, _31659_, _31693_);
  and (_31695_, _31694_, _31673_);
  or (_31696_, _31695_, _03753_);
  and (_31697_, _31696_, _03747_);
  and (_31698_, _31697_, _31692_);
  or (_31699_, _31686_, _13072_);
  and (_31700_, _31699_, _06106_);
  or (_31701_, _31700_, _31659_);
  and (_31703_, _31701_, _03746_);
  or (_31704_, _31703_, _07927_);
  or (_31705_, _31704_, _31698_);
  and (_31706_, _06968_, _05498_);
  or (_31707_, _31633_, _03738_);
  or (_31708_, _31707_, _31706_);
  or (_31709_, _31678_, _07925_);
  and (_31710_, _31709_, _03820_);
  and (_31711_, _31710_, _31708_);
  and (_31712_, _31711_, _31705_);
  and (_31714_, _06515_, \oc8051_golden_model_1.P2 [5]);
  and (_31715_, _06501_, \oc8051_golden_model_1.P0 [5]);
  or (_31716_, _31715_, _13142_);
  or (_31717_, _31716_, _31714_);
  and (_31718_, _06505_, \oc8051_golden_model_1.P1 [5]);
  and (_31719_, _06507_, \oc8051_golden_model_1.P3 [5]);
  or (_31720_, _31719_, _31718_);
  nor (_31721_, _31720_, _13143_);
  nand (_31722_, _31721_, _13151_);
  nor (_31723_, _31722_, _31717_);
  and (_31725_, _31723_, _13139_);
  nand (_31726_, _31725_, _13179_);
  or (_31727_, _31726_, _13136_);
  and (_31728_, _31727_, _05498_);
  or (_31729_, _31728_, _31633_);
  and (_31730_, _31729_, _03455_);
  or (_31731_, _31730_, _03903_);
  or (_31732_, _31731_, _31712_);
  and (_31733_, _31732_, _31643_);
  or (_31734_, _31733_, _03897_);
  nand (_31736_, _11060_, _06411_);
  or (_31737_, _11060_, _06411_);
  and (_31738_, _31737_, _31736_);
  and (_31739_, _31738_, _05498_);
  or (_31740_, _31633_, _04790_);
  or (_31741_, _31740_, _31739_);
  and (_31742_, _31741_, _04792_);
  and (_31743_, _31742_, _31734_);
  or (_31744_, _31743_, _31640_);
  and (_31745_, _31744_, _03909_);
  or (_31747_, _31633_, _11237_);
  and (_31748_, _31642_, _03908_);
  and (_31749_, _31748_, _31747_);
  or (_31750_, _31749_, _31745_);
  and (_31751_, _31750_, _04785_);
  and (_31752_, _31651_, _04027_);
  and (_31753_, _31752_, _31747_);
  or (_31754_, _31753_, _03914_);
  or (_31755_, _31754_, _31751_);
  and (_31756_, _31736_, _05498_);
  or (_31758_, _31633_, _06567_);
  or (_31759_, _31758_, _31756_);
  and (_31760_, _31759_, _06572_);
  and (_31761_, _31760_, _31755_);
  and (_31762_, _31634_, _05498_);
  or (_31763_, _31762_, _31633_);
  and (_31764_, _31763_, _04011_);
  or (_31765_, _31764_, _03773_);
  or (_31766_, _31765_, _31761_);
  or (_31767_, _31648_, _03774_);
  and (_31769_, _31767_, _03375_);
  and (_31770_, _31769_, _31766_);
  and (_31771_, _31688_, _03374_);
  or (_31772_, _31771_, _03772_);
  or (_31773_, _31772_, _31770_);
  nor (_31774_, _11244_, _11237_);
  nor (_31775_, _31774_, _11245_);
  and (_31776_, _31775_, _05498_);
  or (_31777_, _31633_, _04060_);
  or (_31778_, _31777_, _31776_);
  and (_31780_, _31778_, _43152_);
  and (_31781_, _31780_, _31773_);
  nor (_31782_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_31783_, _31782_, _05397_);
  or (_43533_, _31783_, _31781_);
  and (_31784_, _30889_, \oc8051_golden_model_1.P2 [6]);
  nand (_31785_, _11044_, _07036_);
  or (_31786_, _11044_, _07036_);
  and (_31787_, _31786_, _31785_);
  and (_31788_, _31787_, _05498_);
  or (_31790_, _31788_, _31784_);
  and (_31791_, _31790_, _04018_);
  and (_31792_, _13394_, _05498_);
  or (_31793_, _31792_, _31784_);
  or (_31794_, _31793_, _04778_);
  and (_31795_, _30913_, \oc8051_golden_model_1.P2 [6]);
  and (_31796_, _06112_, \oc8051_golden_model_1.P0 [6]);
  and (_31797_, _06106_, \oc8051_golden_model_1.P2 [6]);
  nor (_31798_, _31797_, _31796_);
  and (_31799_, _06114_, \oc8051_golden_model_1.P1 [6]);
  and (_31801_, _06108_, \oc8051_golden_model_1.P3 [6]);
  nor (_31802_, _31801_, _31799_);
  and (_31803_, _31802_, _31798_);
  and (_31804_, _31803_, _10835_);
  and (_31805_, _31804_, _10832_);
  and (_31806_, _31805_, _10822_);
  nor (_31807_, _31806_, _10846_);
  and (_31808_, _31807_, _06106_);
  or (_31809_, _31808_, _31795_);
  and (_31810_, _31809_, _03759_);
  nor (_31812_, _11131_, _11044_);
  or (_31813_, _31812_, _11132_);
  and (_31814_, _31813_, _05498_);
  or (_31815_, _31814_, _31784_);
  or (_31816_, _31815_, _04722_);
  and (_31817_, _05498_, \oc8051_golden_model_1.ACC [6]);
  or (_31818_, _31817_, _31784_);
  and (_31819_, _31818_, _04707_);
  and (_31820_, _04708_, \oc8051_golden_model_1.P2 [6]);
  or (_31821_, _31820_, _03850_);
  or (_31823_, _31821_, _31819_);
  and (_31824_, _31823_, _03764_);
  and (_31825_, _31824_, _31816_);
  nand (_31826_, _31806_, _10847_);
  and (_31827_, _31826_, _06106_);
  or (_31828_, _31827_, _31795_);
  and (_31829_, _31828_, _03763_);
  or (_31830_, _31829_, _03848_);
  or (_31831_, _31830_, _31825_);
  and (_31832_, _06065_, _05498_);
  or (_31834_, _31832_, _31784_);
  or (_31835_, _31834_, _04733_);
  and (_31836_, _31835_, _31831_);
  or (_31837_, _31836_, _03854_);
  or (_31838_, _31818_, _03855_);
  and (_31839_, _31838_, _03760_);
  and (_31840_, _31839_, _31837_);
  or (_31841_, _31840_, _31810_);
  and (_31842_, _31841_, _03753_);
  or (_31843_, _31806_, _10847_);
  or (_31845_, _31795_, _31843_);
  and (_31846_, _31845_, _03752_);
  and (_31847_, _31846_, _31828_);
  or (_31848_, _31847_, _31842_);
  and (_31849_, _31848_, _03747_);
  or (_31850_, _31807_, _13278_);
  and (_31851_, _31850_, _06106_);
  or (_31852_, _31851_, _31795_);
  and (_31853_, _31852_, _03746_);
  or (_31854_, _31853_, _07927_);
  or (_31856_, _31854_, _31849_);
  and (_31857_, _06641_, _05498_);
  or (_31858_, _31784_, _03738_);
  or (_31859_, _31858_, _31857_);
  or (_31860_, _31834_, _07925_);
  and (_31861_, _31860_, _03820_);
  and (_31862_, _31861_, _31859_);
  and (_31863_, _31862_, _31856_);
  and (_31864_, _06505_, \oc8051_golden_model_1.P1 [6]);
  and (_31865_, _06507_, \oc8051_golden_model_1.P3 [6]);
  or (_31867_, _31865_, _31864_);
  or (_31868_, _31867_, _13342_);
  and (_31869_, _06501_, \oc8051_golden_model_1.P0 [6]);
  and (_31870_, _06515_, \oc8051_golden_model_1.P2 [6]);
  or (_31871_, _31870_, _31869_);
  or (_31872_, _31871_, _31868_);
  nor (_31873_, _31872_, _13340_);
  and (_31874_, _31873_, _13363_);
  nand (_31875_, _31874_, _13384_);
  or (_31876_, _31875_, _13339_);
  and (_31878_, _31876_, _05498_);
  or (_31879_, _31878_, _31784_);
  and (_31880_, _31879_, _03455_);
  or (_31881_, _31880_, _03903_);
  or (_31882_, _31881_, _31863_);
  and (_31883_, _31882_, _31794_);
  or (_31884_, _31883_, _03897_);
  nand (_31885_, _11044_, _06379_);
  or (_31886_, _11044_, _06379_);
  and (_31887_, _31886_, _31885_);
  and (_31889_, _31887_, _05498_);
  or (_31890_, _31784_, _04790_);
  or (_31891_, _31890_, _31889_);
  and (_31892_, _31891_, _04792_);
  and (_31893_, _31892_, _31884_);
  or (_31894_, _31893_, _31791_);
  and (_31895_, _31894_, _03909_);
  or (_31896_, _31784_, _11236_);
  and (_31897_, _31793_, _03908_);
  and (_31898_, _31897_, _31896_);
  or (_31900_, _31898_, _31895_);
  and (_31901_, _31900_, _04785_);
  and (_31902_, _31818_, _04027_);
  and (_31903_, _31902_, _31896_);
  or (_31904_, _31903_, _03914_);
  or (_31905_, _31904_, _31901_);
  and (_31906_, _31885_, _05498_);
  or (_31907_, _31784_, _06567_);
  or (_31908_, _31907_, _31906_);
  and (_31909_, _31908_, _06572_);
  and (_31911_, _31909_, _31905_);
  and (_31912_, _31785_, _05498_);
  or (_31913_, _31912_, _31784_);
  and (_31914_, _31913_, _04011_);
  or (_31915_, _31914_, _03773_);
  or (_31916_, _31915_, _31911_);
  or (_31917_, _31815_, _03774_);
  and (_31918_, _31917_, _03375_);
  and (_31919_, _31918_, _31916_);
  and (_31920_, _31809_, _03374_);
  or (_31922_, _31920_, _03772_);
  or (_31923_, _31922_, _31919_);
  or (_31924_, _11245_, _11236_);
  and (_31925_, _31924_, _11246_);
  and (_31926_, _31925_, _05498_);
  or (_31927_, _31784_, _04060_);
  or (_31928_, _31927_, _31926_);
  and (_31929_, _31928_, _43152_);
  and (_31930_, _31929_, _31923_);
  nor (_31931_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_31933_, _31931_, _05397_);
  or (_43534_, _31933_, _31930_);
  nor (_31934_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_31935_, _31934_, _05397_);
  and (_31936_, _11257_, \oc8051_golden_model_1.P3 [0]);
  and (_31937_, _30893_, _05500_);
  or (_31938_, _31937_, _31936_);
  and (_31939_, _31938_, _04018_);
  and (_31940_, _05500_, _06479_);
  or (_31941_, _31940_, _31936_);
  or (_31943_, _31941_, _04778_);
  and (_31944_, _11126_, _05500_);
  or (_31945_, _31944_, _31936_);
  or (_31946_, _31945_, _04722_);
  and (_31947_, _05500_, \oc8051_golden_model_1.ACC [0]);
  or (_31948_, _31947_, _31936_);
  and (_31949_, _31948_, _04707_);
  and (_31950_, _04708_, \oc8051_golden_model_1.P3 [0]);
  or (_31951_, _31950_, _03850_);
  or (_31952_, _31951_, _31949_);
  and (_31954_, _31952_, _03764_);
  and (_31955_, _31954_, _31946_);
  and (_31956_, _11265_, \oc8051_golden_model_1.P3 [0]);
  and (_31957_, _30926_, _06108_);
  or (_31958_, _31957_, _31956_);
  and (_31959_, _31958_, _03763_);
  or (_31960_, _31959_, _31955_);
  and (_31961_, _31960_, _04733_);
  and (_31962_, _05500_, _04700_);
  or (_31963_, _31962_, _31936_);
  and (_31965_, _31963_, _03848_);
  or (_31966_, _31965_, _03854_);
  or (_31967_, _31966_, _31961_);
  or (_31968_, _31948_, _03855_);
  and (_31969_, _31968_, _03760_);
  and (_31970_, _31969_, _31967_);
  and (_31971_, _31936_, _03759_);
  or (_31972_, _31971_, _03752_);
  or (_31973_, _31972_, _31970_);
  or (_31974_, _31945_, _03753_);
  and (_31976_, _31974_, _03747_);
  and (_31977_, _31976_, _31973_);
  or (_31978_, _31956_, _14237_);
  and (_31979_, _31978_, _03746_);
  and (_31980_, _31979_, _31958_);
  or (_31981_, _31980_, _07927_);
  or (_31982_, _31981_, _31977_);
  and (_31983_, _06962_, _05500_);
  or (_31984_, _31936_, _03738_);
  or (_31985_, _31984_, _31983_);
  or (_31987_, _31963_, _07925_);
  and (_31988_, _31987_, _03820_);
  and (_31989_, _31988_, _31985_);
  and (_31990_, _31989_, _31982_);
  and (_31991_, _30976_, _05500_);
  or (_31992_, _31991_, _31936_);
  and (_31993_, _31992_, _03455_);
  or (_31994_, _31993_, _03903_);
  or (_31995_, _31994_, _31990_);
  and (_31996_, _31995_, _31943_);
  or (_31998_, _31996_, _03897_);
  and (_31999_, _30988_, _05500_);
  or (_32000_, _31999_, _31936_);
  or (_32001_, _32000_, _04790_);
  and (_32002_, _32001_, _04792_);
  and (_32003_, _32002_, _31998_);
  or (_32004_, _32003_, _31939_);
  and (_32005_, _32004_, _03909_);
  nand (_32006_, _31941_, _03908_);
  nor (_32007_, _32006_, _31944_);
  or (_32009_, _32007_, _32005_);
  and (_32010_, _32009_, _04785_);
  or (_32011_, _31936_, _31001_);
  and (_32012_, _31948_, _04027_);
  and (_32013_, _32012_, _32011_);
  or (_32014_, _32013_, _03914_);
  or (_32015_, _32014_, _32010_);
  and (_32016_, _30985_, _05500_);
  or (_32017_, _31936_, _06567_);
  or (_32018_, _32017_, _32016_);
  and (_32020_, _32018_, _06572_);
  and (_32021_, _32020_, _32015_);
  and (_32022_, _30891_, _05500_);
  or (_32023_, _32022_, _31936_);
  and (_32024_, _32023_, _04011_);
  or (_32025_, _32024_, _03773_);
  or (_32026_, _32025_, _32021_);
  or (_32027_, _31945_, _03774_);
  and (_32028_, _32027_, _03375_);
  and (_32029_, _32028_, _32026_);
  and (_32031_, _31936_, _03374_);
  or (_32032_, _32031_, _03772_);
  or (_32033_, _32032_, _32029_);
  or (_32034_, _31945_, _04060_);
  and (_32035_, _32034_, _43152_);
  and (_32036_, _32035_, _32033_);
  or (_43535_, _32036_, _31935_);
  or (_32037_, _31030_, _11257_);
  or (_32038_, _05500_, \oc8051_golden_model_1.P3 [1]);
  and (_32039_, _32038_, _03897_);
  and (_32040_, _32039_, _32037_);
  nand (_32041_, _05500_, _04595_);
  and (_32042_, _32038_, _03903_);
  and (_32043_, _32042_, _32041_);
  and (_32044_, _31037_, _05500_);
  not (_32045_, _32044_);
  and (_32046_, _32045_, _32038_);
  or (_32047_, _32046_, _04722_);
  nand (_32048_, _05500_, _03474_);
  and (_32049_, _32048_, _32038_);
  and (_32051_, _32049_, _04707_);
  and (_32052_, _04708_, \oc8051_golden_model_1.P3 [1]);
  or (_32053_, _32052_, _03850_);
  or (_32054_, _32053_, _32051_);
  and (_32055_, _32054_, _03764_);
  and (_32056_, _32055_, _32047_);
  and (_32057_, _31062_, _06108_);
  and (_32058_, _11265_, \oc8051_golden_model_1.P3 [1]);
  or (_32059_, _32058_, _32057_);
  and (_32060_, _32059_, _03763_);
  or (_32062_, _32060_, _03848_);
  or (_32063_, _32062_, _32056_);
  and (_32064_, _11257_, \oc8051_golden_model_1.P3 [1]);
  and (_32065_, _05500_, _04900_);
  or (_32066_, _32065_, _32064_);
  or (_32067_, _32066_, _04733_);
  and (_32068_, _32067_, _32063_);
  or (_32069_, _32068_, _03854_);
  or (_32070_, _32049_, _03855_);
  and (_32071_, _32070_, _03760_);
  and (_32073_, _32071_, _32069_);
  and (_32074_, _31079_, _06108_);
  or (_32075_, _32074_, _32058_);
  and (_32076_, _32075_, _03759_);
  or (_32077_, _32076_, _32073_);
  and (_32078_, _32077_, _31085_);
  or (_32079_, _32058_, _31087_);
  and (_32080_, _32079_, _03752_);
  and (_32081_, _32080_, _32059_);
  and (_32082_, _31093_, _06108_);
  or (_32084_, _32082_, _32058_);
  and (_32085_, _32084_, _03746_);
  or (_32086_, _32085_, _07927_);
  or (_32087_, _32086_, _32081_);
  or (_32088_, _32087_, _32078_);
  and (_32089_, _06961_, _05500_);
  or (_32090_, _32064_, _03738_);
  or (_32091_, _32090_, _32089_);
  or (_32092_, _32066_, _07925_);
  and (_32093_, _32092_, _03820_);
  and (_32095_, _32093_, _32091_);
  and (_32096_, _32095_, _32088_);
  and (_32097_, _31120_, _05500_);
  or (_32098_, _32097_, _32064_);
  and (_32099_, _32098_, _03455_);
  or (_32100_, _32099_, _32096_);
  and (_32101_, _32100_, _04778_);
  or (_32102_, _32101_, _32043_);
  and (_32103_, _32102_, _04790_);
  or (_32104_, _32103_, _32040_);
  and (_32106_, _32104_, _04792_);
  or (_32107_, _31137_, _11257_);
  and (_32108_, _32038_, _04018_);
  and (_32109_, _32108_, _32107_);
  or (_32110_, _32109_, _32106_);
  and (_32111_, _32110_, _03909_);
  or (_32112_, _31029_, _11257_);
  and (_32113_, _32038_, _03908_);
  and (_32114_, _32113_, _32112_);
  or (_32115_, _32114_, _32111_);
  and (_32117_, _32115_, _04785_);
  or (_32118_, _32064_, _31149_);
  and (_32119_, _32049_, _04027_);
  and (_32120_, _32119_, _32118_);
  or (_32121_, _32120_, _32117_);
  and (_32122_, _32121_, _04012_);
  or (_32123_, _32048_, _31149_);
  and (_32124_, _32038_, _04011_);
  and (_32125_, _32124_, _32123_);
  or (_32126_, _32125_, _03773_);
  or (_32128_, _32041_, _31149_);
  and (_32129_, _32038_, _03914_);
  and (_32130_, _32129_, _32128_);
  or (_32131_, _32130_, _32126_);
  or (_32132_, _32131_, _32122_);
  or (_32133_, _32046_, _03774_);
  and (_32134_, _32133_, _03375_);
  and (_32135_, _32134_, _32132_);
  and (_32136_, _32075_, _03374_);
  or (_32137_, _32136_, _03772_);
  or (_32139_, _32137_, _32135_);
  or (_32140_, _32064_, _04060_);
  or (_32141_, _32140_, _32044_);
  and (_32142_, _32141_, _43152_);
  and (_32143_, _32142_, _32139_);
  nor (_32144_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_32145_, _32144_, _05397_);
  or (_43536_, _32145_, _32143_);
  and (_32146_, _11257_, \oc8051_golden_model_1.P3 [2]);
  and (_32147_, _31182_, _05500_);
  or (_32149_, _32147_, _32146_);
  and (_32150_, _32149_, _04018_);
  and (_32151_, _05500_, _06495_);
  or (_32152_, _32151_, _32146_);
  or (_32153_, _32152_, _04778_);
  and (_32154_, _05500_, _05307_);
  or (_32155_, _32154_, _32146_);
  or (_32156_, _32155_, _04733_);
  and (_32157_, _31194_, _05500_);
  or (_32158_, _32157_, _32146_);
  or (_32160_, _32158_, _04722_);
  and (_32161_, _05500_, \oc8051_golden_model_1.ACC [2]);
  or (_32162_, _32161_, _32146_);
  and (_32163_, _32162_, _04707_);
  and (_32164_, _04708_, \oc8051_golden_model_1.P3 [2]);
  or (_32165_, _32164_, _03850_);
  or (_32166_, _32165_, _32163_);
  and (_32167_, _32166_, _03764_);
  and (_32168_, _32167_, _32160_);
  and (_32169_, _11265_, \oc8051_golden_model_1.P3 [2]);
  and (_32171_, _31219_, _06108_);
  or (_32172_, _32171_, _32169_);
  and (_32173_, _32172_, _03763_);
  or (_32174_, _32173_, _03848_);
  or (_32175_, _32174_, _32168_);
  and (_32176_, _32175_, _32156_);
  or (_32177_, _32176_, _03854_);
  or (_32178_, _32162_, _03855_);
  and (_32179_, _32178_, _03760_);
  and (_32180_, _32179_, _32177_);
  and (_32182_, _31231_, _06108_);
  or (_32183_, _32182_, _32169_);
  and (_32184_, _32183_, _03759_);
  or (_32185_, _32184_, _03752_);
  or (_32186_, _32185_, _32180_);
  and (_32187_, _32171_, _31238_);
  or (_32188_, _32169_, _03753_);
  or (_32189_, _32188_, _32187_);
  and (_32190_, _32189_, _03747_);
  and (_32191_, _32190_, _32186_);
  and (_32193_, _31245_, _06108_);
  or (_32194_, _32193_, _32169_);
  and (_32195_, _32194_, _03746_);
  or (_32196_, _32195_, _07927_);
  or (_32197_, _32196_, _32191_);
  and (_32198_, _06965_, _05500_);
  or (_32199_, _32146_, _03738_);
  or (_32200_, _32199_, _32198_);
  or (_32201_, _32155_, _07925_);
  and (_32202_, _32201_, _03820_);
  and (_32204_, _32202_, _32200_);
  and (_32205_, _32204_, _32197_);
  and (_32206_, _31272_, _05500_);
  or (_32207_, _32206_, _32146_);
  and (_32208_, _32207_, _03455_);
  or (_32209_, _32208_, _03903_);
  or (_32210_, _32209_, _32205_);
  and (_32211_, _32210_, _32153_);
  or (_32212_, _32211_, _03897_);
  and (_32213_, _31283_, _05500_);
  or (_32215_, _32146_, _04790_);
  or (_32216_, _32215_, _32213_);
  and (_32217_, _32216_, _04792_);
  and (_32218_, _32217_, _32212_);
  or (_32219_, _32218_, _32150_);
  and (_32220_, _32219_, _03909_);
  or (_32221_, _32146_, _11240_);
  and (_32222_, _32152_, _03908_);
  and (_32223_, _32222_, _32221_);
  or (_32224_, _32223_, _32220_);
  and (_32226_, _32224_, _04785_);
  and (_32227_, _32162_, _04027_);
  and (_32228_, _32227_, _32221_);
  or (_32229_, _32228_, _03914_);
  or (_32230_, _32229_, _32226_);
  and (_32231_, _31281_, _05500_);
  or (_32232_, _32146_, _06567_);
  or (_32233_, _32232_, _32231_);
  and (_32234_, _32233_, _06572_);
  and (_32235_, _32234_, _32230_);
  and (_32236_, _31180_, _05500_);
  or (_32237_, _32236_, _32146_);
  and (_32238_, _32237_, _04011_);
  or (_32239_, _32238_, _03773_);
  or (_32240_, _32239_, _32235_);
  or (_32241_, _32158_, _03774_);
  and (_32242_, _32241_, _03375_);
  and (_32243_, _32242_, _32240_);
  and (_32244_, _32183_, _03374_);
  or (_32245_, _32244_, _03772_);
  or (_32248_, _32245_, _32243_);
  and (_32249_, _31320_, _05500_);
  or (_32250_, _32146_, _04060_);
  or (_32251_, _32250_, _32249_);
  and (_32252_, _32251_, _43152_);
  and (_32253_, _32252_, _32248_);
  nor (_32254_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_32255_, _32254_, _05397_);
  or (_43537_, _32255_, _32253_);
  and (_32256_, _11257_, \oc8051_golden_model_1.P3 [3]);
  and (_32258_, _31332_, _05500_);
  or (_32259_, _32258_, _32256_);
  and (_32260_, _32259_, _04018_);
  and (_32261_, _05500_, _06345_);
  or (_32262_, _32261_, _32256_);
  or (_32263_, _32262_, _04778_);
  and (_32264_, _31340_, _05500_);
  or (_32265_, _32264_, _32256_);
  or (_32266_, _32265_, _04722_);
  and (_32267_, _05500_, \oc8051_golden_model_1.ACC [3]);
  or (_32269_, _32267_, _32256_);
  and (_32270_, _32269_, _04707_);
  and (_32271_, _04708_, \oc8051_golden_model_1.P3 [3]);
  or (_32272_, _32271_, _03850_);
  or (_32273_, _32272_, _32270_);
  and (_32274_, _32273_, _03764_);
  and (_32275_, _32274_, _32266_);
  and (_32276_, _11265_, \oc8051_golden_model_1.P3 [3]);
  and (_32277_, _31366_, _06108_);
  or (_32278_, _32277_, _32276_);
  and (_32280_, _32278_, _03763_);
  or (_32281_, _32280_, _03848_);
  or (_32282_, _32281_, _32275_);
  and (_32283_, _05500_, _05119_);
  or (_32284_, _32283_, _32256_);
  or (_32285_, _32284_, _04733_);
  and (_32286_, _32285_, _32282_);
  or (_32287_, _32286_, _03854_);
  or (_32288_, _32269_, _03855_);
  and (_32289_, _32288_, _03760_);
  and (_32291_, _32289_, _32287_);
  and (_32292_, _31381_, _06108_);
  or (_32293_, _32292_, _32276_);
  and (_32294_, _32293_, _03759_);
  or (_32295_, _32294_, _03752_);
  or (_32296_, _32295_, _32291_);
  or (_32297_, _32276_, _31388_);
  and (_32298_, _32297_, _32278_);
  or (_32299_, _32298_, _03753_);
  and (_32300_, _32299_, _03747_);
  and (_32302_, _32300_, _32296_);
  and (_32303_, _31394_, _06108_);
  or (_32304_, _32303_, _32276_);
  and (_32305_, _32304_, _03746_);
  or (_32306_, _32305_, _07927_);
  or (_32307_, _32306_, _32302_);
  and (_32308_, _06964_, _05500_);
  or (_32309_, _32256_, _03738_);
  or (_32310_, _32309_, _32308_);
  or (_32311_, _32284_, _07925_);
  and (_32313_, _32311_, _03820_);
  and (_32314_, _32313_, _32310_);
  and (_32315_, _32314_, _32307_);
  and (_32316_, _31421_, _05500_);
  or (_32317_, _32316_, _32256_);
  and (_32318_, _32317_, _03455_);
  or (_32319_, _32318_, _03903_);
  or (_32320_, _32319_, _32315_);
  and (_32321_, _32320_, _32263_);
  or (_32322_, _32321_, _03897_);
  and (_32324_, _31432_, _05500_);
  or (_32325_, _32256_, _04790_);
  or (_32326_, _32325_, _32324_);
  and (_32327_, _32326_, _04792_);
  and (_32328_, _32327_, _32322_);
  or (_32329_, _32328_, _32260_);
  and (_32330_, _32329_, _03909_);
  or (_32331_, _32256_, _11239_);
  and (_32332_, _32262_, _03908_);
  and (_32333_, _32332_, _32331_);
  or (_32335_, _32333_, _32330_);
  and (_32336_, _32335_, _04785_);
  and (_32337_, _32269_, _04027_);
  and (_32338_, _32337_, _32331_);
  or (_32339_, _32338_, _03914_);
  or (_32340_, _32339_, _32336_);
  and (_32341_, _31430_, _05500_);
  or (_32342_, _32256_, _06567_);
  or (_32343_, _32342_, _32341_);
  and (_32344_, _32343_, _06572_);
  and (_32346_, _32344_, _32340_);
  and (_32347_, _31329_, _05500_);
  or (_32348_, _32347_, _32256_);
  and (_32349_, _32348_, _04011_);
  or (_32350_, _32349_, _03773_);
  or (_32351_, _32350_, _32346_);
  or (_32352_, _32265_, _03774_);
  and (_32353_, _32352_, _03375_);
  and (_32354_, _32353_, _32351_);
  and (_32355_, _32293_, _03374_);
  or (_32357_, _32355_, _03772_);
  or (_32358_, _32357_, _32354_);
  and (_32359_, _31469_, _05500_);
  or (_32360_, _32256_, _04060_);
  or (_32361_, _32360_, _32359_);
  and (_32362_, _32361_, _43152_);
  and (_32363_, _32362_, _32358_);
  nor (_32364_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_32365_, _32364_, _05397_);
  or (_43538_, _32365_, _32363_);
  and (_32367_, _11257_, \oc8051_golden_model_1.P3 [4]);
  and (_32368_, _31484_, _05500_);
  or (_32369_, _32368_, _32367_);
  and (_32370_, _32369_, _04018_);
  and (_32371_, _06456_, _05500_);
  or (_32372_, _32371_, _32367_);
  or (_32373_, _32372_, _04778_);
  and (_32374_, _31492_, _05500_);
  or (_32375_, _32374_, _32367_);
  or (_32376_, _32375_, _04722_);
  and (_32378_, _05500_, \oc8051_golden_model_1.ACC [4]);
  or (_32379_, _32378_, _32367_);
  and (_32380_, _32379_, _04707_);
  and (_32381_, _04708_, \oc8051_golden_model_1.P3 [4]);
  or (_32382_, _32381_, _03850_);
  or (_32383_, _32382_, _32380_);
  and (_32384_, _32383_, _03764_);
  and (_32385_, _32384_, _32376_);
  and (_32386_, _11265_, \oc8051_golden_model_1.P3 [4]);
  and (_32387_, _31520_, _06108_);
  or (_32389_, _32387_, _32386_);
  and (_32390_, _32389_, _03763_);
  or (_32391_, _32390_, _03848_);
  or (_32392_, _32391_, _32385_);
  and (_32393_, _05950_, _05500_);
  or (_32394_, _32393_, _32367_);
  or (_32395_, _32394_, _04733_);
  and (_32396_, _32395_, _32392_);
  or (_32397_, _32396_, _03854_);
  or (_32398_, _32379_, _03855_);
  and (_32400_, _32398_, _03760_);
  and (_32401_, _32400_, _32397_);
  and (_32402_, _31535_, _06108_);
  or (_32403_, _32402_, _32386_);
  and (_32404_, _32403_, _03759_);
  or (_32405_, _32404_, _03752_);
  or (_32406_, _32405_, _32401_);
  or (_32407_, _32386_, _31542_);
  and (_32408_, _32407_, _32389_);
  or (_32409_, _32408_, _03753_);
  and (_32411_, _32409_, _03747_);
  and (_32412_, _32411_, _32406_);
  and (_32413_, _31548_, _06108_);
  or (_32414_, _32413_, _32386_);
  and (_32415_, _32414_, _03746_);
  or (_32416_, _32415_, _07927_);
  or (_32417_, _32416_, _32412_);
  and (_32418_, _06969_, _05500_);
  or (_32419_, _32367_, _03738_);
  or (_32420_, _32419_, _32418_);
  or (_32422_, _32394_, _07925_);
  and (_32423_, _32422_, _03820_);
  and (_32424_, _32423_, _32420_);
  and (_32425_, _32424_, _32417_);
  and (_32426_, _31578_, _05500_);
  or (_32427_, _32426_, _32367_);
  and (_32428_, _32427_, _03455_);
  or (_32429_, _32428_, _03903_);
  or (_32430_, _32429_, _32425_);
  and (_32431_, _32430_, _32373_);
  or (_32433_, _32431_, _03897_);
  and (_32434_, _31589_, _05500_);
  or (_32435_, _32434_, _32367_);
  or (_32436_, _32435_, _04790_);
  and (_32437_, _32436_, _04792_);
  and (_32438_, _32437_, _32433_);
  or (_32439_, _32438_, _32370_);
  and (_32440_, _32439_, _03909_);
  or (_32441_, _32367_, _11238_);
  and (_32442_, _32372_, _03908_);
  and (_32444_, _32442_, _32441_);
  or (_32445_, _32444_, _32440_);
  and (_32446_, _32445_, _04785_);
  and (_32447_, _32379_, _04027_);
  and (_32448_, _32447_, _32441_);
  or (_32449_, _32448_, _03914_);
  or (_32450_, _32449_, _32446_);
  and (_32451_, _31587_, _05500_);
  or (_32452_, _32367_, _06567_);
  or (_32453_, _32452_, _32451_);
  and (_32455_, _32453_, _06572_);
  and (_32456_, _32455_, _32450_);
  and (_32457_, _31481_, _05500_);
  or (_32458_, _32457_, _32367_);
  and (_32459_, _32458_, _04011_);
  or (_32460_, _32459_, _03773_);
  or (_32461_, _32460_, _32456_);
  or (_32462_, _32375_, _03774_);
  and (_32463_, _32462_, _03375_);
  and (_32464_, _32463_, _32461_);
  and (_32466_, _32403_, _03374_);
  or (_32467_, _32466_, _03772_);
  or (_32468_, _32467_, _32464_);
  and (_32469_, _31627_, _05500_);
  or (_32470_, _32367_, _04060_);
  or (_32471_, _32470_, _32469_);
  and (_32472_, _32471_, _43152_);
  and (_32473_, _32472_, _32468_);
  nor (_32474_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_32475_, _32474_, _05397_);
  or (_43539_, _32475_, _32473_);
  nor (_32477_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_32478_, _32477_, _05397_);
  and (_32479_, _11257_, \oc8051_golden_model_1.P3 [5]);
  and (_32480_, _31637_, _05500_);
  or (_32481_, _32480_, _32479_);
  and (_32482_, _32481_, _04018_);
  and (_32483_, _06447_, _05500_);
  or (_32484_, _32483_, _32479_);
  or (_32485_, _32484_, _04778_);
  and (_32487_, _31645_, _05500_);
  or (_32488_, _32487_, _32479_);
  or (_32489_, _32488_, _04722_);
  and (_32490_, _05500_, \oc8051_golden_model_1.ACC [5]);
  or (_32491_, _32490_, _32479_);
  and (_32492_, _32491_, _04707_);
  and (_32493_, _04708_, \oc8051_golden_model_1.P3 [5]);
  or (_32494_, _32493_, _03850_);
  or (_32495_, _32494_, _32492_);
  and (_32496_, _32495_, _03764_);
  and (_32498_, _32496_, _32489_);
  and (_32499_, _11265_, \oc8051_golden_model_1.P3 [5]);
  and (_32500_, _31671_, _06108_);
  or (_32501_, _32500_, _32499_);
  and (_32502_, _32501_, _03763_);
  or (_32503_, _32502_, _03848_);
  or (_32504_, _32503_, _32498_);
  and (_32505_, _05857_, _05500_);
  or (_32506_, _32505_, _32479_);
  or (_32507_, _32506_, _04733_);
  and (_32509_, _32507_, _32504_);
  or (_32510_, _32509_, _03854_);
  or (_32511_, _32491_, _03855_);
  and (_32512_, _32511_, _03760_);
  and (_32513_, _32512_, _32510_);
  and (_32514_, _31686_, _06108_);
  or (_32515_, _32514_, _32499_);
  and (_32516_, _32515_, _03759_);
  or (_32517_, _32516_, _03752_);
  or (_32518_, _32517_, _32513_);
  or (_32520_, _32499_, _31693_);
  and (_32521_, _32520_, _32501_);
  or (_32522_, _32521_, _03753_);
  and (_32523_, _32522_, _03747_);
  and (_32524_, _32523_, _32518_);
  and (_32525_, _31699_, _06108_);
  or (_32526_, _32525_, _32499_);
  and (_32527_, _32526_, _03746_);
  or (_32528_, _32527_, _07927_);
  or (_32529_, _32528_, _32524_);
  and (_32531_, _06968_, _05500_);
  or (_32532_, _32479_, _03738_);
  or (_32533_, _32532_, _32531_);
  or (_32534_, _32506_, _07925_);
  and (_32535_, _32534_, _03820_);
  and (_32536_, _32535_, _32533_);
  and (_32537_, _32536_, _32529_);
  and (_32538_, _31727_, _05500_);
  or (_32539_, _32538_, _32479_);
  and (_32540_, _32539_, _03455_);
  or (_32541_, _32540_, _03903_);
  or (_32542_, _32541_, _32537_);
  and (_32543_, _32542_, _32485_);
  or (_32544_, _32543_, _03897_);
  and (_32545_, _31738_, _05500_);
  or (_32546_, _32479_, _04790_);
  or (_32547_, _32546_, _32545_);
  and (_32548_, _32547_, _04792_);
  and (_32549_, _32548_, _32544_);
  or (_32550_, _32549_, _32482_);
  and (_32553_, _32550_, _03909_);
  or (_32554_, _32479_, _11237_);
  and (_32555_, _32484_, _03908_);
  and (_32556_, _32555_, _32554_);
  or (_32557_, _32556_, _32553_);
  and (_32558_, _32557_, _04785_);
  and (_32559_, _32491_, _04027_);
  and (_32560_, _32559_, _32554_);
  or (_32561_, _32560_, _03914_);
  or (_32562_, _32561_, _32558_);
  and (_32564_, _31736_, _05500_);
  or (_32565_, _32479_, _06567_);
  or (_32566_, _32565_, _32564_);
  and (_32567_, _32566_, _06572_);
  and (_32568_, _32567_, _32562_);
  and (_32569_, _31634_, _05500_);
  or (_32570_, _32569_, _32479_);
  and (_32571_, _32570_, _04011_);
  or (_32572_, _32571_, _03773_);
  or (_32573_, _32572_, _32568_);
  or (_32575_, _32488_, _03774_);
  and (_32576_, _32575_, _03375_);
  and (_32577_, _32576_, _32573_);
  and (_32578_, _32515_, _03374_);
  or (_32579_, _32578_, _03772_);
  or (_32580_, _32579_, _32577_);
  and (_32581_, _31775_, _05500_);
  or (_32582_, _32479_, _04060_);
  or (_32583_, _32582_, _32581_);
  and (_32584_, _32583_, _43152_);
  and (_32586_, _32584_, _32580_);
  or (_43542_, _32586_, _32478_);
  nor (_32587_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_32588_, _32587_, _05397_);
  and (_32589_, _11257_, \oc8051_golden_model_1.P3 [6]);
  and (_32590_, _31787_, _05500_);
  or (_32591_, _32590_, _32589_);
  and (_32592_, _32591_, _04018_);
  and (_32593_, _13394_, _05500_);
  or (_32594_, _32593_, _32589_);
  or (_32596_, _32594_, _04778_);
  and (_32597_, _11265_, \oc8051_golden_model_1.P3 [6]);
  and (_32598_, _31807_, _06108_);
  or (_32599_, _32598_, _32597_);
  and (_32600_, _32599_, _03759_);
  and (_32601_, _31813_, _05500_);
  or (_32602_, _32601_, _32589_);
  or (_32603_, _32602_, _04722_);
  and (_32604_, _05500_, \oc8051_golden_model_1.ACC [6]);
  or (_32605_, _32604_, _32589_);
  and (_32607_, _32605_, _04707_);
  and (_32608_, _04708_, \oc8051_golden_model_1.P3 [6]);
  or (_32609_, _32608_, _03850_);
  or (_32610_, _32609_, _32607_);
  and (_32611_, _32610_, _03764_);
  and (_32612_, _32611_, _32603_);
  and (_32613_, _31826_, _06108_);
  or (_32614_, _32613_, _32597_);
  and (_32615_, _32614_, _03763_);
  or (_32616_, _32615_, _03848_);
  or (_32618_, _32616_, _32612_);
  and (_32619_, _06065_, _05500_);
  or (_32620_, _32619_, _32589_);
  or (_32621_, _32620_, _04733_);
  and (_32622_, _32621_, _32618_);
  or (_32623_, _32622_, _03854_);
  or (_32624_, _32605_, _03855_);
  and (_32625_, _32624_, _03760_);
  and (_32626_, _32625_, _32623_);
  or (_32627_, _32626_, _32600_);
  and (_32629_, _32627_, _03753_);
  or (_32630_, _32597_, _31843_);
  and (_32631_, _32630_, _03752_);
  and (_32632_, _32631_, _32614_);
  or (_32633_, _32632_, _32629_);
  and (_32634_, _32633_, _03747_);
  and (_32635_, _31850_, _06108_);
  or (_32636_, _32635_, _32597_);
  and (_32637_, _32636_, _03746_);
  or (_32638_, _32637_, _07927_);
  or (_32640_, _32638_, _32634_);
  and (_32641_, _06641_, _05500_);
  or (_32642_, _32589_, _03738_);
  or (_32643_, _32642_, _32641_);
  or (_32644_, _32620_, _07925_);
  and (_32645_, _32644_, _03820_);
  and (_32646_, _32645_, _32643_);
  and (_32647_, _32646_, _32640_);
  and (_32648_, _31876_, _05500_);
  or (_32649_, _32648_, _32589_);
  and (_32651_, _32649_, _03455_);
  or (_32652_, _32651_, _03903_);
  or (_32653_, _32652_, _32647_);
  and (_32654_, _32653_, _32596_);
  or (_32655_, _32654_, _03897_);
  and (_32656_, _31887_, _05500_);
  or (_32657_, _32589_, _04790_);
  or (_32658_, _32657_, _32656_);
  and (_32659_, _32658_, _04792_);
  and (_32660_, _32659_, _32655_);
  or (_32662_, _32660_, _32592_);
  and (_32663_, _32662_, _03909_);
  or (_32664_, _32589_, _11236_);
  and (_32665_, _32594_, _03908_);
  and (_32666_, _32665_, _32664_);
  or (_32667_, _32666_, _32663_);
  and (_32668_, _32667_, _04785_);
  and (_32669_, _32605_, _04027_);
  and (_32670_, _32669_, _32664_);
  or (_32671_, _32670_, _03914_);
  or (_32673_, _32671_, _32668_);
  and (_32674_, _31885_, _05500_);
  or (_32675_, _32589_, _06567_);
  or (_32676_, _32675_, _32674_);
  and (_32677_, _32676_, _06572_);
  and (_32678_, _32677_, _32673_);
  and (_32679_, _31785_, _05500_);
  or (_32680_, _32679_, _32589_);
  and (_32681_, _32680_, _04011_);
  or (_32682_, _32681_, _03773_);
  or (_32684_, _32682_, _32678_);
  or (_32685_, _32602_, _03774_);
  and (_32686_, _32685_, _03375_);
  and (_32687_, _32686_, _32684_);
  and (_32688_, _32599_, _03374_);
  or (_32689_, _32688_, _03772_);
  or (_32690_, _32689_, _32687_);
  and (_32691_, _31925_, _05500_);
  or (_32692_, _32589_, _04060_);
  or (_32693_, _32692_, _32691_);
  and (_32695_, _32693_, _43152_);
  and (_32696_, _32695_, _32690_);
  or (_43543_, _32696_, _32588_);
  nor (_32697_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_32698_, _32697_, _05397_);
  and (_32699_, _11359_, \oc8051_golden_model_1.P0 [0]);
  and (_32700_, _30893_, _05505_);
  or (_32701_, _32700_, _32699_);
  and (_32702_, _32701_, _04018_);
  and (_32703_, _05505_, _06479_);
  or (_32705_, _32703_, _32699_);
  or (_32706_, _32705_, _04778_);
  and (_32707_, _11126_, _05505_);
  or (_32708_, _32707_, _32699_);
  or (_32709_, _32708_, _04722_);
  and (_32710_, _05505_, \oc8051_golden_model_1.ACC [0]);
  or (_32711_, _32710_, _32699_);
  and (_32712_, _32711_, _04707_);
  and (_32713_, _04708_, \oc8051_golden_model_1.P0 [0]);
  or (_32714_, _32713_, _03850_);
  or (_32716_, _32714_, _32712_);
  and (_32717_, _32716_, _03764_);
  and (_32718_, _32717_, _32709_);
  and (_32719_, _11367_, \oc8051_golden_model_1.P0 [0]);
  and (_32720_, _30926_, _06112_);
  or (_32721_, _32720_, _32719_);
  and (_32722_, _32721_, _03763_);
  or (_32723_, _32722_, _32718_);
  and (_32724_, _32723_, _04733_);
  and (_32725_, _05505_, _04700_);
  or (_32727_, _32725_, _32699_);
  and (_32728_, _32727_, _03848_);
  or (_32729_, _32728_, _03854_);
  or (_32730_, _32729_, _32724_);
  or (_32731_, _32711_, _03855_);
  and (_32732_, _32731_, _03760_);
  and (_32733_, _32732_, _32730_);
  and (_32734_, _32699_, _03759_);
  or (_32735_, _32734_, _03752_);
  or (_32736_, _32735_, _32733_);
  or (_32738_, _32708_, _03753_);
  and (_32739_, _32738_, _03747_);
  and (_32740_, _32739_, _32736_);
  or (_32741_, _32719_, _14237_);
  and (_32742_, _32741_, _03746_);
  and (_32743_, _32742_, _32721_);
  or (_32744_, _32743_, _07927_);
  or (_32745_, _32744_, _32740_);
  and (_32746_, _06962_, _05505_);
  or (_32747_, _32699_, _03738_);
  or (_32749_, _32747_, _32746_);
  or (_32750_, _32727_, _07925_);
  and (_32751_, _32750_, _03820_);
  and (_32752_, _32751_, _32749_);
  and (_32753_, _32752_, _32745_);
  and (_32754_, _30976_, _05505_);
  or (_32755_, _32754_, _32699_);
  and (_32756_, _32755_, _03455_);
  or (_32757_, _32756_, _03903_);
  or (_32758_, _32757_, _32753_);
  and (_32760_, _32758_, _32706_);
  or (_32761_, _32760_, _03897_);
  and (_32762_, _30988_, _05505_);
  or (_32763_, _32699_, _04790_);
  or (_32764_, _32763_, _32762_);
  and (_32765_, _32764_, _04792_);
  and (_32766_, _32765_, _32761_);
  or (_32767_, _32766_, _32702_);
  and (_32768_, _32767_, _03909_);
  nand (_32769_, _32705_, _03908_);
  nor (_32771_, _32769_, _32707_);
  or (_32772_, _32771_, _32768_);
  and (_32773_, _32772_, _04785_);
  or (_32774_, _32699_, _31001_);
  and (_32775_, _32711_, _04027_);
  and (_32776_, _32775_, _32774_);
  or (_32777_, _32776_, _03914_);
  or (_32778_, _32777_, _32773_);
  and (_32779_, _30985_, _05505_);
  or (_32780_, _32699_, _06567_);
  or (_32782_, _32780_, _32779_);
  and (_32783_, _32782_, _06572_);
  and (_32784_, _32783_, _32778_);
  and (_32785_, _30891_, _05505_);
  or (_32786_, _32785_, _32699_);
  and (_32787_, _32786_, _04011_);
  or (_32788_, _32787_, _03773_);
  or (_32789_, _32788_, _32784_);
  or (_32790_, _32708_, _03774_);
  and (_32791_, _32790_, _03375_);
  and (_32793_, _32791_, _32789_);
  and (_32794_, _32699_, _03374_);
  or (_32795_, _32794_, _03772_);
  or (_32796_, _32795_, _32793_);
  or (_32797_, _32708_, _04060_);
  and (_32798_, _32797_, _43152_);
  and (_32799_, _32798_, _32796_);
  or (_43544_, _32799_, _32698_);
  nor (_32800_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_32801_, _32800_, _05397_);
  or (_32803_, _05505_, \oc8051_golden_model_1.P0 [1]);
  and (_32804_, _31037_, _05505_);
  not (_32805_, _32804_);
  and (_32806_, _32805_, _32803_);
  or (_32807_, _32806_, _04722_);
  nand (_32808_, _05505_, _03474_);
  and (_32809_, _32808_, _32803_);
  and (_32810_, _32809_, _04707_);
  and (_32811_, _04708_, \oc8051_golden_model_1.P0 [1]);
  or (_32812_, _32811_, _03850_);
  or (_32814_, _32812_, _32810_);
  and (_32815_, _32814_, _03764_);
  and (_32816_, _32815_, _32807_);
  and (_32817_, _31062_, _06112_);
  and (_32818_, _11367_, \oc8051_golden_model_1.P0 [1]);
  or (_32819_, _32818_, _32817_);
  and (_32820_, _32819_, _03763_);
  or (_32821_, _32820_, _03848_);
  or (_32822_, _32821_, _32816_);
  and (_32823_, _11359_, \oc8051_golden_model_1.P0 [1]);
  and (_32824_, _05505_, _04900_);
  or (_32825_, _32824_, _32823_);
  or (_32826_, _32825_, _04733_);
  and (_32827_, _32826_, _32822_);
  or (_32828_, _32827_, _03854_);
  or (_32829_, _32809_, _03855_);
  and (_32830_, _32829_, _03760_);
  and (_32831_, _32830_, _32828_);
  and (_32832_, _31079_, _06112_);
  or (_32833_, _32832_, _32818_);
  and (_32835_, _32833_, _03759_);
  or (_32836_, _32835_, _32831_);
  and (_32837_, _32836_, _31085_);
  or (_32838_, _32818_, _31087_);
  and (_32839_, _32838_, _03752_);
  and (_32840_, _32839_, _32819_);
  and (_32841_, _31093_, _06112_);
  or (_32842_, _32841_, _32818_);
  and (_32843_, _32842_, _03746_);
  or (_32844_, _32843_, _07927_);
  or (_32846_, _32844_, _32840_);
  or (_32847_, _32846_, _32837_);
  and (_32848_, _06961_, _05505_);
  or (_32849_, _32823_, _03738_);
  or (_32850_, _32849_, _32848_);
  or (_32851_, _32825_, _07925_);
  and (_32852_, _32851_, _03820_);
  and (_32853_, _32852_, _32850_);
  and (_32854_, _32853_, _32847_);
  and (_32855_, _31120_, _05505_);
  or (_32857_, _32855_, _32823_);
  and (_32858_, _32857_, _03455_);
  or (_32859_, _32858_, _32854_);
  and (_32860_, _32859_, _04778_);
  nand (_32861_, _05505_, _04595_);
  and (_32862_, _32803_, _03903_);
  and (_32863_, _32862_, _32861_);
  or (_32864_, _32863_, _32860_);
  and (_32865_, _32864_, _04790_);
  or (_32866_, _31030_, _11359_);
  and (_32868_, _32803_, _03897_);
  and (_32869_, _32868_, _32866_);
  or (_32870_, _32869_, _32865_);
  and (_32871_, _32870_, _04792_);
  or (_32872_, _31137_, _11359_);
  and (_32873_, _32803_, _04018_);
  and (_32874_, _32873_, _32872_);
  or (_32875_, _32874_, _32871_);
  and (_32876_, _32875_, _03909_);
  or (_32877_, _31029_, _11359_);
  and (_32879_, _32803_, _03908_);
  and (_32880_, _32879_, _32877_);
  or (_32881_, _32880_, _32876_);
  and (_32882_, _32881_, _04785_);
  or (_32883_, _32823_, _31149_);
  and (_32884_, _32809_, _04027_);
  and (_32885_, _32884_, _32883_);
  or (_32886_, _32885_, _32882_);
  and (_32887_, _32886_, _04012_);
  or (_32888_, _31134_, _11359_);
  and (_32889_, _32803_, _04011_);
  and (_32890_, _32889_, _32888_);
  or (_32891_, _32890_, _03773_);
  or (_32892_, _32861_, _31149_);
  and (_32893_, _32803_, _03914_);
  and (_32894_, _32893_, _32892_);
  or (_32895_, _32894_, _32891_);
  or (_32896_, _32895_, _32887_);
  or (_32897_, _32806_, _03774_);
  and (_32898_, _32897_, _03375_);
  and (_32901_, _32898_, _32896_);
  and (_32902_, _32833_, _03374_);
  or (_32903_, _32902_, _03772_);
  or (_32904_, _32903_, _32901_);
  or (_32905_, _32823_, _04060_);
  or (_32906_, _32905_, _32804_);
  and (_32907_, _32906_, _43152_);
  and (_32908_, _32907_, _32904_);
  or (_43547_, _32908_, _32801_);
  and (_32909_, _11359_, \oc8051_golden_model_1.P0 [2]);
  and (_32911_, _31182_, _05505_);
  or (_32912_, _32911_, _32909_);
  and (_32913_, _32912_, _04018_);
  and (_32914_, _05505_, _06495_);
  or (_32915_, _32914_, _32909_);
  or (_32916_, _32915_, _04778_);
  and (_32917_, _05505_, _05307_);
  or (_32918_, _32917_, _32909_);
  or (_32919_, _32918_, _04733_);
  and (_32920_, _31194_, _05505_);
  or (_32922_, _32920_, _32909_);
  or (_32923_, _32922_, _04722_);
  and (_32924_, _05505_, \oc8051_golden_model_1.ACC [2]);
  or (_32925_, _32924_, _32909_);
  and (_32926_, _32925_, _04707_);
  and (_32927_, _04708_, \oc8051_golden_model_1.P0 [2]);
  or (_32928_, _32927_, _03850_);
  or (_32929_, _32928_, _32926_);
  and (_32930_, _32929_, _03764_);
  and (_32931_, _32930_, _32923_);
  and (_32933_, _11367_, \oc8051_golden_model_1.P0 [2]);
  and (_32934_, _31219_, _06112_);
  or (_32935_, _32934_, _32933_);
  and (_32936_, _32935_, _03763_);
  or (_32937_, _32936_, _03848_);
  or (_32938_, _32937_, _32931_);
  and (_32939_, _32938_, _32919_);
  or (_32940_, _32939_, _03854_);
  or (_32941_, _32925_, _03855_);
  and (_32942_, _32941_, _03760_);
  and (_32944_, _32942_, _32940_);
  and (_32945_, _31231_, _06112_);
  or (_32946_, _32945_, _32933_);
  and (_32947_, _32946_, _03759_);
  or (_32948_, _32947_, _03752_);
  or (_32949_, _32948_, _32944_);
  and (_32950_, _32934_, _31238_);
  or (_32951_, _32933_, _03753_);
  or (_32952_, _32951_, _32950_);
  and (_32953_, _32952_, _03747_);
  and (_32955_, _32953_, _32949_);
  and (_32956_, _31245_, _06112_);
  or (_32957_, _32956_, _32933_);
  and (_32958_, _32957_, _03746_);
  or (_32959_, _32958_, _07927_);
  or (_32960_, _32959_, _32955_);
  and (_32961_, _06965_, _05505_);
  or (_32962_, _32909_, _03738_);
  or (_32963_, _32962_, _32961_);
  or (_32964_, _32918_, _07925_);
  and (_32966_, _32964_, _03820_);
  and (_32967_, _32966_, _32963_);
  and (_32968_, _32967_, _32960_);
  and (_32969_, _31272_, _05505_);
  or (_32970_, _32969_, _32909_);
  and (_32971_, _32970_, _03455_);
  or (_32972_, _32971_, _03903_);
  or (_32973_, _32972_, _32968_);
  and (_32974_, _32973_, _32916_);
  or (_32975_, _32974_, _03897_);
  and (_32977_, _31283_, _05505_);
  or (_32978_, _32977_, _32909_);
  or (_32979_, _32978_, _04790_);
  and (_32980_, _32979_, _04792_);
  and (_32981_, _32980_, _32975_);
  or (_32982_, _32981_, _32913_);
  and (_32983_, _32982_, _03909_);
  or (_32984_, _32909_, _11240_);
  and (_32985_, _32915_, _03908_);
  and (_32986_, _32985_, _32984_);
  or (_32988_, _32986_, _32983_);
  and (_32989_, _32988_, _04785_);
  and (_32990_, _32925_, _04027_);
  and (_32991_, _32990_, _32984_);
  or (_32992_, _32991_, _03914_);
  or (_32993_, _32992_, _32989_);
  and (_32994_, _31281_, _05505_);
  or (_32995_, _32909_, _06567_);
  or (_32996_, _32995_, _32994_);
  and (_32997_, _32996_, _06572_);
  and (_32999_, _32997_, _32993_);
  and (_33000_, _31180_, _05505_);
  or (_33001_, _33000_, _32909_);
  and (_33002_, _33001_, _04011_);
  or (_33003_, _33002_, _03773_);
  or (_33004_, _33003_, _32999_);
  or (_33005_, _32922_, _03774_);
  and (_33006_, _33005_, _03375_);
  and (_33007_, _33006_, _33004_);
  and (_33008_, _32946_, _03374_);
  or (_33010_, _33008_, _03772_);
  or (_33011_, _33010_, _33007_);
  and (_33012_, _31320_, _05505_);
  or (_33013_, _32909_, _04060_);
  or (_33014_, _33013_, _33012_);
  and (_33015_, _33014_, _43152_);
  and (_33016_, _33015_, _33011_);
  nor (_33017_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_33018_, _33017_, _05397_);
  or (_43548_, _33018_, _33016_);
  and (_33020_, _11359_, \oc8051_golden_model_1.P0 [3]);
  and (_33021_, _31332_, _05505_);
  or (_33022_, _33021_, _33020_);
  and (_33023_, _33022_, _04018_);
  and (_33024_, _05505_, _06345_);
  or (_33025_, _33024_, _33020_);
  or (_33026_, _33025_, _04778_);
  and (_33027_, _31340_, _05505_);
  or (_33028_, _33027_, _33020_);
  or (_33029_, _33028_, _04722_);
  and (_33031_, _05505_, \oc8051_golden_model_1.ACC [3]);
  or (_33032_, _33031_, _33020_);
  and (_33033_, _33032_, _04707_);
  and (_33034_, _04708_, \oc8051_golden_model_1.P0 [3]);
  or (_33035_, _33034_, _03850_);
  or (_33036_, _33035_, _33033_);
  and (_33037_, _33036_, _03764_);
  and (_33038_, _33037_, _33029_);
  and (_33039_, _11367_, \oc8051_golden_model_1.P0 [3]);
  and (_33040_, _31366_, _06112_);
  or (_33042_, _33040_, _33039_);
  and (_33043_, _33042_, _03763_);
  or (_33044_, _33043_, _03848_);
  or (_33045_, _33044_, _33038_);
  and (_33046_, _05505_, _05119_);
  or (_33047_, _33046_, _33020_);
  or (_33048_, _33047_, _04733_);
  and (_33049_, _33048_, _33045_);
  or (_33050_, _33049_, _03854_);
  or (_33051_, _33032_, _03855_);
  and (_33053_, _33051_, _03760_);
  and (_33054_, _33053_, _33050_);
  and (_33055_, _31381_, _06112_);
  or (_33056_, _33055_, _33039_);
  and (_33057_, _33056_, _03759_);
  or (_33058_, _33057_, _03752_);
  or (_33059_, _33058_, _33054_);
  or (_33060_, _33039_, _31388_);
  and (_33061_, _33060_, _33042_);
  or (_33062_, _33061_, _03753_);
  and (_33064_, _33062_, _03747_);
  and (_33065_, _33064_, _33059_);
  and (_33066_, _31394_, _06112_);
  or (_33067_, _33066_, _33039_);
  and (_33068_, _33067_, _03746_);
  or (_33069_, _33068_, _07927_);
  or (_33070_, _33069_, _33065_);
  and (_33071_, _06964_, _05505_);
  or (_33072_, _33020_, _03738_);
  or (_33073_, _33072_, _33071_);
  or (_33075_, _33047_, _07925_);
  and (_33076_, _33075_, _03820_);
  and (_33077_, _33076_, _33073_);
  and (_33078_, _33077_, _33070_);
  and (_33079_, _31421_, _05505_);
  or (_33080_, _33079_, _33020_);
  and (_33081_, _33080_, _03455_);
  or (_33082_, _33081_, _03903_);
  or (_33083_, _33082_, _33078_);
  and (_33084_, _33083_, _33026_);
  or (_33086_, _33084_, _03897_);
  and (_33087_, _31432_, _05505_);
  or (_33088_, _33087_, _33020_);
  or (_33089_, _33088_, _04790_);
  and (_33090_, _33089_, _04792_);
  and (_33091_, _33090_, _33086_);
  or (_33092_, _33091_, _33023_);
  and (_33093_, _33092_, _03909_);
  or (_33094_, _33020_, _11239_);
  and (_33095_, _33025_, _03908_);
  and (_33097_, _33095_, _33094_);
  or (_33098_, _33097_, _33093_);
  and (_33099_, _33098_, _04785_);
  and (_33100_, _33032_, _04027_);
  and (_33101_, _33100_, _33094_);
  or (_33102_, _33101_, _03914_);
  or (_33103_, _33102_, _33099_);
  and (_33104_, _31430_, _05505_);
  or (_33105_, _33020_, _06567_);
  or (_33106_, _33105_, _33104_);
  and (_33108_, _33106_, _06572_);
  and (_33109_, _33108_, _33103_);
  and (_33110_, _31329_, _05505_);
  or (_33111_, _33110_, _33020_);
  and (_33112_, _33111_, _04011_);
  or (_33113_, _33112_, _03773_);
  or (_33114_, _33113_, _33109_);
  or (_33115_, _33028_, _03774_);
  and (_33116_, _33115_, _03375_);
  and (_33117_, _33116_, _33114_);
  and (_33119_, _33056_, _03374_);
  or (_33120_, _33119_, _03772_);
  or (_33121_, _33120_, _33117_);
  and (_33122_, _31469_, _05505_);
  or (_33123_, _33020_, _04060_);
  or (_33124_, _33123_, _33122_);
  and (_33125_, _33124_, _43152_);
  and (_33126_, _33125_, _33121_);
  nor (_33127_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_33128_, _33127_, _05397_);
  or (_43549_, _33128_, _33126_);
  and (_33130_, _11359_, \oc8051_golden_model_1.P0 [4]);
  and (_33131_, _31484_, _05505_);
  or (_33132_, _33131_, _33130_);
  and (_33133_, _33132_, _04018_);
  and (_33134_, _06456_, _05505_);
  or (_33135_, _33134_, _33130_);
  or (_33136_, _33135_, _04778_);
  and (_33137_, _31492_, _05505_);
  or (_33138_, _33137_, _33130_);
  or (_33140_, _33138_, _04722_);
  and (_33141_, _05505_, \oc8051_golden_model_1.ACC [4]);
  or (_33142_, _33141_, _33130_);
  and (_33143_, _33142_, _04707_);
  and (_33144_, _04708_, \oc8051_golden_model_1.P0 [4]);
  or (_33145_, _33144_, _03850_);
  or (_33146_, _33145_, _33143_);
  and (_33147_, _33146_, _03764_);
  and (_33148_, _33147_, _33140_);
  and (_33149_, _11367_, \oc8051_golden_model_1.P0 [4]);
  and (_33151_, _31520_, _06112_);
  or (_33152_, _33151_, _33149_);
  and (_33153_, _33152_, _03763_);
  or (_33154_, _33153_, _03848_);
  or (_33155_, _33154_, _33148_);
  and (_33156_, _05950_, _05505_);
  or (_33157_, _33156_, _33130_);
  or (_33158_, _33157_, _04733_);
  and (_33159_, _33158_, _33155_);
  or (_33160_, _33159_, _03854_);
  or (_33162_, _33142_, _03855_);
  and (_33163_, _33162_, _03760_);
  and (_33164_, _33163_, _33160_);
  and (_33165_, _31535_, _06112_);
  or (_33166_, _33165_, _33149_);
  and (_33167_, _33166_, _03759_);
  or (_33168_, _33167_, _03752_);
  or (_33169_, _33168_, _33164_);
  or (_33170_, _33149_, _31542_);
  and (_33171_, _33170_, _33152_);
  or (_33173_, _33171_, _03753_);
  and (_33174_, _33173_, _03747_);
  and (_33175_, _33174_, _33169_);
  and (_33176_, _31548_, _06112_);
  or (_33177_, _33176_, _33149_);
  and (_33178_, _33177_, _03746_);
  or (_33179_, _33178_, _07927_);
  or (_33180_, _33179_, _33175_);
  and (_33181_, _06969_, _05505_);
  or (_33182_, _33130_, _03738_);
  or (_33184_, _33182_, _33181_);
  or (_33185_, _33157_, _07925_);
  and (_33186_, _33185_, _03820_);
  and (_33187_, _33186_, _33184_);
  and (_33188_, _33187_, _33180_);
  and (_33189_, _31578_, _05505_);
  or (_33190_, _33189_, _33130_);
  and (_33191_, _33190_, _03455_);
  or (_33192_, _33191_, _03903_);
  or (_33193_, _33192_, _33188_);
  and (_33195_, _33193_, _33136_);
  or (_33196_, _33195_, _03897_);
  and (_33197_, _31589_, _05505_);
  or (_33198_, _33130_, _04790_);
  or (_33199_, _33198_, _33197_);
  and (_33200_, _33199_, _04792_);
  and (_33201_, _33200_, _33196_);
  or (_33202_, _33201_, _33133_);
  and (_33203_, _33202_, _03909_);
  or (_33204_, _33130_, _11238_);
  and (_33206_, _33135_, _03908_);
  and (_33207_, _33206_, _33204_);
  or (_33208_, _33207_, _33203_);
  and (_33209_, _33208_, _04785_);
  and (_33210_, _33142_, _04027_);
  and (_33211_, _33210_, _33204_);
  or (_33212_, _33211_, _03914_);
  or (_33213_, _33212_, _33209_);
  and (_33214_, _31587_, _05505_);
  or (_33215_, _33130_, _06567_);
  or (_33217_, _33215_, _33214_);
  and (_33218_, _33217_, _06572_);
  and (_33219_, _33218_, _33213_);
  and (_33220_, _31481_, _05505_);
  or (_33221_, _33220_, _33130_);
  and (_33222_, _33221_, _04011_);
  or (_33223_, _33222_, _03773_);
  or (_33224_, _33223_, _33219_);
  or (_33225_, _33138_, _03774_);
  and (_33226_, _33225_, _03375_);
  and (_33228_, _33226_, _33224_);
  and (_33229_, _33166_, _03374_);
  or (_33230_, _33229_, _03772_);
  or (_33231_, _33230_, _33228_);
  and (_33232_, _31627_, _05505_);
  or (_33233_, _33130_, _04060_);
  or (_33234_, _33233_, _33232_);
  and (_33235_, _33234_, _43152_);
  and (_33236_, _33235_, _33231_);
  nor (_33237_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_33239_, _33237_, _05397_);
  or (_43550_, _33239_, _33236_);
  and (_33240_, _11359_, \oc8051_golden_model_1.P0 [5]);
  and (_33241_, _31637_, _05505_);
  or (_33242_, _33241_, _33240_);
  and (_33243_, _33242_, _04018_);
  and (_33244_, _06447_, _05505_);
  or (_33245_, _33244_, _33240_);
  or (_33246_, _33245_, _04778_);
  and (_33247_, _31645_, _05505_);
  or (_33249_, _33247_, _33240_);
  or (_33250_, _33249_, _04722_);
  and (_33251_, _05505_, \oc8051_golden_model_1.ACC [5]);
  or (_33252_, _33251_, _33240_);
  and (_33253_, _33252_, _04707_);
  and (_33254_, _04708_, \oc8051_golden_model_1.P0 [5]);
  or (_33255_, _33254_, _03850_);
  or (_33256_, _33255_, _33253_);
  and (_33257_, _33256_, _03764_);
  and (_33258_, _33257_, _33250_);
  and (_33259_, _11367_, \oc8051_golden_model_1.P0 [5]);
  and (_33260_, _31671_, _06112_);
  or (_33261_, _33260_, _33259_);
  and (_33262_, _33261_, _03763_);
  or (_33263_, _33262_, _03848_);
  or (_33264_, _33263_, _33258_);
  and (_33265_, _05857_, _05505_);
  or (_33266_, _33265_, _33240_);
  or (_33267_, _33266_, _04733_);
  and (_33268_, _33267_, _33264_);
  or (_33271_, _33268_, _03854_);
  or (_33272_, _33252_, _03855_);
  and (_33273_, _33272_, _03760_);
  and (_33274_, _33273_, _33271_);
  and (_33275_, _31686_, _06112_);
  or (_33276_, _33275_, _33259_);
  and (_33277_, _33276_, _03759_);
  or (_33278_, _33277_, _03752_);
  or (_33279_, _33278_, _33274_);
  or (_33280_, _33259_, _31693_);
  and (_33282_, _33280_, _33261_);
  or (_33283_, _33282_, _03753_);
  and (_33284_, _33283_, _03747_);
  and (_33285_, _33284_, _33279_);
  and (_33286_, _31699_, _06112_);
  or (_33287_, _33286_, _33259_);
  and (_33288_, _33287_, _03746_);
  or (_33289_, _33288_, _07927_);
  or (_33290_, _33289_, _33285_);
  and (_33291_, _06968_, _05505_);
  or (_33293_, _33240_, _03738_);
  or (_33294_, _33293_, _33291_);
  or (_33295_, _33266_, _07925_);
  and (_33296_, _33295_, _03820_);
  and (_33297_, _33296_, _33294_);
  and (_33298_, _33297_, _33290_);
  and (_33299_, _31727_, _05505_);
  or (_33300_, _33299_, _33240_);
  and (_33301_, _33300_, _03455_);
  or (_33302_, _33301_, _03903_);
  or (_33304_, _33302_, _33298_);
  and (_33305_, _33304_, _33246_);
  or (_33306_, _33305_, _03897_);
  and (_33307_, _31738_, _05505_);
  or (_33308_, _33307_, _33240_);
  or (_33309_, _33308_, _04790_);
  and (_33310_, _33309_, _04792_);
  and (_33311_, _33310_, _33306_);
  or (_33312_, _33311_, _33243_);
  and (_33313_, _33312_, _03909_);
  or (_33315_, _33240_, _11237_);
  and (_33316_, _33245_, _03908_);
  and (_33317_, _33316_, _33315_);
  or (_33318_, _33317_, _33313_);
  and (_33319_, _33318_, _04785_);
  and (_33320_, _33252_, _04027_);
  and (_33321_, _33320_, _33315_);
  or (_33322_, _33321_, _03914_);
  or (_33323_, _33322_, _33319_);
  and (_33324_, _31736_, _05505_);
  or (_33326_, _33240_, _06567_);
  or (_33327_, _33326_, _33324_);
  and (_33328_, _33327_, _06572_);
  and (_33329_, _33328_, _33323_);
  and (_33330_, _31634_, _05505_);
  or (_33331_, _33330_, _33240_);
  and (_33332_, _33331_, _04011_);
  or (_33333_, _33332_, _03773_);
  or (_33334_, _33333_, _33329_);
  or (_33335_, _33249_, _03774_);
  and (_33337_, _33335_, _03375_);
  and (_33338_, _33337_, _33334_);
  and (_33339_, _33276_, _03374_);
  or (_33340_, _33339_, _03772_);
  or (_33341_, _33340_, _33338_);
  and (_33342_, _31775_, _05505_);
  or (_33343_, _33240_, _04060_);
  or (_33344_, _33343_, _33342_);
  and (_33345_, _33344_, _43152_);
  and (_33346_, _33345_, _33341_);
  nor (_33348_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_33349_, _33348_, _05397_);
  or (_43551_, _33349_, _33346_);
  nor (_33350_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_33351_, _33350_, _05397_);
  and (_33352_, _11359_, \oc8051_golden_model_1.P0 [6]);
  and (_33353_, _31787_, _05505_);
  or (_33354_, _33353_, _33352_);
  and (_33355_, _33354_, _04018_);
  and (_33356_, _13394_, _05505_);
  or (_33358_, _33356_, _33352_);
  or (_33359_, _33358_, _04778_);
  and (_33360_, _11367_, \oc8051_golden_model_1.P0 [6]);
  and (_33361_, _31807_, _06112_);
  or (_33362_, _33361_, _33360_);
  and (_33363_, _33362_, _03759_);
  and (_33364_, _31813_, _05505_);
  or (_33365_, _33364_, _33352_);
  or (_33366_, _33365_, _04722_);
  and (_33367_, _05505_, \oc8051_golden_model_1.ACC [6]);
  or (_33369_, _33367_, _33352_);
  and (_33370_, _33369_, _04707_);
  and (_33371_, _04708_, \oc8051_golden_model_1.P0 [6]);
  or (_33372_, _33371_, _03850_);
  or (_33373_, _33372_, _33370_);
  and (_33374_, _33373_, _03764_);
  and (_33375_, _33374_, _33366_);
  and (_33376_, _31826_, _06112_);
  or (_33377_, _33376_, _33360_);
  and (_33378_, _33377_, _03763_);
  or (_33380_, _33378_, _03848_);
  or (_33381_, _33380_, _33375_);
  and (_33382_, _06065_, _05505_);
  or (_33383_, _33382_, _33352_);
  or (_33384_, _33383_, _04733_);
  and (_33385_, _33384_, _33381_);
  or (_33386_, _33385_, _03854_);
  or (_33387_, _33369_, _03855_);
  and (_33388_, _33387_, _03760_);
  and (_33389_, _33388_, _33386_);
  or (_33391_, _33389_, _33363_);
  and (_33392_, _33391_, _03753_);
  or (_33393_, _33360_, _31843_);
  and (_33394_, _33393_, _03752_);
  and (_33395_, _33394_, _33377_);
  or (_33396_, _33395_, _33392_);
  and (_33397_, _33396_, _03747_);
  and (_33398_, _31850_, _06112_);
  or (_33399_, _33398_, _33360_);
  and (_33400_, _33399_, _03746_);
  or (_33402_, _33400_, _07927_);
  or (_33403_, _33402_, _33397_);
  and (_33404_, _06641_, _05505_);
  or (_33405_, _33352_, _03738_);
  or (_33406_, _33405_, _33404_);
  or (_33407_, _33383_, _07925_);
  and (_33408_, _33407_, _03820_);
  and (_33409_, _33408_, _33406_);
  and (_33410_, _33409_, _33403_);
  and (_33411_, _31876_, _05505_);
  or (_33413_, _33411_, _33352_);
  and (_33414_, _33413_, _03455_);
  or (_33415_, _33414_, _03903_);
  or (_33416_, _33415_, _33410_);
  and (_33417_, _33416_, _33359_);
  or (_33418_, _33417_, _03897_);
  and (_33419_, _31887_, _05505_);
  or (_33420_, _33352_, _04790_);
  or (_33421_, _33420_, _33419_);
  and (_33422_, _33421_, _04792_);
  and (_33424_, _33422_, _33418_);
  or (_33425_, _33424_, _33355_);
  and (_33426_, _33425_, _03909_);
  or (_33427_, _33352_, _11236_);
  and (_33428_, _33358_, _03908_);
  and (_33429_, _33428_, _33427_);
  or (_33430_, _33429_, _33426_);
  and (_33431_, _33430_, _04785_);
  and (_33432_, _33369_, _04027_);
  and (_33433_, _33432_, _33427_);
  or (_33435_, _33433_, _03914_);
  or (_33436_, _33435_, _33431_);
  and (_33437_, _31885_, _05505_);
  or (_33438_, _33352_, _06567_);
  or (_33439_, _33438_, _33437_);
  and (_33440_, _33439_, _06572_);
  and (_33441_, _33440_, _33436_);
  and (_33442_, _31785_, _05505_);
  or (_33443_, _33442_, _33352_);
  and (_33444_, _33443_, _04011_);
  or (_33446_, _33444_, _03773_);
  or (_33447_, _33446_, _33441_);
  or (_33448_, _33365_, _03774_);
  and (_33449_, _33448_, _03375_);
  and (_33450_, _33449_, _33447_);
  and (_33451_, _33362_, _03374_);
  or (_33452_, _33451_, _03772_);
  or (_33453_, _33452_, _33450_);
  and (_33454_, _31925_, _05505_);
  or (_33455_, _33352_, _04060_);
  or (_33457_, _33455_, _33454_);
  and (_33458_, _33457_, _43152_);
  and (_33459_, _33458_, _33453_);
  or (_43552_, _33459_, _33351_);
  and (_33460_, _11461_, \oc8051_golden_model_1.P1 [0]);
  and (_33461_, _30893_, _05455_);
  or (_33462_, _33461_, _33460_);
  and (_33463_, _33462_, _04018_);
  and (_33464_, _05455_, _06479_);
  or (_33465_, _33464_, _33460_);
  or (_33467_, _33465_, _04778_);
  and (_33468_, _11469_, \oc8051_golden_model_1.P1 [0]);
  and (_33469_, _30926_, _06114_);
  or (_33470_, _33469_, _33468_);
  or (_33471_, _33470_, _03764_);
  and (_33472_, _11126_, _05455_);
  or (_33473_, _33472_, _33460_);
  and (_33474_, _33473_, _03850_);
  and (_33475_, _04708_, \oc8051_golden_model_1.P1 [0]);
  and (_33476_, _05455_, \oc8051_golden_model_1.ACC [0]);
  or (_33478_, _33476_, _33460_);
  and (_33479_, _33478_, _04707_);
  or (_33480_, _33479_, _33475_);
  and (_33481_, _33480_, _04722_);
  or (_33482_, _33481_, _03763_);
  or (_33483_, _33482_, _33474_);
  and (_33484_, _33483_, _33471_);
  and (_33485_, _33484_, _04733_);
  and (_33486_, _05455_, _04700_);
  or (_33487_, _33486_, _33460_);
  and (_33489_, _33487_, _03848_);
  or (_33490_, _33489_, _03854_);
  or (_33491_, _33490_, _33485_);
  or (_33492_, _33478_, _03855_);
  and (_33493_, _33492_, _03760_);
  and (_33494_, _33493_, _33491_);
  and (_33495_, _33460_, _03759_);
  or (_33496_, _33495_, _03752_);
  or (_33497_, _33496_, _33494_);
  or (_33498_, _33473_, _03753_);
  and (_33500_, _33498_, _03747_);
  and (_33501_, _33500_, _33497_);
  or (_33502_, _33468_, _14237_);
  and (_33503_, _33502_, _03746_);
  and (_33504_, _33503_, _33470_);
  or (_33505_, _33504_, _07927_);
  or (_33506_, _33505_, _33501_);
  and (_33507_, _06962_, _05455_);
  or (_33508_, _33460_, _03738_);
  or (_33509_, _33508_, _33507_);
  or (_33511_, _33487_, _07925_);
  and (_33512_, _33511_, _03820_);
  and (_33513_, _33512_, _33509_);
  and (_33514_, _33513_, _33506_);
  and (_33515_, _30976_, _05455_);
  or (_33516_, _33515_, _33460_);
  and (_33517_, _33516_, _03455_);
  or (_33518_, _33517_, _03903_);
  or (_33519_, _33518_, _33514_);
  and (_33520_, _33519_, _33467_);
  or (_33522_, _33520_, _03897_);
  and (_33523_, _30988_, _05455_);
  or (_33524_, _33523_, _33460_);
  or (_33525_, _33524_, _04790_);
  and (_33526_, _33525_, _04792_);
  and (_33527_, _33526_, _33522_);
  or (_33528_, _33527_, _33463_);
  and (_33529_, _33528_, _03909_);
  nand (_33530_, _33465_, _03908_);
  nor (_33531_, _33530_, _33472_);
  or (_33533_, _33531_, _33529_);
  and (_33534_, _33533_, _04785_);
  or (_33535_, _33460_, _31001_);
  and (_33536_, _33478_, _04027_);
  and (_33537_, _33536_, _33535_);
  or (_33538_, _33537_, _03914_);
  or (_33539_, _33538_, _33534_);
  and (_33540_, _30985_, _05455_);
  or (_33541_, _33460_, _06567_);
  or (_33542_, _33541_, _33540_);
  and (_33544_, _33542_, _06572_);
  and (_33545_, _33544_, _33539_);
  and (_33546_, _30891_, _05455_);
  or (_33547_, _33546_, _33460_);
  and (_33548_, _33547_, _04011_);
  or (_33549_, _33548_, _03773_);
  or (_33550_, _33549_, _33545_);
  or (_33551_, _33473_, _03774_);
  and (_33552_, _33551_, _03375_);
  and (_33553_, _33552_, _33550_);
  and (_33554_, _33460_, _03374_);
  or (_33555_, _33554_, _03772_);
  or (_33556_, _33555_, _33553_);
  or (_33557_, _33473_, _04060_);
  and (_33558_, _33557_, _43152_);
  and (_33559_, _33558_, _33556_);
  nor (_33560_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_33561_, _33560_, _05397_);
  or (_43553_, _33561_, _33559_);
  or (_33562_, _31030_, _11461_);
  or (_33564_, _05455_, \oc8051_golden_model_1.P1 [1]);
  and (_33565_, _33564_, _03897_);
  and (_33566_, _33565_, _33562_);
  nand (_33567_, _05455_, _04595_);
  and (_33568_, _33564_, _03903_);
  and (_33569_, _33568_, _33567_);
  and (_33570_, _11469_, \oc8051_golden_model_1.P1 [1]);
  and (_33571_, _31079_, _06114_);
  or (_33572_, _33571_, _33570_);
  and (_33573_, _33572_, _03759_);
  and (_33575_, _31037_, _05455_);
  not (_33576_, _33575_);
  and (_33577_, _33576_, _33564_);
  or (_33578_, _33577_, _04722_);
  nand (_33579_, _05455_, _03474_);
  and (_33580_, _33579_, _33564_);
  and (_33581_, _33580_, _04707_);
  and (_33582_, _04708_, \oc8051_golden_model_1.P1 [1]);
  or (_33583_, _33582_, _03850_);
  or (_33584_, _33583_, _33581_);
  and (_33586_, _33584_, _03764_);
  and (_33587_, _33586_, _33578_);
  and (_33588_, _31062_, _06114_);
  or (_33589_, _33588_, _33570_);
  and (_33590_, _33589_, _03763_);
  or (_33591_, _33590_, _03848_);
  or (_33592_, _33591_, _33587_);
  and (_33593_, _11461_, \oc8051_golden_model_1.P1 [1]);
  and (_33594_, _05455_, _04900_);
  or (_33595_, _33594_, _33593_);
  or (_33597_, _33595_, _04733_);
  and (_33598_, _33597_, _33592_);
  or (_33599_, _33598_, _03854_);
  or (_33600_, _33580_, _03855_);
  and (_33601_, _33600_, _03760_);
  and (_33602_, _33601_, _33599_);
  or (_33603_, _33602_, _33573_);
  and (_33604_, _33603_, _31085_);
  or (_33605_, _33570_, _31087_);
  and (_33606_, _33605_, _03752_);
  and (_33608_, _33606_, _33589_);
  and (_33609_, _31093_, _06114_);
  or (_33610_, _33609_, _33570_);
  and (_33611_, _33610_, _03746_);
  or (_33612_, _33611_, _07927_);
  or (_33613_, _33612_, _33608_);
  or (_33614_, _33613_, _33604_);
  and (_33615_, _06961_, _05455_);
  or (_33616_, _33593_, _03738_);
  or (_33617_, _33616_, _33615_);
  or (_33619_, _33595_, _07925_);
  and (_33620_, _33619_, _03820_);
  and (_33621_, _33620_, _33617_);
  and (_33622_, _33621_, _33614_);
  and (_33623_, _31120_, _05455_);
  or (_33624_, _33623_, _33593_);
  and (_33625_, _33624_, _03455_);
  or (_33626_, _33625_, _33622_);
  and (_33627_, _33626_, _04778_);
  or (_33628_, _33627_, _33569_);
  and (_33630_, _33628_, _04790_);
  or (_33631_, _33630_, _33566_);
  and (_33632_, _33631_, _04792_);
  or (_33633_, _31137_, _11461_);
  and (_33634_, _33564_, _04018_);
  and (_33635_, _33634_, _33633_);
  or (_33636_, _33635_, _33632_);
  and (_33637_, _33636_, _03909_);
  or (_33638_, _31029_, _11461_);
  and (_33639_, _33564_, _03908_);
  and (_33641_, _33639_, _33638_);
  or (_33642_, _33641_, _33637_);
  and (_33643_, _33642_, _04785_);
  or (_33644_, _33593_, _31149_);
  and (_33645_, _33580_, _04027_);
  and (_33646_, _33645_, _33644_);
  or (_33647_, _33646_, _33643_);
  and (_33648_, _33647_, _04012_);
  or (_33649_, _33567_, _31149_);
  and (_33650_, _33564_, _03914_);
  and (_33652_, _33650_, _33649_);
  or (_33653_, _33579_, _31149_);
  and (_33654_, _33564_, _04011_);
  and (_33655_, _33654_, _33653_);
  or (_33656_, _33655_, _03773_);
  or (_33657_, _33656_, _33652_);
  or (_33658_, _33657_, _33648_);
  or (_33659_, _33577_, _03774_);
  and (_33660_, _33659_, _03375_);
  and (_33661_, _33660_, _33658_);
  and (_33663_, _33572_, _03374_);
  or (_33664_, _33663_, _03772_);
  or (_33665_, _33664_, _33661_);
  or (_33666_, _33593_, _04060_);
  or (_33667_, _33666_, _33575_);
  and (_33668_, _33667_, _43152_);
  and (_33669_, _33668_, _33665_);
  nor (_33670_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_33671_, _33670_, _05397_);
  or (_43554_, _33671_, _33669_);
  and (_33673_, _11461_, \oc8051_golden_model_1.P1 [2]);
  and (_33674_, _31182_, _05455_);
  or (_33675_, _33674_, _33673_);
  and (_33676_, _33675_, _04018_);
  and (_33677_, _05455_, _06495_);
  or (_33678_, _33677_, _33673_);
  or (_33679_, _33678_, _04778_);
  and (_33680_, _05455_, _05307_);
  or (_33681_, _33680_, _33673_);
  or (_33682_, _33681_, _04733_);
  and (_33684_, _31194_, _05455_);
  or (_33685_, _33684_, _33673_);
  or (_33686_, _33685_, _04722_);
  and (_33687_, _05455_, \oc8051_golden_model_1.ACC [2]);
  or (_33688_, _33687_, _33673_);
  and (_33689_, _33688_, _04707_);
  and (_33690_, _04708_, \oc8051_golden_model_1.P1 [2]);
  or (_33691_, _33690_, _03850_);
  or (_33692_, _33691_, _33689_);
  and (_33693_, _33692_, _03764_);
  and (_33695_, _33693_, _33686_);
  and (_33696_, _11469_, \oc8051_golden_model_1.P1 [2]);
  and (_33697_, _31219_, _06114_);
  or (_33698_, _33697_, _33696_);
  and (_33699_, _33698_, _03763_);
  or (_33700_, _33699_, _03848_);
  or (_33701_, _33700_, _33695_);
  and (_33702_, _33701_, _33682_);
  or (_33703_, _33702_, _03854_);
  or (_33704_, _33688_, _03855_);
  and (_33706_, _33704_, _03760_);
  and (_33707_, _33706_, _33703_);
  and (_33708_, _31231_, _06114_);
  or (_33709_, _33708_, _33696_);
  and (_33710_, _33709_, _03759_);
  or (_33711_, _33710_, _03752_);
  or (_33712_, _33711_, _33707_);
  and (_33713_, _33697_, _31238_);
  or (_33714_, _33696_, _03753_);
  or (_33715_, _33714_, _33713_);
  and (_33717_, _33715_, _03747_);
  and (_33718_, _33717_, _33712_);
  and (_33719_, _31245_, _06114_);
  or (_33720_, _33719_, _33696_);
  and (_33721_, _33720_, _03746_);
  or (_33722_, _33721_, _07927_);
  or (_33723_, _33722_, _33718_);
  and (_33724_, _06965_, _05455_);
  or (_33725_, _33673_, _03738_);
  or (_33726_, _33725_, _33724_);
  or (_33728_, _33681_, _07925_);
  and (_33729_, _33728_, _03820_);
  and (_33730_, _33729_, _33726_);
  and (_33731_, _33730_, _33723_);
  and (_33732_, _31272_, _05455_);
  or (_33733_, _33732_, _33673_);
  and (_33734_, _33733_, _03455_);
  or (_33735_, _33734_, _03903_);
  or (_33736_, _33735_, _33731_);
  and (_33737_, _33736_, _33679_);
  or (_33739_, _33737_, _03897_);
  and (_33740_, _31283_, _05455_);
  or (_33741_, _33673_, _04790_);
  or (_33742_, _33741_, _33740_);
  and (_33743_, _33742_, _04792_);
  and (_33744_, _33743_, _33739_);
  or (_33745_, _33744_, _33676_);
  and (_33746_, _33745_, _03909_);
  or (_33747_, _33673_, _11240_);
  and (_33748_, _33678_, _03908_);
  and (_33750_, _33748_, _33747_);
  or (_33751_, _33750_, _33746_);
  and (_33752_, _33751_, _04785_);
  and (_33753_, _33688_, _04027_);
  and (_33754_, _33753_, _33747_);
  or (_33755_, _33754_, _03914_);
  or (_33756_, _33755_, _33752_);
  and (_33757_, _31281_, _05455_);
  or (_33758_, _33673_, _06567_);
  or (_33759_, _33758_, _33757_);
  and (_33761_, _33759_, _06572_);
  and (_33762_, _33761_, _33756_);
  and (_33763_, _31180_, _05455_);
  or (_33764_, _33763_, _33673_);
  and (_33765_, _33764_, _04011_);
  or (_33766_, _33765_, _03773_);
  or (_33767_, _33766_, _33762_);
  or (_33768_, _33685_, _03774_);
  and (_33769_, _33768_, _03375_);
  and (_33770_, _33769_, _33767_);
  and (_33772_, _33709_, _03374_);
  or (_33773_, _33772_, _03772_);
  or (_33774_, _33773_, _33770_);
  and (_33775_, _31320_, _05455_);
  or (_33776_, _33673_, _04060_);
  or (_33777_, _33776_, _33775_);
  and (_33778_, _33777_, _43152_);
  and (_33779_, _33778_, _33774_);
  nor (_33780_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_33781_, _33780_, _05397_);
  or (_43555_, _33781_, _33779_);
  and (_33782_, _11461_, \oc8051_golden_model_1.P1 [3]);
  and (_33783_, _31332_, _05455_);
  or (_33784_, _33783_, _33782_);
  and (_33785_, _33784_, _04018_);
  and (_33786_, _05455_, _06345_);
  or (_33787_, _33786_, _33782_);
  or (_33788_, _33787_, _04778_);
  and (_33789_, _31340_, _05455_);
  or (_33790_, _33789_, _33782_);
  or (_33793_, _33790_, _04722_);
  and (_33794_, _05455_, \oc8051_golden_model_1.ACC [3]);
  or (_33795_, _33794_, _33782_);
  and (_33796_, _33795_, _04707_);
  and (_33797_, _04708_, \oc8051_golden_model_1.P1 [3]);
  or (_33798_, _33797_, _03850_);
  or (_33799_, _33798_, _33796_);
  and (_33800_, _33799_, _03764_);
  and (_33801_, _33800_, _33793_);
  and (_33802_, _11469_, \oc8051_golden_model_1.P1 [3]);
  and (_33804_, _31366_, _06114_);
  or (_33805_, _33804_, _33802_);
  and (_33806_, _33805_, _03763_);
  or (_33807_, _33806_, _03848_);
  or (_33808_, _33807_, _33801_);
  and (_33809_, _05455_, _05119_);
  or (_33810_, _33809_, _33782_);
  or (_33811_, _33810_, _04733_);
  and (_33812_, _33811_, _33808_);
  or (_33813_, _33812_, _03854_);
  or (_33815_, _33795_, _03855_);
  and (_33816_, _33815_, _03760_);
  and (_33817_, _33816_, _33813_);
  and (_33818_, _31381_, _06114_);
  or (_33819_, _33818_, _33802_);
  and (_33820_, _33819_, _03759_);
  or (_33821_, _33820_, _03752_);
  or (_33822_, _33821_, _33817_);
  or (_33823_, _33802_, _31388_);
  and (_33824_, _33823_, _33805_);
  or (_33826_, _33824_, _03753_);
  and (_33827_, _33826_, _03747_);
  and (_33828_, _33827_, _33822_);
  and (_33829_, _31394_, _06114_);
  or (_33830_, _33829_, _33802_);
  and (_33831_, _33830_, _03746_);
  or (_33832_, _33831_, _07927_);
  or (_33833_, _33832_, _33828_);
  and (_33834_, _06964_, _05455_);
  or (_33835_, _33782_, _03738_);
  or (_33837_, _33835_, _33834_);
  or (_33838_, _33810_, _07925_);
  and (_33839_, _33838_, _03820_);
  and (_33840_, _33839_, _33837_);
  and (_33841_, _33840_, _33833_);
  and (_33842_, _31421_, _05455_);
  or (_33843_, _33842_, _33782_);
  and (_33844_, _33843_, _03455_);
  or (_33845_, _33844_, _03903_);
  or (_33846_, _33845_, _33841_);
  and (_33848_, _33846_, _33788_);
  or (_33849_, _33848_, _03897_);
  and (_33850_, _31432_, _05455_);
  or (_33851_, _33850_, _33782_);
  or (_33852_, _33851_, _04790_);
  and (_33853_, _33852_, _04792_);
  and (_33854_, _33853_, _33849_);
  or (_33855_, _33854_, _33785_);
  and (_33856_, _33855_, _03909_);
  or (_33857_, _33782_, _11239_);
  and (_33859_, _33787_, _03908_);
  and (_33860_, _33859_, _33857_);
  or (_33861_, _33860_, _33856_);
  and (_33862_, _33861_, _04785_);
  and (_33863_, _33795_, _04027_);
  and (_33864_, _33863_, _33857_);
  or (_33865_, _33864_, _03914_);
  or (_33866_, _33865_, _33862_);
  and (_33867_, _31430_, _05455_);
  or (_33868_, _33782_, _06567_);
  or (_33870_, _33868_, _33867_);
  and (_33871_, _33870_, _06572_);
  and (_33872_, _33871_, _33866_);
  and (_33873_, _31329_, _05455_);
  or (_33874_, _33873_, _33782_);
  and (_33875_, _33874_, _04011_);
  or (_33876_, _33875_, _03773_);
  or (_33877_, _33876_, _33872_);
  or (_33878_, _33790_, _03774_);
  and (_33879_, _33878_, _03375_);
  and (_33881_, _33879_, _33877_);
  and (_33882_, _33819_, _03374_);
  or (_33883_, _33882_, _03772_);
  or (_33884_, _33883_, _33881_);
  and (_33885_, _31469_, _05455_);
  or (_33886_, _33782_, _04060_);
  or (_33887_, _33886_, _33885_);
  and (_33888_, _33887_, _43152_);
  and (_33889_, _33888_, _33884_);
  nor (_33890_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_33892_, _33890_, _05397_);
  or (_43556_, _33892_, _33889_);
  nor (_33893_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_33894_, _33893_, _05397_);
  and (_33895_, _11461_, \oc8051_golden_model_1.P1 [4]);
  and (_33896_, _31484_, _05455_);
  or (_33897_, _33896_, _33895_);
  and (_33898_, _33897_, _04018_);
  and (_33899_, _06456_, _05455_);
  or (_33900_, _33899_, _33895_);
  or (_33902_, _33900_, _04778_);
  and (_33903_, _31492_, _05455_);
  or (_33904_, _33903_, _33895_);
  or (_33905_, _33904_, _04722_);
  and (_33906_, _05455_, \oc8051_golden_model_1.ACC [4]);
  or (_33907_, _33906_, _33895_);
  and (_33908_, _33907_, _04707_);
  and (_33909_, _04708_, \oc8051_golden_model_1.P1 [4]);
  or (_33910_, _33909_, _03850_);
  or (_33911_, _33910_, _33908_);
  and (_33913_, _33911_, _03764_);
  and (_33914_, _33913_, _33905_);
  and (_33915_, _11469_, \oc8051_golden_model_1.P1 [4]);
  and (_33916_, _31520_, _06114_);
  or (_33917_, _33916_, _33915_);
  and (_33918_, _33917_, _03763_);
  or (_33919_, _33918_, _03848_);
  or (_33920_, _33919_, _33914_);
  and (_33921_, _05950_, _05455_);
  or (_33922_, _33921_, _33895_);
  or (_33924_, _33922_, _04733_);
  and (_33925_, _33924_, _33920_);
  or (_33926_, _33925_, _03854_);
  or (_33927_, _33907_, _03855_);
  and (_33928_, _33927_, _03760_);
  and (_33929_, _33928_, _33926_);
  and (_33930_, _31535_, _06114_);
  or (_33931_, _33930_, _33915_);
  and (_33932_, _33931_, _03759_);
  or (_33933_, _33932_, _03752_);
  or (_33935_, _33933_, _33929_);
  or (_33936_, _33915_, _31542_);
  and (_33937_, _33936_, _33917_);
  or (_33938_, _33937_, _03753_);
  and (_33939_, _33938_, _03747_);
  and (_33940_, _33939_, _33935_);
  and (_33941_, _31548_, _06114_);
  or (_33942_, _33941_, _33915_);
  and (_33943_, _33942_, _03746_);
  or (_33944_, _33943_, _07927_);
  or (_33946_, _33944_, _33940_);
  and (_33947_, _06969_, _05455_);
  or (_33948_, _33895_, _03738_);
  or (_33949_, _33948_, _33947_);
  or (_33950_, _33922_, _07925_);
  and (_33951_, _33950_, _03820_);
  and (_33952_, _33951_, _33949_);
  and (_33953_, _33952_, _33946_);
  and (_33954_, _31578_, _05455_);
  or (_33955_, _33954_, _33895_);
  and (_33957_, _33955_, _03455_);
  or (_33958_, _33957_, _03903_);
  or (_33959_, _33958_, _33953_);
  and (_33960_, _33959_, _33902_);
  or (_33961_, _33960_, _03897_);
  and (_33962_, _31589_, _05455_);
  or (_33963_, _33895_, _04790_);
  or (_33964_, _33963_, _33962_);
  and (_33965_, _33964_, _04792_);
  and (_33966_, _33965_, _33961_);
  or (_33968_, _33966_, _33898_);
  and (_33969_, _33968_, _03909_);
  or (_33970_, _33895_, _11238_);
  and (_33971_, _33900_, _03908_);
  and (_33972_, _33971_, _33970_);
  or (_33973_, _33972_, _33969_);
  and (_33974_, _33973_, _04785_);
  and (_33975_, _33907_, _04027_);
  and (_33976_, _33975_, _33970_);
  or (_33977_, _33976_, _03914_);
  or (_33979_, _33977_, _33974_);
  and (_33980_, _31587_, _05455_);
  or (_33981_, _33895_, _06567_);
  or (_33982_, _33981_, _33980_);
  and (_33983_, _33982_, _06572_);
  and (_33984_, _33983_, _33979_);
  and (_33985_, _31481_, _05455_);
  or (_33986_, _33985_, _33895_);
  and (_33987_, _33986_, _04011_);
  or (_33988_, _33987_, _03773_);
  or (_33990_, _33988_, _33984_);
  or (_33991_, _33904_, _03774_);
  and (_33992_, _33991_, _03375_);
  and (_33993_, _33992_, _33990_);
  and (_33994_, _33931_, _03374_);
  or (_33995_, _33994_, _03772_);
  or (_33996_, _33995_, _33993_);
  and (_33997_, _31627_, _05455_);
  or (_33998_, _33895_, _04060_);
  or (_33999_, _33998_, _33997_);
  and (_34001_, _33999_, _43152_);
  and (_34002_, _34001_, _33996_);
  or (_43557_, _34002_, _33894_);
  and (_34003_, _11461_, \oc8051_golden_model_1.P1 [5]);
  and (_34004_, _31637_, _05455_);
  or (_34005_, _34004_, _34003_);
  and (_34006_, _34005_, _04018_);
  and (_34007_, _06447_, _05455_);
  or (_34008_, _34007_, _34003_);
  or (_34009_, _34008_, _04778_);
  and (_34011_, _31645_, _05455_);
  or (_34012_, _34011_, _34003_);
  or (_34013_, _34012_, _04722_);
  and (_34014_, _05455_, \oc8051_golden_model_1.ACC [5]);
  or (_34015_, _34014_, _34003_);
  and (_34016_, _34015_, _04707_);
  and (_34017_, _04708_, \oc8051_golden_model_1.P1 [5]);
  or (_34018_, _34017_, _03850_);
  or (_34019_, _34018_, _34016_);
  and (_34020_, _34019_, _03764_);
  and (_34022_, _34020_, _34013_);
  and (_34023_, _11469_, \oc8051_golden_model_1.P1 [5]);
  and (_34024_, _31671_, _06114_);
  or (_34025_, _34024_, _34023_);
  and (_34026_, _34025_, _03763_);
  or (_34027_, _34026_, _03848_);
  or (_34028_, _34027_, _34022_);
  and (_34029_, _05857_, _05455_);
  or (_34030_, _34029_, _34003_);
  or (_34031_, _34030_, _04733_);
  and (_34033_, _34031_, _34028_);
  or (_34034_, _34033_, _03854_);
  or (_34035_, _34015_, _03855_);
  and (_34036_, _34035_, _03760_);
  and (_34037_, _34036_, _34034_);
  and (_34038_, _31686_, _06114_);
  or (_34039_, _34038_, _34023_);
  and (_34040_, _34039_, _03759_);
  or (_34041_, _34040_, _03752_);
  or (_34042_, _34041_, _34037_);
  or (_34044_, _34023_, _31693_);
  and (_34045_, _34044_, _34025_);
  or (_34046_, _34045_, _03753_);
  and (_34047_, _34046_, _03747_);
  and (_34048_, _34047_, _34042_);
  and (_34049_, _31699_, _06114_);
  or (_34050_, _34049_, _34023_);
  and (_34051_, _34050_, _03746_);
  or (_34052_, _34051_, _08474_);
  or (_34053_, _34052_, _34048_);
  or (_34054_, _34030_, _07925_);
  and (_34055_, _34054_, _34053_);
  or (_34056_, _34055_, _03737_);
  and (_34057_, _06968_, _05455_);
  or (_34058_, _34003_, _03738_);
  or (_34059_, _34058_, _34057_);
  and (_34060_, _34059_, _03820_);
  and (_34061_, _34060_, _34056_);
  and (_34062_, _31727_, _05455_);
  or (_34063_, _34062_, _34003_);
  and (_34066_, _34063_, _03455_);
  or (_34067_, _34066_, _03903_);
  or (_34068_, _34067_, _34061_);
  and (_34069_, _34068_, _34009_);
  or (_34070_, _34069_, _03897_);
  and (_34071_, _31738_, _05455_);
  or (_34072_, _34071_, _34003_);
  or (_34073_, _34072_, _04790_);
  and (_34074_, _34073_, _04792_);
  and (_34075_, _34074_, _34070_);
  or (_34077_, _34075_, _34006_);
  and (_34078_, _34077_, _03909_);
  or (_34079_, _34003_, _11237_);
  and (_34080_, _34008_, _03908_);
  and (_34081_, _34080_, _34079_);
  or (_34082_, _34081_, _34078_);
  and (_34083_, _34082_, _04785_);
  and (_34084_, _34015_, _04027_);
  and (_34085_, _34084_, _34079_);
  or (_34086_, _34085_, _03914_);
  or (_34088_, _34086_, _34083_);
  and (_34089_, _31736_, _05455_);
  or (_34090_, _34003_, _06567_);
  or (_34091_, _34090_, _34089_);
  and (_34092_, _34091_, _06572_);
  and (_34093_, _34092_, _34088_);
  and (_34094_, _31634_, _05455_);
  or (_34095_, _34094_, _34003_);
  and (_34096_, _34095_, _04011_);
  or (_34097_, _34096_, _03773_);
  or (_34099_, _34097_, _34093_);
  or (_34100_, _34012_, _03774_);
  and (_34101_, _34100_, _03375_);
  and (_34102_, _34101_, _34099_);
  and (_34103_, _34039_, _03374_);
  or (_34104_, _34103_, _03772_);
  or (_34105_, _34104_, _34102_);
  and (_34106_, _31775_, _05455_);
  or (_34107_, _34003_, _04060_);
  or (_34108_, _34107_, _34106_);
  and (_34110_, _34108_, _43152_);
  and (_34111_, _34110_, _34105_);
  nor (_34112_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_34113_, _34112_, _05397_);
  or (_43558_, _34113_, _34111_);
  and (_34114_, _11461_, \oc8051_golden_model_1.P1 [6]);
  and (_34115_, _31787_, _05455_);
  or (_34116_, _34115_, _34114_);
  and (_34117_, _34116_, _04018_);
  and (_34118_, _13394_, _05455_);
  or (_34120_, _34118_, _34114_);
  or (_34121_, _34120_, _04778_);
  and (_34122_, _11469_, \oc8051_golden_model_1.P1 [6]);
  and (_34123_, _31807_, _06114_);
  or (_34124_, _34123_, _34122_);
  and (_34125_, _34124_, _03759_);
  and (_34126_, _31813_, _05455_);
  or (_34127_, _34126_, _34114_);
  or (_34128_, _34127_, _04722_);
  and (_34129_, _05455_, \oc8051_golden_model_1.ACC [6]);
  or (_34131_, _34129_, _34114_);
  and (_34132_, _34131_, _04707_);
  and (_34133_, _04708_, \oc8051_golden_model_1.P1 [6]);
  or (_34134_, _34133_, _03850_);
  or (_34135_, _34134_, _34132_);
  and (_34136_, _34135_, _03764_);
  and (_34137_, _34136_, _34128_);
  and (_34138_, _31826_, _06114_);
  or (_34139_, _34138_, _34122_);
  and (_34140_, _34139_, _03763_);
  or (_34142_, _34140_, _03848_);
  or (_34143_, _34142_, _34137_);
  and (_34144_, _06065_, _05455_);
  or (_34145_, _34144_, _34114_);
  or (_34146_, _34145_, _04733_);
  and (_34147_, _34146_, _34143_);
  or (_34148_, _34147_, _03854_);
  or (_34149_, _34131_, _03855_);
  and (_34150_, _34149_, _03760_);
  and (_34151_, _34150_, _34148_);
  or (_34153_, _34151_, _34125_);
  and (_34154_, _34153_, _03753_);
  or (_34155_, _34122_, _31843_);
  and (_34156_, _34139_, _03752_);
  and (_34157_, _34156_, _34155_);
  or (_34158_, _34157_, _34154_);
  and (_34159_, _34158_, _03747_);
  and (_34160_, _31850_, _06114_);
  or (_34161_, _34160_, _34122_);
  and (_34162_, _34161_, _03746_);
  or (_34164_, _34162_, _07927_);
  or (_34165_, _34164_, _34159_);
  and (_34166_, _06641_, _05455_);
  or (_34167_, _34114_, _03738_);
  or (_34168_, _34167_, _34166_);
  or (_34169_, _34145_, _07925_);
  and (_34170_, _34169_, _03820_);
  and (_34171_, _34170_, _34168_);
  and (_34172_, _34171_, _34165_);
  and (_34173_, _31876_, _05455_);
  or (_34175_, _34173_, _34114_);
  and (_34176_, _34175_, _03455_);
  or (_34177_, _34176_, _03903_);
  or (_34178_, _34177_, _34172_);
  and (_34179_, _34178_, _34121_);
  or (_34180_, _34179_, _03897_);
  and (_34181_, _31887_, _05455_);
  or (_34182_, _34114_, _04790_);
  or (_34183_, _34182_, _34181_);
  and (_34184_, _34183_, _04792_);
  and (_34186_, _34184_, _34180_);
  or (_34187_, _34186_, _34117_);
  and (_34188_, _34187_, _03909_);
  or (_34189_, _34114_, _11236_);
  and (_34190_, _34120_, _03908_);
  and (_34191_, _34190_, _34189_);
  or (_34192_, _34191_, _34188_);
  and (_34193_, _34192_, _04785_);
  and (_34194_, _34131_, _04027_);
  and (_34195_, _34194_, _34189_);
  or (_34197_, _34195_, _03914_);
  or (_34198_, _34197_, _34193_);
  and (_34199_, _31885_, _05455_);
  or (_34200_, _34114_, _06567_);
  or (_34201_, _34200_, _34199_);
  and (_34202_, _34201_, _06572_);
  and (_34203_, _34202_, _34198_);
  and (_34204_, _31785_, _05455_);
  or (_34205_, _34204_, _34114_);
  and (_34206_, _34205_, _04011_);
  or (_34208_, _34206_, _03773_);
  or (_34209_, _34208_, _34203_);
  or (_34210_, _34127_, _03774_);
  and (_34211_, _34210_, _03375_);
  and (_34212_, _34211_, _34209_);
  and (_34213_, _34124_, _03374_);
  or (_34214_, _34213_, _03772_);
  or (_34215_, _34214_, _34212_);
  and (_34216_, _31925_, _05455_);
  or (_34217_, _34114_, _04060_);
  or (_34219_, _34217_, _34216_);
  and (_34220_, _34219_, _43152_);
  and (_34221_, _34220_, _34215_);
  nor (_34222_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_34223_, _34222_, _05397_);
  or (_43559_, _34223_, _34221_);
  and (_34224_, _05516_, _04700_);
  nor (_34225_, _05516_, _03683_);
  or (_34226_, _34225_, _07925_);
  or (_34227_, _34226_, _34224_);
  and (_34229_, _05716_, _05516_);
  or (_34230_, _34229_, _34225_);
  or (_34231_, _34230_, _04722_);
  and (_34232_, _05516_, \oc8051_golden_model_1.ACC [0]);
  or (_34233_, _34232_, _34225_);
  and (_34234_, _34233_, _04707_);
  nor (_34235_, _04707_, _03683_);
  or (_34236_, _34235_, _03850_);
  or (_34237_, _34236_, _34234_);
  and (_34238_, _34237_, _04733_);
  and (_34240_, _34238_, _34231_);
  or (_34241_, _04288_, _03854_);
  or (_34242_, _34241_, _34240_);
  or (_34243_, _34233_, _03855_);
  and (_34244_, _34243_, _04845_);
  and (_34245_, _34244_, _34242_);
  nand (_34246_, _07925_, _04750_);
  or (_34247_, _34246_, _34245_);
  and (_34248_, _34247_, _34227_);
  or (_34249_, _34248_, _03737_);
  and (_34251_, _06962_, _05516_);
  or (_34252_, _34225_, _03738_);
  or (_34253_, _34252_, _34251_);
  and (_34254_, _34253_, _34249_);
  or (_34255_, _34254_, _03455_);
  nor (_34256_, _12164_, _11630_);
  or (_34257_, _34225_, _03820_);
  or (_34258_, _34257_, _34256_);
  and (_34259_, _34258_, _04778_);
  and (_34260_, _34259_, _34255_);
  and (_34262_, _05516_, _06479_);
  or (_34263_, _34262_, _34225_);
  and (_34264_, _34263_, _03903_);
  or (_34265_, _34264_, _03897_);
  or (_34266_, _34265_, _34260_);
  and (_34267_, _12178_, _05516_);
  or (_34268_, _34225_, _04790_);
  or (_34269_, _34268_, _34267_);
  and (_34270_, _34269_, _04792_);
  and (_34271_, _34270_, _34266_);
  nor (_34273_, _10488_, _11630_);
  or (_34274_, _34273_, _34225_);
  nand (_34275_, _08753_, _05516_);
  and (_34276_, _34275_, _04018_);
  and (_34277_, _34276_, _34274_);
  or (_34278_, _34277_, _34271_);
  and (_34279_, _34278_, _03909_);
  nand (_34280_, _34263_, _03908_);
  nor (_34281_, _34280_, _34229_);
  or (_34282_, _34281_, _04027_);
  or (_34283_, _34282_, _34279_);
  nor (_34284_, _34225_, _04785_);
  nand (_34285_, _34284_, _34275_);
  and (_34286_, _34285_, _34283_);
  or (_34287_, _34286_, _03914_);
  nor (_34288_, _12177_, _11630_);
  or (_34289_, _34225_, _06567_);
  or (_34290_, _34289_, _34288_);
  and (_34291_, _34290_, _06572_);
  and (_34292_, _34291_, _34287_);
  and (_34294_, _34274_, _04011_);
  or (_34295_, _34294_, _17157_);
  or (_34296_, _34295_, _34292_);
  or (_34297_, _34230_, _04144_);
  and (_34298_, _34297_, _43152_);
  and (_34299_, _34298_, _34296_);
  nor (_34300_, _43152_, _03683_);
  or (_34301_, _34300_, rst);
  or (_43562_, _34301_, _34299_);
  nor (_34302_, _05516_, _04605_);
  and (_34304_, _12262_, _05516_);
  or (_34305_, _34304_, _34302_);
  and (_34306_, _34305_, _03772_);
  not (_34307_, _34304_);
  or (_34308_, _05516_, \oc8051_golden_model_1.SP [1]);
  and (_34309_, _34308_, _34307_);
  or (_34310_, _34309_, _04722_);
  nand (_34311_, _03768_, \oc8051_golden_model_1.SP [1]);
  and (_34312_, _05516_, \oc8051_golden_model_1.ACC [1]);
  or (_34313_, _34312_, _34302_);
  and (_34315_, _34313_, _04707_);
  nor (_34316_, _04707_, _04605_);
  or (_34317_, _34316_, _03768_);
  or (_34318_, _34317_, _34315_);
  and (_34319_, _34318_, _34311_);
  or (_34320_, _34319_, _03850_);
  and (_34321_, _34320_, _03431_);
  and (_34322_, _34321_, _34310_);
  nor (_34323_, _03431_, \oc8051_golden_model_1.SP [1]);
  or (_34324_, _34323_, _03848_);
  or (_34326_, _34324_, _34322_);
  nand (_34327_, _04840_, _03848_);
  and (_34328_, _34327_, _34326_);
  or (_34329_, _34328_, _03854_);
  or (_34330_, _34313_, _03855_);
  and (_34331_, _34330_, _04845_);
  and (_34332_, _34331_, _34329_);
  not (_34333_, _05050_);
  or (_34334_, _34333_, _04844_);
  or (_34335_, _34334_, _34332_);
  or (_34337_, _05050_, _04605_);
  and (_34338_, _34337_, _07925_);
  and (_34339_, _34338_, _34335_);
  or (_34340_, _11630_, _04900_);
  and (_34341_, _34308_, _08474_);
  and (_34342_, _34341_, _34340_);
  or (_34343_, _34342_, _03737_);
  or (_34344_, _34343_, _34339_);
  and (_34345_, _06961_, _05516_);
  or (_34346_, _34302_, _03738_);
  or (_34348_, _34346_, _34345_);
  and (_34349_, _34348_, _03820_);
  and (_34350_, _34349_, _34344_);
  nor (_34351_, _12352_, _11630_);
  or (_34352_, _34351_, _34302_);
  and (_34353_, _34352_, _03455_);
  or (_34354_, _34353_, _34350_);
  and (_34355_, _34354_, _04778_);
  nand (_34356_, _05516_, _04595_);
  and (_34357_, _34308_, _03903_);
  and (_34359_, _34357_, _34356_);
  or (_34360_, _34359_, _03401_);
  or (_34361_, _34360_, _34355_);
  nand (_34362_, _03401_, \oc8051_golden_model_1.SP [1]);
  and (_34363_, _34362_, _04790_);
  and (_34364_, _34363_, _34361_);
  or (_34365_, _12366_, _11630_);
  and (_34366_, _34308_, _03897_);
  and (_34367_, _34366_, _34365_);
  or (_34368_, _34367_, _04018_);
  or (_34370_, _34368_, _34364_);
  nor (_34371_, _08751_, _11630_);
  or (_34372_, _34371_, _34302_);
  nand (_34373_, _08750_, _05516_);
  and (_34374_, _34373_, _34372_);
  or (_34375_, _34374_, _04792_);
  and (_34376_, _34375_, _03909_);
  and (_34377_, _34376_, _34370_);
  or (_34378_, _12244_, _11630_);
  and (_34379_, _34308_, _03908_);
  and (_34381_, _34379_, _34378_);
  or (_34382_, _34381_, _04027_);
  or (_34383_, _34382_, _34377_);
  nor (_34384_, _34302_, _04785_);
  nand (_34385_, _34384_, _34373_);
  and (_34386_, _34385_, _34383_);
  or (_34387_, _34386_, _03388_);
  nand (_34388_, _03388_, \oc8051_golden_model_1.SP [1]);
  and (_34389_, _34388_, _06567_);
  and (_34390_, _34389_, _34387_);
  or (_34392_, _34356_, _08366_);
  and (_34393_, _34308_, _03914_);
  and (_34394_, _34393_, _34392_);
  or (_34395_, _34394_, _34390_);
  and (_34396_, _34395_, _06572_);
  and (_34397_, _34372_, _04011_);
  or (_34398_, _34397_, _04034_);
  nor (_34399_, _34398_, _34396_);
  or (_34400_, _34399_, _04618_);
  nor (_34401_, _03777_, _03383_);
  nand (_34403_, _34401_, _34400_);
  or (_34404_, _34401_, _04605_);
  and (_34405_, _34404_, _03774_);
  and (_34406_, _34405_, _34403_);
  and (_34407_, _34309_, _03773_);
  or (_34408_, _34407_, _05223_);
  or (_34409_, _34408_, _34406_);
  or (_34410_, _04819_, _04605_);
  and (_34411_, _34410_, _04060_);
  and (_34412_, _34411_, _34409_);
  or (_34414_, _34412_, _34306_);
  and (_34415_, _34414_, _43152_);
  nor (_34416_, \oc8051_golden_model_1.SP [1], rst);
  nor (_34417_, _34416_, _00000_);
  or (_43563_, _34417_, _34415_);
  nor (_34418_, _43152_, _04182_);
  or (_34419_, _34418_, rst);
  nand (_34420_, _13842_, _03401_);
  and (_34421_, _05516_, _05307_);
  nor (_34422_, _05516_, _04182_);
  or (_34424_, _34422_, _07925_);
  or (_34425_, _34424_, _34421_);
  nor (_34426_, _12471_, _11630_);
  or (_34427_, _34426_, _34422_);
  or (_34428_, _34427_, _04722_);
  and (_34429_, _05516_, \oc8051_golden_model_1.ACC [2]);
  or (_34430_, _34429_, _34422_);
  or (_34431_, _34430_, _04708_);
  or (_34432_, _04707_, \oc8051_golden_model_1.SP [2]);
  and (_34433_, _34432_, _03770_);
  and (_34435_, _34433_, _34431_);
  and (_34436_, _05393_, _03768_);
  or (_34437_, _34436_, _03850_);
  or (_34438_, _34437_, _34435_);
  and (_34439_, _34438_, _03431_);
  and (_34440_, _34439_, _34428_);
  nor (_34441_, _13842_, _03431_);
  or (_34442_, _34441_, _03848_);
  or (_34443_, _34442_, _34440_);
  nand (_34444_, _06178_, _03848_);
  and (_34446_, _34444_, _34443_);
  or (_34447_, _34446_, _03854_);
  or (_34448_, _34430_, _03855_);
  and (_34449_, _34448_, _04845_);
  and (_34450_, _34449_, _34447_);
  or (_34451_, _05253_, _05049_);
  or (_34452_, _34451_, _34450_);
  nor (_34453_, _05393_, _03428_);
  nor (_34454_, _34453_, _03456_);
  and (_34455_, _34454_, _34452_);
  nand (_34457_, _05393_, _03456_);
  nand (_34458_, _34457_, _07925_);
  or (_34459_, _34458_, _34455_);
  and (_34460_, _34459_, _34425_);
  or (_34461_, _34460_, _03737_);
  and (_34462_, _06965_, _05516_);
  or (_34463_, _34422_, _03738_);
  or (_34464_, _34463_, _34462_);
  and (_34465_, _34464_, _03820_);
  and (_34466_, _34465_, _34461_);
  nor (_34468_, _12572_, _11630_);
  or (_34469_, _34468_, _34422_);
  and (_34470_, _34469_, _03455_);
  or (_34471_, _34470_, _03903_);
  or (_34472_, _34471_, _34466_);
  and (_34473_, _05516_, _06495_);
  or (_34474_, _34473_, _34422_);
  or (_34475_, _34474_, _04778_);
  and (_34476_, _34475_, _34472_);
  or (_34477_, _34476_, _03401_);
  and (_34479_, _34477_, _34420_);
  or (_34480_, _34479_, _03897_);
  and (_34481_, _12586_, _05516_);
  or (_34482_, _34422_, _04790_);
  or (_34483_, _34482_, _34481_);
  and (_34484_, _34483_, _04792_);
  and (_34485_, _34484_, _34480_);
  and (_34486_, _08748_, _05516_);
  or (_34487_, _34486_, _34422_);
  and (_34488_, _34487_, _04018_);
  or (_34490_, _34488_, _34485_);
  and (_34491_, _34490_, _03909_);
  or (_34492_, _34422_, _05765_);
  and (_34493_, _34474_, _03908_);
  and (_34494_, _34493_, _34492_);
  or (_34495_, _34494_, _34491_);
  and (_34496_, _34495_, _10076_);
  and (_34497_, _34430_, _04027_);
  and (_34498_, _34497_, _34492_);
  and (_34499_, _05393_, _03388_);
  or (_34501_, _34499_, _03914_);
  or (_34502_, _34501_, _34498_);
  or (_34503_, _34502_, _34496_);
  nor (_34504_, _12585_, _11630_);
  or (_34505_, _34422_, _06567_);
  or (_34506_, _34505_, _34504_);
  and (_34507_, _34506_, _34503_);
  or (_34508_, _34507_, _04011_);
  nor (_34509_, _08747_, _11630_);
  or (_34510_, _34509_, _34422_);
  or (_34512_, _34510_, _06572_);
  and (_34513_, _34512_, _10704_);
  and (_34514_, _34513_, _34508_);
  and (_34515_, _13842_, _04034_);
  or (_34516_, _34515_, _03383_);
  or (_34517_, _34516_, _34514_);
  nand (_34518_, _13842_, _03383_);
  and (_34519_, _34518_, _03778_);
  and (_34520_, _34519_, _34517_);
  and (_34521_, _13842_, _03777_);
  or (_34523_, _34521_, _03773_);
  or (_34524_, _34523_, _34520_);
  or (_34525_, _34427_, _03774_);
  and (_34526_, _34525_, _04819_);
  and (_34527_, _34526_, _34524_);
  nor (_34528_, _13842_, _04819_);
  or (_34529_, _34528_, _03772_);
  or (_34530_, _34529_, _34527_);
  and (_34531_, _12642_, _05516_);
  or (_34532_, _34422_, _04060_);
  or (_34534_, _34532_, _34531_);
  and (_34535_, _34534_, _43152_);
  and (_34536_, _34535_, _34530_);
  or (_43564_, _34536_, _34419_);
  nor (_34537_, _43152_, _03847_);
  or (_34538_, _05396_, _04819_);
  nand (_34539_, _13648_, _03383_);
  or (_34540_, _05396_, _05050_);
  nor (_34541_, _05516_, _03847_);
  nor (_34542_, _12681_, _11630_);
  or (_34544_, _34542_, _34541_);
  or (_34545_, _34544_, _04722_);
  and (_34546_, _05516_, \oc8051_golden_model_1.ACC [3]);
  or (_34547_, _34546_, _34541_);
  or (_34548_, _34547_, _04708_);
  or (_34549_, _04707_, \oc8051_golden_model_1.SP [3]);
  and (_34550_, _34549_, _03770_);
  and (_34551_, _34550_, _34548_);
  and (_34552_, _05396_, _03768_);
  or (_34553_, _34552_, _03850_);
  or (_34555_, _34553_, _34551_);
  and (_34556_, _34555_, _03431_);
  and (_34557_, _34556_, _34545_);
  nor (_34558_, _13648_, _03431_);
  or (_34559_, _34558_, _03848_);
  or (_34560_, _34559_, _34557_);
  nand (_34561_, _06168_, _03848_);
  and (_34562_, _34561_, _34560_);
  or (_34563_, _34562_, _03854_);
  or (_34564_, _34547_, _03855_);
  and (_34566_, _34564_, _04845_);
  and (_34567_, _34566_, _34563_);
  or (_34568_, _05173_, _34333_);
  or (_34569_, _34568_, _34567_);
  and (_34570_, _34569_, _34540_);
  or (_34571_, _34570_, _07927_);
  and (_34572_, _06964_, _05516_);
  or (_34573_, _34541_, _03738_);
  or (_34574_, _34573_, _34572_);
  and (_34575_, _05516_, _05119_);
  or (_34577_, _34541_, _07925_);
  or (_34578_, _34577_, _34575_);
  and (_34579_, _34578_, _03820_);
  and (_34580_, _34579_, _34574_);
  and (_34581_, _34580_, _34571_);
  nor (_34582_, _12775_, _11630_);
  or (_34583_, _34582_, _34541_);
  and (_34584_, _34583_, _03455_);
  or (_34585_, _34584_, _03903_);
  or (_34586_, _34585_, _34581_);
  and (_34588_, _05516_, _06345_);
  or (_34589_, _34588_, _34541_);
  or (_34590_, _34589_, _04778_);
  and (_34591_, _34590_, _11641_);
  and (_34592_, _34591_, _34586_);
  and (_34593_, _05396_, _03401_);
  or (_34594_, _34593_, _03897_);
  or (_34595_, _34594_, _34592_);
  and (_34596_, _12789_, _05516_);
  or (_34597_, _34541_, _04790_);
  or (_34599_, _34597_, _34596_);
  and (_34600_, _34599_, _04792_);
  and (_34601_, _34600_, _34595_);
  and (_34602_, _10491_, _05516_);
  or (_34603_, _34602_, _34541_);
  and (_34604_, _34603_, _04018_);
  or (_34605_, _34604_, _34601_);
  and (_34606_, _34605_, _03909_);
  or (_34607_, _34541_, _05622_);
  and (_34608_, _34589_, _03908_);
  and (_34610_, _34608_, _34607_);
  or (_34611_, _34610_, _34606_);
  and (_34612_, _34611_, _10076_);
  and (_34613_, _34547_, _04027_);
  and (_34614_, _34613_, _34607_);
  and (_34615_, _05396_, _03388_);
  or (_34616_, _34615_, _03914_);
  or (_34617_, _34616_, _34614_);
  or (_34618_, _34617_, _34612_);
  nor (_34619_, _12788_, _11630_);
  or (_34621_, _34619_, _34541_);
  or (_34622_, _34621_, _06567_);
  and (_34623_, _34622_, _34618_);
  or (_34624_, _34623_, _04011_);
  nor (_34625_, _08742_, _11630_);
  or (_34626_, _34625_, _34541_);
  or (_34627_, _34626_, _06572_);
  and (_34628_, _34627_, _10704_);
  and (_34629_, _34628_, _34624_);
  nor (_34630_, _06165_, _03847_);
  or (_34632_, _34630_, _06166_);
  and (_34633_, _34632_, _04034_);
  or (_34634_, _34633_, _03383_);
  or (_34635_, _34634_, _34629_);
  and (_34636_, _34635_, _34539_);
  or (_34637_, _34636_, _03777_);
  or (_34638_, _34632_, _03778_);
  and (_34639_, _34638_, _03774_);
  and (_34640_, _34639_, _34637_);
  and (_34641_, _34544_, _03773_);
  or (_34643_, _34641_, _05223_);
  or (_34644_, _34643_, _34640_);
  and (_34645_, _34644_, _34538_);
  or (_34646_, _34645_, _03772_);
  and (_34647_, _12848_, _05516_);
  or (_34648_, _34541_, _04060_);
  or (_34649_, _34648_, _34647_);
  and (_34650_, _34649_, _43152_);
  and (_34651_, _34650_, _34646_);
  or (_34652_, _34651_, _34537_);
  and (_43567_, _34652_, _41894_);
  nor (_34654_, _43152_, _11599_);
  nor (_34655_, _05127_, \oc8051_golden_model_1.SP [4]);
  nor (_34656_, _34655_, _11565_);
  or (_34657_, _34656_, _04819_);
  or (_34658_, _34656_, _03384_);
  or (_34659_, _34656_, _05050_);
  nor (_34660_, _05516_, _11599_);
  nor (_34661_, _12891_, _11630_);
  or (_34662_, _34661_, _34660_);
  or (_34664_, _34662_, _04722_);
  and (_34665_, _05516_, \oc8051_golden_model_1.ACC [4]);
  or (_34666_, _34665_, _34660_);
  or (_34667_, _34666_, _04708_);
  or (_34668_, _04707_, \oc8051_golden_model_1.SP [4]);
  and (_34669_, _34668_, _03770_);
  and (_34670_, _34669_, _34667_);
  and (_34671_, _34656_, _03768_);
  or (_34672_, _34671_, _03850_);
  or (_34673_, _34672_, _34670_);
  and (_34674_, _34673_, _03431_);
  and (_34675_, _34674_, _34664_);
  and (_34676_, _34656_, _05045_);
  or (_34677_, _34676_, _03848_);
  or (_34678_, _34677_, _34675_);
  and (_34679_, _11600_, _03683_);
  nor (_34680_, _06167_, _11599_);
  nor (_34681_, _34680_, _34679_);
  nand (_34682_, _34681_, _03848_);
  and (_34683_, _34682_, _34678_);
  or (_34686_, _34683_, _03854_);
  or (_34687_, _34666_, _03855_);
  and (_34688_, _34687_, _04845_);
  and (_34689_, _34688_, _34686_);
  and (_34690_, _05128_, \oc8051_golden_model_1.SP [4]);
  nor (_34691_, _05128_, \oc8051_golden_model_1.SP [4]);
  nor (_34692_, _34691_, _34690_);
  nand (_34693_, _34692_, _03758_);
  nand (_34694_, _34693_, _05050_);
  or (_34695_, _34694_, _34689_);
  and (_34697_, _34695_, _34659_);
  or (_34698_, _34697_, _08474_);
  and (_34699_, _05950_, _05516_);
  or (_34700_, _34660_, _07925_);
  or (_34701_, _34700_, _34699_);
  and (_34702_, _34701_, _34698_);
  or (_34703_, _34702_, _03737_);
  and (_34704_, _06969_, _05516_);
  or (_34705_, _34660_, _03738_);
  or (_34706_, _34705_, _34704_);
  and (_34708_, _34706_, _34703_);
  or (_34709_, _34708_, _03455_);
  nor (_34710_, _12982_, _11630_);
  or (_34711_, _34660_, _03820_);
  or (_34712_, _34711_, _34710_);
  and (_34713_, _34712_, _04778_);
  and (_34714_, _34713_, _34709_);
  and (_34715_, _06456_, _05516_);
  or (_34716_, _34715_, _34660_);
  and (_34717_, _34716_, _03903_);
  or (_34719_, _34717_, _03401_);
  or (_34720_, _34719_, _34714_);
  or (_34721_, _34656_, _11641_);
  and (_34722_, _34721_, _34720_);
  or (_34723_, _34722_, _03897_);
  and (_34724_, _12997_, _05516_);
  or (_34725_, _34660_, _04790_);
  or (_34726_, _34725_, _34724_);
  and (_34727_, _34726_, _04792_);
  and (_34728_, _34727_, _34723_);
  and (_34730_, _08741_, _05516_);
  or (_34731_, _34730_, _34660_);
  and (_34732_, _34731_, _04018_);
  or (_34733_, _34732_, _34728_);
  and (_34734_, _34733_, _03909_);
  or (_34735_, _34660_, _08336_);
  and (_34736_, _34716_, _03908_);
  and (_34737_, _34736_, _34735_);
  or (_34738_, _34737_, _34734_);
  and (_34739_, _34738_, _10076_);
  and (_34741_, _34666_, _04027_);
  and (_34742_, _34741_, _34735_);
  and (_34743_, _34656_, _03388_);
  or (_34744_, _34743_, _03914_);
  or (_34745_, _34744_, _34742_);
  or (_34746_, _34745_, _34739_);
  nor (_34747_, _12996_, _11630_);
  or (_34748_, _34660_, _06567_);
  or (_34749_, _34748_, _34747_);
  and (_34750_, _34749_, _34746_);
  or (_34752_, _34750_, _04011_);
  nor (_34753_, _08740_, _11630_);
  or (_34754_, _34753_, _34660_);
  or (_34755_, _34754_, _06572_);
  and (_34756_, _34755_, _10704_);
  and (_34757_, _34756_, _34752_);
  nor (_34758_, _06166_, _11599_);
  or (_34759_, _34758_, _11600_);
  and (_34760_, _34759_, _04034_);
  or (_34761_, _34760_, _03383_);
  or (_34763_, _34761_, _34757_);
  and (_34764_, _34763_, _34658_);
  or (_34765_, _34764_, _03777_);
  or (_34766_, _34759_, _03778_);
  and (_34767_, _34766_, _03774_);
  and (_34768_, _34767_, _34765_);
  and (_34769_, _34662_, _03773_);
  or (_34770_, _34769_, _05223_);
  or (_34771_, _34770_, _34768_);
  and (_34772_, _34771_, _34657_);
  or (_34774_, _34772_, _03772_);
  and (_34775_, _13056_, _05516_);
  or (_34776_, _34660_, _04060_);
  or (_34777_, _34776_, _34775_);
  and (_34778_, _34777_, _43152_);
  and (_34779_, _34778_, _34774_);
  or (_34780_, _34779_, _34654_);
  and (_43568_, _34780_, _41894_);
  nor (_34781_, _43152_, _11598_);
  nor (_34782_, _11565_, \oc8051_golden_model_1.SP [5]);
  nor (_34784_, _34782_, _11566_);
  or (_34785_, _34784_, _04819_);
  or (_34786_, _34784_, _03384_);
  or (_34787_, _34784_, _05050_);
  nor (_34788_, _05516_, _11598_);
  nor (_34789_, _13090_, _11630_);
  or (_34790_, _34789_, _34788_);
  or (_34791_, _34790_, _04722_);
  and (_34792_, _05516_, \oc8051_golden_model_1.ACC [5]);
  or (_34793_, _34792_, _34788_);
  or (_34795_, _34793_, _04708_);
  or (_34796_, _04707_, \oc8051_golden_model_1.SP [5]);
  and (_34797_, _34796_, _03770_);
  and (_34798_, _34797_, _34795_);
  and (_34799_, _34784_, _03768_);
  or (_34800_, _34799_, _03850_);
  or (_34801_, _34800_, _34798_);
  and (_34802_, _34801_, _03431_);
  and (_34803_, _34802_, _34791_);
  and (_34804_, _34784_, _05045_);
  or (_34806_, _34804_, _03848_);
  or (_34807_, _34806_, _34803_);
  and (_34808_, _11601_, _03683_);
  nor (_34809_, _34679_, _11598_);
  nor (_34810_, _34809_, _34808_);
  nand (_34811_, _34810_, _03848_);
  and (_34812_, _34811_, _34807_);
  or (_34813_, _34812_, _03854_);
  or (_34814_, _34793_, _03855_);
  and (_34815_, _34814_, _04845_);
  and (_34817_, _34815_, _34813_);
  nor (_34818_, _34690_, \oc8051_golden_model_1.SP [5]);
  nor (_34819_, _34818_, _11613_);
  nand (_34820_, _34819_, _03758_);
  nand (_34821_, _34820_, _05050_);
  or (_34822_, _34821_, _34817_);
  and (_34823_, _34822_, _34787_);
  or (_34824_, _34823_, _08474_);
  and (_34825_, _05857_, _05516_);
  or (_34826_, _34788_, _07925_);
  or (_34828_, _34826_, _34825_);
  and (_34829_, _34828_, _34824_);
  or (_34830_, _34829_, _03737_);
  and (_34831_, _06968_, _05516_);
  or (_34832_, _34788_, _03738_);
  or (_34833_, _34832_, _34831_);
  and (_34834_, _34833_, _03820_);
  and (_34835_, _34834_, _34830_);
  nor (_34836_, _13182_, _11630_);
  or (_34837_, _34836_, _34788_);
  and (_34839_, _34837_, _03455_);
  or (_34840_, _34839_, _03903_);
  or (_34841_, _34840_, _34835_);
  and (_34842_, _06447_, _05516_);
  or (_34843_, _34842_, _34788_);
  or (_34844_, _34843_, _04778_);
  and (_34845_, _34844_, _34841_);
  or (_34846_, _34845_, _03401_);
  or (_34847_, _34784_, _11641_);
  and (_34848_, _34847_, _34846_);
  or (_34850_, _34848_, _03897_);
  and (_34851_, _13196_, _05516_);
  or (_34852_, _34788_, _04790_);
  or (_34853_, _34852_, _34851_);
  and (_34854_, _34853_, _04792_);
  and (_34855_, _34854_, _34850_);
  and (_34856_, _10493_, _05516_);
  or (_34857_, _34856_, _34788_);
  and (_34858_, _34857_, _04018_);
  or (_34859_, _34858_, _34855_);
  and (_34861_, _34859_, _03909_);
  or (_34862_, _34788_, _08335_);
  and (_34863_, _34843_, _03908_);
  and (_34864_, _34863_, _34862_);
  or (_34865_, _34864_, _34861_);
  and (_34866_, _34865_, _10076_);
  and (_34867_, _34793_, _04027_);
  and (_34868_, _34867_, _34862_);
  and (_34869_, _34784_, _03388_);
  or (_34870_, _34869_, _03914_);
  or (_34872_, _34870_, _34868_);
  or (_34873_, _34872_, _34866_);
  nor (_34874_, _13195_, _11630_);
  or (_34875_, _34788_, _06567_);
  or (_34876_, _34875_, _34874_);
  and (_34877_, _34876_, _34873_);
  or (_34878_, _34877_, _04011_);
  nor (_34879_, _08738_, _11630_);
  or (_34880_, _34879_, _34788_);
  or (_34881_, _34880_, _06572_);
  and (_34883_, _34881_, _10704_);
  and (_34884_, _34883_, _34878_);
  nor (_34885_, _11600_, _11598_);
  or (_34886_, _34885_, _11601_);
  and (_34887_, _34886_, _04034_);
  or (_34888_, _34887_, _03383_);
  or (_34889_, _34888_, _34884_);
  and (_34890_, _34889_, _34786_);
  or (_34891_, _34890_, _03777_);
  or (_34892_, _34886_, _03778_);
  and (_34894_, _34892_, _03774_);
  and (_34895_, _34894_, _34891_);
  and (_34896_, _34790_, _03773_);
  or (_34897_, _34896_, _05223_);
  or (_34898_, _34897_, _34895_);
  and (_34899_, _34898_, _34785_);
  or (_34900_, _34899_, _03772_);
  and (_34901_, _13255_, _05516_);
  or (_34902_, _34788_, _04060_);
  or (_34903_, _34902_, _34901_);
  and (_34905_, _34903_, _43152_);
  and (_34906_, _34905_, _34900_);
  or (_34907_, _34906_, _34781_);
  and (_43569_, _34907_, _41894_);
  nor (_34908_, _43152_, _11597_);
  nor (_34909_, _05516_, _11597_);
  nor (_34910_, _13293_, _11630_);
  or (_34911_, _34910_, _34909_);
  or (_34912_, _34911_, _04722_);
  and (_34913_, _05516_, \oc8051_golden_model_1.ACC [6]);
  nor (_34915_, _34913_, _34909_);
  nand (_34916_, _34915_, _04707_);
  or (_34917_, _04707_, \oc8051_golden_model_1.SP [6]);
  and (_34918_, _34917_, _03770_);
  and (_34919_, _34918_, _34916_);
  nor (_34920_, _11566_, \oc8051_golden_model_1.SP [6]);
  nor (_34921_, _34920_, _11567_);
  and (_34922_, _34921_, _03768_);
  or (_34923_, _34922_, _03850_);
  or (_34924_, _34923_, _34919_);
  and (_34926_, _34924_, _03431_);
  and (_34927_, _34926_, _34912_);
  and (_34928_, _34921_, _05045_);
  or (_34929_, _34928_, _03848_);
  or (_34930_, _34929_, _34927_);
  nor (_34931_, _34808_, _11597_);
  nor (_34932_, _34931_, _11603_);
  nand (_34933_, _34932_, _03848_);
  nand (_34934_, _34933_, _34930_);
  and (_34935_, _34934_, _03855_);
  and (_34937_, _34915_, _03854_);
  or (_34938_, _34937_, _03758_);
  or (_34939_, _34938_, _34935_);
  nor (_34940_, _11613_, \oc8051_golden_model_1.SP [6]);
  nor (_34941_, _34940_, _11614_);
  nand (_34942_, _34941_, _03758_);
  and (_34943_, _34942_, _34939_);
  nor (_34944_, _34943_, _34333_);
  nand (_34945_, _34921_, _34333_);
  nand (_34946_, _34945_, _07925_);
  or (_34948_, _34946_, _34944_);
  and (_34949_, _06065_, _05516_);
  or (_34950_, _34909_, _07925_);
  or (_34951_, _34950_, _34949_);
  and (_34952_, _34951_, _34948_);
  or (_34953_, _34952_, _03737_);
  and (_34954_, _06641_, _05516_);
  or (_34955_, _34909_, _03738_);
  or (_34956_, _34955_, _34954_);
  and (_34957_, _34956_, _03820_);
  and (_34959_, _34957_, _34953_);
  nor (_34960_, _13387_, _11630_);
  or (_34961_, _34960_, _34909_);
  and (_34962_, _34961_, _03455_);
  or (_34963_, _34962_, _03903_);
  or (_34964_, _34963_, _34959_);
  and (_34965_, _13394_, _05516_);
  or (_34966_, _34965_, _34909_);
  or (_34967_, _34966_, _04778_);
  and (_34968_, _34967_, _34964_);
  or (_34970_, _34968_, _03401_);
  or (_34971_, _34921_, _11641_);
  and (_34972_, _34971_, _34970_);
  or (_34973_, _34972_, _03897_);
  and (_34974_, _13402_, _05516_);
  or (_34975_, _34974_, _34909_);
  or (_34976_, _34975_, _04790_);
  and (_34977_, _34976_, _04792_);
  and (_34978_, _34977_, _34973_);
  and (_34979_, _08736_, _05516_);
  or (_34981_, _34979_, _34909_);
  and (_34982_, _34981_, _04018_);
  or (_34983_, _34982_, _34978_);
  and (_34984_, _34983_, _03909_);
  or (_34985_, _34909_, _08322_);
  and (_34986_, _34966_, _03908_);
  and (_34987_, _34986_, _34985_);
  or (_34988_, _34987_, _34984_);
  and (_34989_, _34988_, _10076_);
  nor (_34990_, _34915_, _04785_);
  and (_34992_, _34990_, _34985_);
  and (_34993_, _34921_, _03388_);
  or (_34994_, _34993_, _03914_);
  or (_34995_, _34994_, _34992_);
  or (_34996_, _34995_, _34989_);
  nor (_34997_, _13401_, _11630_);
  or (_34998_, _34909_, _06567_);
  or (_34999_, _34998_, _34997_);
  and (_35000_, _34999_, _34996_);
  or (_35001_, _35000_, _04011_);
  nor (_35003_, _08735_, _11630_);
  or (_35004_, _35003_, _34909_);
  or (_35005_, _35004_, _06572_);
  and (_35006_, _35005_, _10704_);
  and (_35007_, _35006_, _35001_);
  nor (_35008_, _11601_, _11597_);
  or (_35009_, _35008_, _11602_);
  and (_35010_, _35009_, _04034_);
  or (_35011_, _35010_, _03383_);
  or (_35012_, _35011_, _35007_);
  or (_35014_, _34921_, _03384_);
  and (_35015_, _35014_, _03778_);
  and (_35016_, _35015_, _35012_);
  and (_35017_, _35009_, _03777_);
  or (_35018_, _35017_, _03773_);
  or (_35019_, _35018_, _35016_);
  or (_35020_, _34911_, _03774_);
  and (_35021_, _35020_, _04819_);
  and (_35022_, _35021_, _35019_);
  and (_35023_, _34921_, _05223_);
  or (_35025_, _35023_, _03772_);
  or (_35026_, _35025_, _35022_);
  nor (_35027_, _13460_, _11630_);
  or (_35028_, _34909_, _04060_);
  or (_35029_, _35028_, _35027_);
  and (_35030_, _35029_, _43152_);
  and (_35031_, _35030_, _35026_);
  or (_35032_, _35031_, _34908_);
  and (_43570_, _35032_, _41894_);
  not (_35033_, \oc8051_golden_model_1.PSW [0]);
  nor (_35035_, _43152_, _35033_);
  and (_35036_, _03767_, _03412_);
  nor (_35037_, _07134_, _07133_);
  nor (_35038_, _35037_, _07036_);
  and (_35039_, _35037_, _07036_);
  nor (_35040_, _35039_, _35038_);
  nor (_35041_, _07055_, _07053_);
  nor (_35042_, _35041_, _15483_);
  and (_35043_, _35041_, _15483_);
  nor (_35044_, _35043_, _35042_);
  and (_35046_, _35044_, _35040_);
  nor (_35047_, _35044_, _35040_);
  nor (_35048_, _35047_, _35046_);
  or (_35049_, _35048_, _06554_);
  nand (_35050_, _35048_, _06554_);
  and (_35051_, _35050_, _35049_);
  and (_35052_, _35051_, _04197_);
  or (_35053_, _35051_, _04819_);
  nor (_35054_, _15000_, _08636_);
  not (_35055_, _15000_);
  nor (_35057_, _15451_, _35055_);
  nor (_35058_, _35057_, _35054_);
  nor (_35059_, _35058_, _15507_);
  and (_35060_, _35058_, _15507_);
  nor (_35061_, _35060_, _35059_);
  nor (_35062_, _35061_, _16075_);
  and (_35063_, _35061_, _16075_);
  or (_35064_, _35063_, _35062_);
  and (_35065_, _35064_, _16409_);
  nor (_35066_, _35064_, _16409_);
  or (_35068_, _35066_, _35065_);
  nor (_35069_, _35068_, _16758_);
  and (_35070_, _35068_, _16758_);
  or (_35071_, _35070_, _35069_);
  nor (_35072_, _35071_, _17089_);
  and (_35073_, _35071_, _17089_);
  or (_35074_, _35073_, _35072_);
  or (_35075_, _35074_, _08653_);
  nand (_35076_, _35074_, _08653_);
  and (_35077_, _35076_, _35075_);
  or (_35079_, _35077_, _04023_);
  and (_35080_, _35079_, _08659_);
  and (_35081_, _10065_, _10064_);
  nor (_35082_, _15009_, _08020_);
  and (_35083_, _15009_, _08020_);
  nor (_35084_, _35083_, _35082_);
  and (_35085_, _35084_, _08016_);
  nor (_35086_, _35084_, _08016_);
  or (_35087_, _35086_, _35085_);
  and (_35088_, _35087_, _08014_);
  nor (_35090_, _35087_, _08014_);
  or (_35091_, _35090_, _35088_);
  not (_35092_, _08007_);
  nor (_35093_, _08011_, _08004_);
  and (_35094_, _08011_, _08004_);
  nor (_35095_, _35094_, _35093_);
  nor (_35096_, _35095_, _35092_);
  and (_35097_, _35095_, _35092_);
  nor (_35098_, _35097_, _35096_);
  not (_35099_, _35098_);
  nor (_35101_, _35099_, _35091_);
  and (_35102_, _35099_, _35091_);
  nor (_35103_, _35102_, _35101_);
  nand (_35104_, _35103_, _08000_);
  or (_35105_, _35103_, _08000_);
  and (_35106_, _35105_, _35104_);
  and (_35107_, _35106_, _16374_);
  and (_35108_, _14996_, _08713_);
  nor (_35109_, _35108_, _15602_);
  and (_35110_, _35109_, _08704_);
  nor (_35112_, _35109_, _08704_);
  nor (_35113_, _35112_, _35110_);
  not (_35114_, _08697_);
  and (_35115_, _35114_, _08526_);
  nor (_35116_, _35114_, _08526_);
  nor (_35117_, _35116_, _35115_);
  nor (_35118_, _15841_, _08709_);
  and (_35119_, _15841_, _08709_);
  nor (_35120_, _35119_, _35118_);
  nor (_35121_, _35120_, _08700_);
  and (_35123_, _35120_, _08700_);
  nor (_35124_, _35123_, _35121_);
  and (_35125_, _35124_, _35117_);
  nor (_35126_, _35124_, _35117_);
  nor (_35127_, _35126_, _35125_);
  and (_35128_, _35127_, _35113_);
  nor (_35129_, _35127_, _35113_);
  or (_35130_, _35129_, _08520_);
  or (_35131_, _35130_, _35128_);
  and (_35132_, _04253_, _03757_);
  and (_35134_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_35135_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_35136_, _35135_, _35134_);
  and (_35137_, _35136_, _15276_);
  nor (_35138_, _35136_, _15276_);
  nor (_35139_, _35138_, _35137_);
  nor (_35140_, _15882_, _07090_);
  and (_35141_, _15882_, _07090_);
  nor (_35142_, _35141_, _35140_);
  and (_35143_, _35142_, _35139_);
  nor (_35145_, _35142_, _35139_);
  nor (_35146_, _35145_, _35143_);
  nor (_35147_, _35146_, _16541_);
  and (_35148_, _35146_, _16541_);
  nor (_35149_, _35148_, _35147_);
  nor (_35150_, _16885_, _08204_);
  and (_35151_, _16885_, _08204_);
  nor (_35152_, _35151_, _35150_);
  not (_35153_, _35152_);
  nor (_35154_, _35153_, _35149_);
  and (_35156_, _35153_, _35149_);
  or (_35157_, _35156_, _35154_);
  or (_35158_, _35157_, _11751_);
  or (_35159_, _06966_, _06825_);
  nand (_35160_, _35159_, _12240_);
  or (_35161_, _35159_, _12240_);
  nand (_35162_, _35161_, _35160_);
  nor (_35163_, _06970_, _06919_);
  nand (_35164_, _35163_, _06641_);
  or (_35165_, _35163_, _06641_);
  and (_35167_, _35165_, _35164_);
  nand (_35168_, _35167_, _35162_);
  or (_35169_, _35167_, _35162_);
  nand (_35170_, _35169_, _35168_);
  nor (_35171_, _35170_, _06248_);
  and (_35172_, _35170_, _06248_);
  or (_35173_, _35172_, _35171_);
  or (_35174_, _35173_, _08160_);
  and (_35175_, _04266_, _03436_);
  nor (_35176_, _06946_, _06126_);
  and (_35178_, _35176_, _12254_);
  nor (_35179_, _35176_, _12254_);
  nor (_35180_, _35179_, _35178_);
  nor (_35181_, _06948_, _06124_);
  nor (_35182_, _35181_, _06954_);
  and (_35183_, _35181_, _06954_);
  nor (_35184_, _35183_, _35182_);
  and (_35185_, _35184_, _35180_);
  nor (_35186_, _35184_, _35180_);
  or (_35187_, _35186_, _35185_);
  or (_35189_, _35187_, _10400_);
  and (_35190_, _26138_, _03770_);
  nand (_35191_, _35190_, _35033_);
  or (_35192_, _35190_, _35051_);
  and (_35193_, _35192_, _35191_);
  or (_35194_, _35193_, _08169_);
  and (_35195_, _35194_, _35189_);
  or (_35196_, _35195_, _08159_);
  and (_35197_, _35196_, _35175_);
  and (_35198_, _35197_, _35174_);
  and (_35200_, _35051_, _04267_);
  or (_35201_, _35200_, _04716_);
  or (_35202_, _35201_, _35198_);
  and (_35203_, _35161_, _35160_);
  nor (_35204_, _35041_, \oc8051_golden_model_1.ACC [6]);
  and (_35205_, _35041_, \oc8051_golden_model_1.ACC [6]);
  nor (_35206_, _35205_, _35204_);
  nor (_35207_, _35206_, \oc8051_golden_model_1.ACC [7]);
  and (_35208_, _35206_, \oc8051_golden_model_1.ACC [7]);
  nor (_35209_, _35208_, _35207_);
  nor (_35211_, _35209_, _35203_);
  and (_35212_, _35209_, _35203_);
  or (_35213_, _35212_, _35211_);
  or (_35214_, _35213_, _04717_);
  and (_35215_, _35214_, _04722_);
  and (_35216_, _35215_, _35202_);
  nor (_35217_, _16170_, _15876_);
  and (_35218_, _16170_, _15876_);
  nor (_35219_, _35218_, _35217_);
  and (_35220_, _35219_, _16878_);
  nor (_35222_, _35219_, _16878_);
  nor (_35223_, _35222_, _35220_);
  not (_35224_, _15038_);
  nor (_35225_, _15270_, _35224_);
  and (_35226_, _15270_, _35224_);
  nor (_35227_, _35226_, _35225_);
  and (_35228_, _35227_, _15529_);
  nor (_35229_, _35227_, _15529_);
  nor (_35230_, _35229_, _35228_);
  nor (_35231_, _35230_, _16534_);
  and (_35233_, _35230_, _16534_);
  or (_35234_, _35233_, _35231_);
  and (_35235_, _35234_, _08181_);
  nor (_35236_, _35234_, _08181_);
  or (_35237_, _35236_, _35235_);
  nand (_35238_, _35237_, _35223_);
  or (_35239_, _35237_, _35223_);
  and (_35240_, _35239_, _35238_);
  and (_35241_, _35240_, _03850_);
  or (_35242_, _35241_, _08179_);
  or (_35244_, _35242_, _35216_);
  and (_35245_, _35244_, _35158_);
  or (_35246_, _35245_, _10411_);
  or (_35247_, _35051_, _11764_);
  and (_35248_, _35247_, _03764_);
  and (_35249_, _35248_, _35246_);
  and (_35250_, _15283_, _15044_);
  nor (_35251_, _15283_, _15044_);
  or (_35252_, _35251_, _35250_);
  nor (_35253_, _15887_, _15543_);
  and (_35255_, _15887_, _15543_);
  nor (_35256_, _35255_, _35253_);
  not (_35257_, _35256_);
  and (_35258_, _35257_, _35252_);
  nor (_35259_, _35257_, _35252_);
  nor (_35260_, _35259_, _35258_);
  not (_35261_, _16892_);
  nor (_35262_, _16545_, _16182_);
  and (_35263_, _16545_, _16182_);
  nor (_35264_, _35263_, _35262_);
  nor (_35266_, _35264_, _35261_);
  and (_35267_, _35264_, _35261_);
  nor (_35268_, _35267_, _35266_);
  nor (_35269_, _35268_, _35260_);
  and (_35270_, _35268_, _35260_);
  nor (_35271_, _35270_, _35269_);
  and (_35272_, _35271_, _08210_);
  nor (_35273_, _35271_, _08210_);
  or (_35274_, _35273_, _35272_);
  and (_35275_, _35274_, _03763_);
  or (_35277_, _35275_, _05045_);
  or (_35278_, _35277_, _35249_);
  or (_35279_, _35051_, _03431_);
  and (_35280_, _35279_, _35278_);
  or (_35281_, _35280_, _03848_);
  not (_35282_, _16895_);
  and (_35283_, _35282_, _08214_);
  nor (_35284_, _35282_, _08214_);
  nor (_35285_, _35284_, _35283_);
  and (_35286_, _15286_, _15049_);
  nor (_35288_, _15286_, _15049_);
  nor (_35289_, _35288_, _35286_);
  not (_35290_, _15892_);
  and (_35291_, _35290_, _15546_);
  nor (_35292_, _35290_, _15546_);
  nor (_35293_, _35292_, _35291_);
  nor (_35294_, _35293_, _35289_);
  and (_35295_, _35293_, _35289_);
  or (_35296_, _35295_, _35294_);
  not (_35297_, _16549_);
  and (_35299_, _35297_, _16186_);
  nor (_35300_, _35297_, _16186_);
  nor (_35301_, _35300_, _35299_);
  and (_35302_, _35301_, _35296_);
  nor (_35303_, _35301_, _35296_);
  nor (_35304_, _35303_, _35302_);
  or (_35305_, _35304_, _35285_);
  nand (_35306_, _35304_, _35285_);
  and (_35307_, _35306_, _35305_);
  or (_35308_, _35307_, _04733_);
  and (_35310_, _35308_, _08157_);
  and (_35311_, _35310_, _35281_);
  and (_35312_, _04760_, _03757_);
  and (_35313_, _35187_, _08212_);
  or (_35314_, _35313_, _35312_);
  or (_35315_, _35314_, _35311_);
  not (_35316_, _35312_);
  or (_35317_, _35173_, _35316_);
  and (_35318_, _35317_, _35315_);
  or (_35319_, _35318_, _35132_);
  not (_35321_, _35132_);
  or (_35322_, _35173_, _35321_);
  and (_35323_, _35322_, _03855_);
  and (_35324_, _35323_, _35319_);
  nor (_35325_, _12262_, _05764_);
  and (_35326_, _12262_, _05764_);
  nor (_35327_, _35326_, _35325_);
  nor (_35328_, _06152_, _05955_);
  nor (_35329_, _35328_, _05622_);
  and (_35330_, _35328_, _05622_);
  nor (_35332_, _35330_, _35329_);
  nor (_35333_, _35332_, _06073_);
  and (_35334_, _35332_, _06073_);
  nor (_35335_, _35334_, _35333_);
  not (_35336_, _35335_);
  nand (_35337_, _35336_, _35327_);
  or (_35338_, _35336_, _35327_);
  and (_35339_, _35338_, _03854_);
  and (_35340_, _35339_, _35337_);
  or (_35341_, _35340_, _10434_);
  or (_35343_, _35341_, _35324_);
  or (_35344_, _35051_, _10431_);
  and (_35345_, _35344_, _03760_);
  and (_35346_, _35345_, _35343_);
  not (_35347_, _15908_);
  and (_35348_, _35347_, _15563_);
  nor (_35349_, _35347_, _15563_);
  nor (_35350_, _35349_, _35348_);
  nor (_35351_, _16567_, _16204_);
  and (_35352_, _16567_, _16204_);
  nor (_35354_, _35352_, _35351_);
  nor (_35355_, _35354_, _35350_);
  and (_35356_, _35354_, _35350_);
  nor (_35357_, _35356_, _35355_);
  nor (_35358_, _15303_, _15003_);
  and (_35359_, _15303_, _15003_);
  nor (_35360_, _35359_, _35358_);
  nor (_35361_, _16914_, _08232_);
  and (_35362_, _16914_, _08232_);
  nor (_35363_, _35362_, _35361_);
  not (_35365_, _35363_);
  and (_35366_, _35365_, _35360_);
  nor (_35367_, _35365_, _35360_);
  nor (_35368_, _35367_, _35366_);
  and (_35369_, _35368_, _35357_);
  nor (_35370_, _35368_, _35357_);
  or (_35371_, _35370_, _35369_);
  nand (_35372_, _35371_, _03759_);
  not (_35373_, _03911_);
  and (_35374_, _10256_, _35373_);
  nand (_35376_, _35374_, _35372_);
  or (_35377_, _35376_, _35346_);
  nor (_35378_, _35374_, _35051_);
  nor (_35379_, _35378_, _03896_);
  and (_35380_, _35379_, _35377_);
  and (_35381_, _35051_, _03896_);
  and (_35382_, _03822_, _03751_);
  and (_35383_, _03825_, _03751_);
  nor (_35384_, _35383_, _35382_);
  and (_35385_, _03834_, _03751_);
  nor (_35387_, _03927_, _35385_);
  nand (_35388_, _35387_, _35384_);
  or (_35389_, _35388_, _35381_);
  or (_35390_, _35389_, _35380_);
  not (_35391_, _35388_);
  or (_35392_, _35391_, _35051_);
  nor (_35393_, _03925_, _03868_);
  and (_35394_, _35393_, _26577_);
  and (_35395_, _35394_, _35392_);
  and (_35396_, _35395_, _35390_);
  not (_35399_, _35394_);
  and (_35400_, _35399_, _35051_);
  or (_35401_, _35400_, _27224_);
  or (_35402_, _35401_, _35396_);
  or (_35403_, _35051_, _10486_);
  and (_35404_, _35403_, _03753_);
  and (_35405_, _35404_, _35402_);
  not (_35406_, _15568_);
  and (_35407_, _35406_, _15308_);
  nor (_35408_, _35406_, _15308_);
  nor (_35410_, _35408_, _35407_);
  and (_35411_, _35410_, _16519_);
  nor (_35412_, _35410_, _16519_);
  or (_35413_, _35412_, _35411_);
  nor (_35414_, _15858_, _35224_);
  and (_35415_, _15858_, _35224_);
  nor (_35416_, _35415_, _35414_);
  and (_35417_, _35416_, _16210_);
  nor (_35418_, _35416_, _16210_);
  nor (_35419_, _35418_, _35417_);
  nor (_35422_, _35419_, _35413_);
  and (_35423_, _35419_, _35413_);
  nor (_35424_, _35423_, _35422_);
  not (_35425_, _16920_);
  and (_35426_, _35425_, _08237_);
  nor (_35427_, _35425_, _08237_);
  nor (_35428_, _35427_, _35426_);
  nand (_35429_, _35428_, _35424_);
  or (_35430_, _35428_, _35424_);
  and (_35431_, _35430_, _03752_);
  nand (_35433_, _35431_, _35429_);
  and (_35434_, _03910_, _03821_);
  not (_35435_, _35434_);
  nor (_35436_, _03843_, _05049_);
  and (_35437_, _35436_, _35435_);
  nand (_35438_, _35437_, _35433_);
  or (_35439_, _35438_, _35405_);
  and (_35440_, _03895_, _03821_);
  nor (_35441_, _35437_, _35051_);
  nor (_35442_, _35441_, _35440_);
  and (_35445_, _35442_, _35439_);
  nand (_35446_, _35051_, _35440_);
  not (_35447_, _03824_);
  and (_35448_, _03838_, _35447_);
  nand (_35449_, _35448_, _35446_);
  or (_35450_, _35449_, _35445_);
  nor (_35451_, _35448_, _35051_);
  nor (_35452_, _35451_, _03826_);
  and (_35453_, _35452_, _35450_);
  nand (_35454_, _35051_, _03826_);
  nor (_35456_, _04939_, _03832_);
  and (_35457_, _35456_, _10090_);
  nand (_35458_, _35457_, _35454_);
  or (_35459_, _35458_, _35453_);
  or (_35460_, _35457_, _35051_);
  and (_35461_, _35460_, _07405_);
  and (_35462_, _35461_, _35459_);
  and (_35463_, _10531_, _09879_);
  nor (_35464_, _15314_, _15070_);
  and (_35465_, _15314_, _15070_);
  or (_35468_, _35465_, _35464_);
  not (_35469_, _35468_);
  nor (_35470_, _35469_, _15573_);
  and (_35471_, _35469_, _15573_);
  nor (_35472_, _35471_, _35470_);
  or (_35473_, _35472_, _15853_);
  nand (_35474_, _35472_, _15853_);
  and (_35475_, _35474_, _35473_);
  nor (_35476_, _35475_, _16215_);
  and (_35477_, _35475_, _16215_);
  or (_35479_, _35477_, _35476_);
  nor (_35480_, _35479_, _16575_);
  and (_35481_, _35479_, _16575_);
  or (_35482_, _35481_, _35480_);
  nor (_35483_, _35482_, _16925_);
  and (_35484_, _35482_, _16925_);
  or (_35485_, _35484_, _35483_);
  or (_35486_, _35485_, _08242_);
  nand (_35487_, _35485_, _08242_);
  and (_35488_, _35487_, _07399_);
  nand (_35490_, _35488_, _35486_);
  nand (_35491_, _35490_, _35463_);
  or (_35492_, _35491_, _35462_);
  or (_35493_, _35463_, _35051_);
  and (_35494_, _35493_, _08152_);
  and (_35495_, _35494_, _35492_);
  not (_35496_, _08149_);
  not (_35497_, _08147_);
  not (_35498_, _16234_);
  or (_35499_, _15322_, _15020_);
  nand (_35501_, _15322_, _15020_);
  and (_35502_, _35501_, _35499_);
  nor (_35503_, _35502_, _15591_);
  and (_35504_, _35502_, _15591_);
  nor (_35505_, _35504_, _35503_);
  and (_35506_, _35505_, _15926_);
  nor (_35507_, _35505_, _15926_);
  or (_35508_, _35507_, _35506_);
  and (_35509_, _35508_, _35498_);
  nor (_35510_, _35508_, _35498_);
  nor (_35512_, _35510_, _35509_);
  nor (_35513_, _35512_, _16593_);
  and (_35514_, _35512_, _16593_);
  nor (_35515_, _35514_, _35513_);
  nor (_35516_, _35515_, _16942_);
  and (_35517_, _35515_, _16942_);
  or (_35518_, _35517_, _35516_);
  or (_35519_, _35518_, _35497_);
  nand (_35520_, _35518_, _35497_);
  and (_35521_, _35520_, _35519_);
  or (_35523_, _35521_, _35496_);
  and (_35524_, _35523_, _15513_);
  or (_35525_, _35524_, _35495_);
  or (_35526_, _35521_, _08149_);
  nand (_35527_, _04330_, _03420_);
  and (_35528_, _35527_, _35526_);
  and (_35529_, _35528_, _35525_);
  not (_35530_, _16253_);
  nor (_35531_, _15253_, _15077_);
  and (_35532_, _15253_, _15077_);
  or (_35534_, _35532_, _35531_);
  and (_35535_, _35534_, _15609_);
  nor (_35536_, _35534_, _15609_);
  or (_35537_, _35536_, _35535_);
  and (_35538_, _35537_, _15850_);
  nor (_35539_, _35537_, _15850_);
  or (_35540_, _35539_, _35538_);
  and (_35541_, _35540_, _35530_);
  nor (_35542_, _35540_, _35530_);
  nor (_35543_, _35542_, _35541_);
  and (_35545_, _35543_, _16514_);
  nor (_35546_, _35543_, _16514_);
  nor (_35547_, _35546_, _35545_);
  nor (_35548_, _35547_, _16862_);
  and (_35549_, _35547_, _16862_);
  or (_35550_, _35549_, _35548_);
  or (_35551_, _35550_, _08316_);
  nand (_35552_, _35550_, _08316_);
  and (_35553_, _35552_, _35551_);
  and (_35554_, _35553_, _04330_);
  or (_35556_, _35554_, _04331_);
  or (_35557_, _35556_, _35529_);
  or (_35558_, _35553_, _04332_);
  and (_35559_, _35558_, _03888_);
  and (_35560_, _35559_, _35557_);
  nor (_35561_, _15332_, _15000_);
  and (_35562_, _15332_, _15000_);
  or (_35563_, _35562_, _35561_);
  and (_35564_, _35563_, _15624_);
  nor (_35565_, _35563_, _15624_);
  or (_35567_, _35565_, _35564_);
  nor (_35568_, _35567_, _15947_);
  and (_35569_, _35567_, _15947_);
  nor (_35570_, _35569_, _35568_);
  or (_35571_, _35570_, _16268_);
  nand (_35572_, _35570_, _16268_);
  and (_35573_, _35572_, _35571_);
  nor (_35574_, _35573_, _16616_);
  and (_35575_, _35573_, _16616_);
  or (_35576_, _35575_, _35574_);
  nor (_35578_, _35576_, _16958_);
  and (_35579_, _35576_, _16958_);
  nor (_35580_, _35579_, _35578_);
  or (_35581_, _35580_, _08390_);
  nand (_35582_, _35580_, _08390_);
  and (_35583_, _35582_, _35581_);
  and (_35584_, _35583_, _03883_);
  or (_35585_, _35584_, _08320_);
  or (_35586_, _35585_, _35560_);
  not (_35587_, _16285_);
  nand (_35589_, _15340_, _15085_);
  or (_35590_, _15340_, _15085_);
  and (_35591_, _35590_, _35589_);
  and (_35592_, _35591_, _15638_);
  nor (_35593_, _35591_, _15638_);
  or (_35594_, _35593_, _35592_);
  and (_35595_, _35594_, _15961_);
  nor (_35596_, _35594_, _15961_);
  or (_35597_, _35596_, _35595_);
  and (_35598_, _35597_, _35587_);
  nor (_35600_, _35597_, _35587_);
  nor (_35601_, _35600_, _35598_);
  or (_35602_, _35601_, _16633_);
  nand (_35603_, _35601_, _16633_);
  and (_35604_, _35603_, _35602_);
  nor (_35605_, _35604_, _16972_);
  and (_35606_, _35604_, _16972_);
  nor (_35607_, _35606_, _35605_);
  nor (_35608_, _35607_, _08458_);
  and (_35609_, _35607_, _08458_);
  or (_35611_, _35609_, _35608_);
  or (_35612_, _35611_, _08321_);
  and (_35613_, _35612_, _35586_);
  or (_35614_, _35613_, _03425_);
  nor (_35615_, _05434_, _03811_);
  nor (_35616_, _05427_, _05420_);
  nor (_35617_, _05417_, _05457_);
  nor (_35618_, _05449_, _05416_);
  nor (_35619_, _35618_, _35617_);
  and (_35620_, _35618_, _35617_);
  nor (_35622_, _35620_, _35619_);
  nor (_35623_, _35622_, _35616_);
  and (_35624_, _35622_, _35616_);
  nor (_35625_, _35624_, _35623_);
  not (_35626_, _35625_);
  nor (_35627_, _35626_, _35615_);
  and (_35628_, _35626_, _35615_);
  or (_35629_, _35628_, _35627_);
  or (_35630_, _35629_, _03426_);
  and (_35631_, _35630_, _03747_);
  and (_35633_, _35631_, _35614_);
  not (_35634_, _15969_);
  and (_35635_, _35634_, _15647_);
  nor (_35636_, _35634_, _15647_);
  nor (_35637_, _35636_, _35635_);
  nor (_35638_, _16642_, _16294_);
  and (_35639_, _16642_, _16294_);
  nor (_35640_, _35639_, _35638_);
  nor (_35641_, _35640_, _35637_);
  and (_35642_, _35640_, _35637_);
  nor (_35644_, _35642_, _35641_);
  and (_35645_, _15348_, _15093_);
  nor (_35646_, _15348_, _15093_);
  or (_35647_, _35646_, _35645_);
  and (_35648_, _16981_, _08467_);
  nor (_35649_, _16981_, _08467_);
  nor (_35650_, _35649_, _35648_);
  not (_35651_, _35650_);
  and (_35652_, _35651_, _35647_);
  nor (_35653_, _35651_, _35647_);
  or (_35655_, _35653_, _35652_);
  not (_35656_, _35655_);
  nand (_35657_, _35656_, _35644_);
  or (_35658_, _35656_, _35644_);
  and (_35659_, _35658_, _03746_);
  nand (_35660_, _35659_, _35657_);
  nand (_35661_, _35660_, _28767_);
  or (_35662_, _35661_, _35633_);
  or (_35663_, _35051_, _28767_);
  and (_35664_, _35663_, _07920_);
  and (_35666_, _35664_, _35662_);
  or (_35667_, _35307_, _07923_);
  and (_35668_, _35667_, _08474_);
  or (_35669_, _35668_, _35666_);
  or (_35670_, _35307_, _07924_);
  and (_35671_, _35670_, _03738_);
  and (_35672_, _35671_, _35669_);
  not (_35673_, _16987_);
  and (_35674_, _35673_, _08472_);
  nor (_35675_, _35673_, _08472_);
  nor (_35677_, _35675_, _35674_);
  not (_35678_, _16648_);
  and (_35679_, _35678_, _16299_);
  nor (_35680_, _35678_, _16299_);
  nor (_35681_, _35680_, _35679_);
  and (_35682_, _15353_, _15098_);
  nor (_35683_, _15353_, _15098_);
  nor (_35684_, _35683_, _35682_);
  not (_35685_, _35684_);
  not (_35686_, _15974_);
  and (_35688_, _35686_, _15652_);
  nor (_35689_, _35686_, _15652_);
  nor (_35690_, _35689_, _35688_);
  and (_35691_, _35690_, _35685_);
  nor (_35692_, _35690_, _35685_);
  nor (_35693_, _35692_, _35691_);
  nor (_35694_, _35693_, _35681_);
  and (_35695_, _35693_, _35681_);
  nor (_35696_, _35695_, _35694_);
  or (_35697_, _35696_, _35677_);
  nand (_35699_, _35696_, _35677_);
  and (_35700_, _35699_, _35697_);
  and (_35701_, _35700_, _03737_);
  or (_35702_, _35701_, _35672_);
  and (_35703_, _35702_, _03820_);
  not (_35704_, _16994_);
  not (_35705_, _16655_);
  and (_35706_, _35705_, _16307_);
  nor (_35707_, _35705_, _16307_);
  nor (_35708_, _35707_, _35706_);
  not (_35710_, _35708_);
  and (_35711_, _15360_, _15105_);
  nor (_35712_, _15360_, _15105_);
  nor (_35713_, _35712_, _35711_);
  and (_35714_, _35713_, _15659_);
  nor (_35715_, _35713_, _15659_);
  or (_35716_, _35715_, _35714_);
  nand (_35717_, _35716_, _15981_);
  or (_35718_, _35716_, _15981_);
  and (_35719_, _35718_, _35717_);
  nor (_35721_, _35719_, _35710_);
  and (_35722_, _35719_, _35710_);
  nor (_35723_, _35722_, _35721_);
  nor (_35724_, _35723_, _35704_);
  and (_35725_, _35723_, _35704_);
  or (_35726_, _35725_, _35724_);
  and (_35727_, _35726_, _08481_);
  nor (_35728_, _35726_, _08481_);
  or (_35729_, _35728_, _35727_);
  and (_35730_, _35729_, _03455_);
  or (_35732_, _35730_, _07010_);
  or (_35733_, _35732_, _35703_);
  and (_35734_, _07069_, _17000_);
  nor (_35735_, _07069_, _17000_);
  nor (_35736_, _35735_, _35734_);
  not (_35737_, _35736_);
  nor (_35738_, _07151_, _07103_);
  and (_35739_, _07151_, _07103_);
  nor (_35740_, _35739_, _35738_);
  not (_35741_, _35740_);
  and (_35743_, _35741_, _07204_);
  nor (_35744_, _35741_, _07204_);
  nor (_35745_, _35744_, _35743_);
  and (_35746_, _35745_, _35737_);
  nor (_35747_, _35745_, _35737_);
  nor (_35748_, _35747_, _35746_);
  nand (_35749_, _35748_, _08485_);
  or (_35750_, _35748_, _08485_);
  and (_35751_, _35750_, _35749_);
  nor (_35752_, _35751_, _07269_);
  and (_35754_, _35751_, _07269_);
  nor (_35755_, _35754_, _35752_);
  not (_35756_, _35755_);
  nand (_35757_, _35756_, _07364_);
  or (_35758_, _35756_, _07364_);
  and (_35759_, _35758_, _35757_);
  or (_35760_, _35759_, _07011_);
  and (_35761_, _35760_, _35733_);
  or (_35762_, _35761_, _03469_);
  or (_35763_, _35629_, _03479_);
  and (_35765_, _35763_, _27373_);
  and (_35766_, _35765_, _35762_);
  nand (_35767_, _35051_, _03816_);
  and (_35768_, _25974_, _06138_);
  nand (_35769_, _35768_, _35767_);
  or (_35770_, _35769_, _35766_);
  or (_35771_, _35768_, _35051_);
  and (_35772_, _35771_, _04778_);
  and (_35773_, _35772_, _35770_);
  nor (_35774_, _15371_, _15115_);
  and (_35776_, _15371_, _15115_);
  or (_35777_, _35776_, _35774_);
  nor (_35778_, _15992_, _15670_);
  and (_35779_, _15992_, _15670_);
  nor (_35780_, _35779_, _35778_);
  nor (_35781_, _35780_, _35777_);
  and (_35782_, _35780_, _35777_);
  or (_35783_, _35782_, _35781_);
  nor (_35784_, _16668_, _16319_);
  and (_35785_, _16668_, _16319_);
  nor (_35787_, _35785_, _35784_);
  and (_35788_, _35787_, _16836_);
  nor (_35789_, _35787_, _16836_);
  nor (_35790_, _35789_, _35788_);
  and (_35791_, _35790_, _35783_);
  nor (_35792_, _35790_, _35783_);
  or (_35793_, _35792_, _35791_);
  or (_35794_, _35793_, _08495_);
  nand (_35795_, _35793_, _08495_);
  and (_35796_, _35795_, _03903_);
  and (_35798_, _35796_, _35794_);
  or (_35799_, _35798_, _35773_);
  and (_35800_, _35799_, _08493_);
  nand (_35801_, _35629_, _08492_);
  nor (_35802_, _10620_, _10580_);
  and (_35803_, _35802_, _10583_);
  nand (_35804_, _35803_, _35801_);
  or (_35805_, _35804_, _35800_);
  or (_35806_, _35803_, _35051_);
  and (_35807_, _35806_, _15999_);
  and (_35809_, _35807_, _35805_);
  and (_35810_, _16846_, _08002_);
  nor (_35811_, _16846_, _08002_);
  nor (_35812_, _35811_, _35810_);
  and (_35813_, _15122_, _08021_);
  nor (_35814_, _35813_, _15584_);
  and (_35815_, _15825_, _08017_);
  nor (_35816_, _15825_, _08017_);
  nor (_35817_, _35816_, _35815_);
  nor (_35818_, _35817_, _35814_);
  and (_35820_, _35817_, _35814_);
  nor (_35821_, _35820_, _35818_);
  and (_35822_, _08012_, _08008_);
  nor (_35823_, _08012_, _08008_);
  nor (_35824_, _35823_, _35822_);
  nor (_35825_, _35824_, _35821_);
  and (_35826_, _35824_, _35821_);
  nor (_35827_, _35826_, _35825_);
  nor (_35828_, _35827_, _35812_);
  and (_35829_, _35827_, _35812_);
  or (_35831_, _35829_, _35828_);
  and (_35832_, _35831_, _16001_);
  or (_35833_, _35832_, _08519_);
  or (_35834_, _35833_, _35809_);
  and (_35835_, _35834_, _35131_);
  or (_35836_, _35835_, _04016_);
  not (_35837_, _10489_);
  and (_35838_, _35837_, _08752_);
  nor (_35839_, _35838_, _10490_);
  nor (_35840_, _10493_, _06557_);
  and (_35842_, _10493_, _06557_);
  nor (_35843_, _35842_, _35840_);
  nor (_35844_, _35843_, _35839_);
  and (_35845_, _35843_, _35839_);
  nor (_35846_, _35845_, _35844_);
  and (_35847_, _10491_, _08748_);
  nor (_35848_, _35847_, _10492_);
  nor (_35849_, _08736_, _08741_);
  and (_35850_, _08736_, _08741_);
  nor (_35851_, _35850_, _35849_);
  nor (_35853_, _35851_, _35848_);
  and (_35854_, _35851_, _35848_);
  nor (_35855_, _35854_, _35853_);
  nand (_35856_, _35855_, _35846_);
  or (_35857_, _35855_, _35846_);
  and (_35858_, _35857_, _35856_);
  or (_35859_, _35858_, _04017_);
  and (_35860_, _35859_, _08531_);
  and (_35861_, _35860_, _35836_);
  and (_35862_, _08776_, _08537_);
  nor (_35864_, _35862_, _10512_);
  and (_35865_, _08779_, _08783_);
  nor (_35866_, _35865_, _10511_);
  not (_35867_, _35866_);
  and (_35868_, _10509_, _08788_);
  nor (_35869_, _35868_, _10510_);
  not (_35870_, _35869_);
  and (_35871_, _10507_, _08792_);
  nor (_35872_, _35871_, _10508_);
  and (_35873_, _35872_, _35870_);
  nor (_35875_, _35872_, _35870_);
  nor (_35876_, _35875_, _35873_);
  nor (_35877_, _35876_, _35867_);
  and (_35878_, _35876_, _35867_);
  nor (_35879_, _35878_, _35877_);
  not (_35880_, _35879_);
  nor (_35881_, _35880_, _35864_);
  and (_35882_, _35880_, _35864_);
  or (_35883_, _35882_, _35881_);
  and (_35884_, _35883_, _08530_);
  or (_35886_, _35884_, _03897_);
  or (_35887_, _35886_, _35861_);
  not (_35888_, _16840_);
  not (_35889_, _16496_);
  and (_35890_, _35889_, _16153_);
  nor (_35891_, _35889_, _16153_);
  nor (_35892_, _35891_, _35890_);
  not (_35893_, _35892_);
  and (_35894_, _15244_, _15016_);
  nor (_35895_, _15244_, _15016_);
  nor (_35897_, _35895_, _35894_);
  and (_35898_, _15836_, _15699_);
  nor (_35899_, _15836_, _15699_);
  nor (_35900_, _35899_, _35898_);
  nor (_35901_, _35900_, _35897_);
  and (_35902_, _35900_, _35897_);
  nor (_35903_, _35902_, _35901_);
  nor (_35904_, _35903_, _35893_);
  and (_35905_, _35903_, _35893_);
  nor (_35906_, _35905_, _35904_);
  nor (_35908_, _35906_, _35888_);
  and (_35909_, _35906_, _35888_);
  or (_35910_, _35909_, _35908_);
  and (_35911_, _35910_, _08126_);
  nor (_35912_, _35910_, _08126_);
  or (_35913_, _35912_, _35911_);
  or (_35914_, _35913_, _04790_);
  and (_35915_, _35914_, _10639_);
  and (_35916_, _35915_, _35887_);
  nand (_35917_, _35051_, _04018_);
  nor (_35919_, _35917_, _05429_);
  or (_35920_, _35919_, _35916_);
  and (_35921_, _35920_, _10644_);
  not (_35922_, _29486_);
  and (_35923_, _35051_, _35922_);
  or (_35924_, _35923_, _04599_);
  or (_35925_, _35924_, _35921_);
  and (_35926_, _03767_, _03387_);
  not (_35927_, _04599_);
  or (_35928_, _08022_, _08019_);
  nand (_35930_, _08022_, _08019_);
  and (_35931_, _35930_, _35928_);
  and (_35932_, _15708_, _08013_);
  nor (_35933_, _15708_, _08013_);
  nor (_35934_, _35933_, _35932_);
  and (_35935_, _35934_, _35931_);
  nor (_35936_, _35934_, _35931_);
  nor (_35937_, _35936_, _35935_);
  nor (_35938_, _08010_, _08003_);
  and (_35939_, _08010_, _08003_);
  nor (_35941_, _35939_, _35938_);
  nor (_35942_, _35941_, _16490_);
  and (_35943_, _35941_, _16490_);
  nor (_35944_, _35943_, _35942_);
  and (_35945_, _35944_, _35937_);
  nor (_35946_, _35944_, _35937_);
  or (_35947_, _35946_, _35945_);
  and (_35948_, _35947_, _08001_);
  nor (_35949_, _35947_, _08001_);
  or (_35950_, _35949_, _35948_);
  nor (_35952_, _35950_, _35927_);
  nor (_35953_, _35952_, _35926_);
  and (_35954_, _35953_, _35925_);
  and (_35955_, _35950_, _35926_);
  or (_35956_, _35955_, _04406_);
  or (_35957_, _35956_, _35954_);
  nand (_35958_, _03825_, _03387_);
  and (_35959_, _35958_, _16019_);
  or (_35960_, _35950_, _04407_);
  and (_35961_, _35960_, _35959_);
  and (_35963_, _35961_, _35957_);
  or (_35964_, _35950_, _03308_);
  and (_35965_, _35964_, _16355_);
  or (_35966_, _35965_, _35963_);
  nor (_35967_, _35950_, _15715_);
  and (_35968_, _08547_, _03420_);
  nor (_35969_, _35968_, _35967_);
  and (_35970_, _35969_, _35966_);
  not (_35971_, _08707_);
  or (_35972_, _08714_, _08711_);
  nand (_35974_, _08714_, _08711_);
  and (_35975_, _35974_, _35972_);
  nand (_35976_, _35975_, _35971_);
  or (_35977_, _35975_, _35971_);
  and (_35978_, _35977_, _35976_);
  nor (_35979_, _35978_, _08705_);
  and (_35980_, _35978_, _08705_);
  or (_35981_, _35980_, _35979_);
  nor (_35982_, _08698_, _08702_);
  and (_35983_, _08698_, _08702_);
  nor (_35985_, _35983_, _35982_);
  and (_35986_, _08695_, _08525_);
  nor (_35987_, _35986_, _11998_);
  nor (_35988_, _35987_, _35985_);
  and (_35989_, _35987_, _35985_);
  nor (_35990_, _35989_, _35988_);
  or (_35991_, _35990_, _35981_);
  nand (_35992_, _35990_, _35981_);
  and (_35993_, _35992_, _35991_);
  and (_35994_, _35993_, _35968_);
  or (_35996_, _35994_, _04413_);
  or (_35997_, _35996_, _35970_);
  not (_35998_, _04413_);
  or (_35999_, _35993_, _35998_);
  and (_36000_, _35999_, _04026_);
  and (_36001_, _36000_, _35997_);
  or (_36002_, _08753_, _08750_);
  nand (_36003_, _08753_, _08750_);
  and (_36004_, _36003_, _36002_);
  and (_36005_, _08745_, _08746_);
  nor (_36007_, _08745_, _08746_);
  nor (_36008_, _36007_, _36005_);
  and (_36009_, _36008_, _36004_);
  nor (_36010_, _36008_, _36004_);
  nor (_36011_, _36010_, _36009_);
  or (_36012_, _36011_, _08739_);
  nand (_36013_, _36011_, _08739_);
  and (_36014_, _36013_, _36012_);
  or (_36015_, _36014_, _08737_);
  nand (_36016_, _36014_, _08737_);
  and (_36018_, _36016_, _36015_);
  or (_36019_, _36018_, _08734_);
  nand (_36020_, _36018_, _08734_);
  and (_36021_, _36020_, _36019_);
  or (_36022_, _36021_, _12005_);
  nand (_36023_, _36021_, _12005_);
  and (_36024_, _36023_, _04025_);
  and (_36025_, _36024_, _36022_);
  or (_36026_, _36025_, _08553_);
  or (_36027_, _36026_, _36001_);
  or (_36029_, _08793_, _08790_);
  nand (_36030_, _08793_, _08790_);
  and (_36031_, _36030_, _36029_);
  not (_36032_, _08784_);
  and (_36033_, _36032_, _08786_);
  nor (_36034_, _36032_, _08786_);
  nor (_36035_, _36034_, _36033_);
  and (_36036_, _36035_, _36031_);
  nor (_36037_, _36035_, _36031_);
  nor (_36038_, _36037_, _36036_);
  nor (_36040_, _08774_, _08536_);
  and (_36041_, _08774_, _08536_);
  nor (_36042_, _36041_, _36040_);
  nor (_36043_, _08777_, _08781_);
  and (_36044_, _08777_, _08781_);
  nor (_36045_, _36044_, _36043_);
  and (_36046_, _36045_, _36042_);
  nor (_36047_, _36045_, _36042_);
  nor (_36048_, _36047_, _36046_);
  and (_36049_, _36048_, _36038_);
  nor (_36051_, _36048_, _36038_);
  or (_36052_, _36051_, _36049_);
  or (_36053_, _36052_, _08557_);
  and (_36054_, _36053_, _03909_);
  and (_36055_, _36054_, _36027_);
  and (_36056_, _10076_, _10075_);
  nor (_36057_, _15728_, _15152_);
  and (_36058_, _15728_, _15152_);
  nor (_36059_, _36058_, _36057_);
  nor (_36060_, _16837_, _16375_);
  and (_36062_, _16837_, _16375_);
  nor (_36063_, _36062_, _36060_);
  and (_36064_, _36063_, _36059_);
  nor (_36065_, _36063_, _36059_);
  nor (_36066_, _36065_, _36064_);
  nor (_36067_, _16041_, _15414_);
  and (_36068_, _16041_, _15414_);
  nor (_36069_, _36068_, _36067_);
  nor (_36070_, _16721_, _08561_);
  and (_36071_, _16721_, _08561_);
  nor (_36073_, _36071_, _36070_);
  and (_36074_, _36073_, _36069_);
  nor (_36075_, _36073_, _36069_);
  nor (_36076_, _36075_, _36074_);
  not (_36077_, _36076_);
  nand (_36078_, _36077_, _36066_);
  or (_36079_, _36077_, _36066_);
  and (_36080_, _36079_, _03908_);
  nand (_36081_, _36080_, _36078_);
  nand (_36082_, _36081_, _36056_);
  or (_36084_, _36082_, _36055_);
  or (_36085_, _35051_, _36056_);
  and (_36086_, _36085_, _10071_);
  and (_36087_, _36086_, _36084_);
  or (_36088_, _36087_, _35107_);
  and (_36089_, _36088_, _08569_);
  and (_36090_, _35106_, _08568_);
  or (_36091_, _36090_, _08573_);
  or (_36092_, _36091_, _36089_);
  not (_36093_, _08524_);
  nor (_36095_, _14995_, _08712_);
  and (_36096_, _14995_, _08712_);
  nor (_36097_, _36096_, _36095_);
  and (_36098_, _36097_, _08708_);
  nor (_36099_, _36097_, _08708_);
  or (_36100_, _36099_, _36098_);
  nand (_36101_, _36100_, _08706_);
  or (_36102_, _36100_, _08706_);
  and (_36103_, _36102_, _36101_);
  nor (_36104_, _08703_, _08696_);
  and (_36106_, _08703_, _08696_);
  nor (_36107_, _36106_, _36104_);
  and (_36108_, _36107_, _08699_);
  nor (_36109_, _36107_, _08699_);
  nor (_36110_, _36109_, _36108_);
  and (_36111_, _36110_, _36103_);
  nor (_36112_, _36110_, _36103_);
  or (_36113_, _36112_, _36111_);
  and (_36114_, _36113_, _36093_);
  or (_36115_, _36113_, _36093_);
  nand (_36117_, _36115_, _08573_);
  or (_36118_, _36117_, _36114_);
  and (_36119_, _36118_, _04014_);
  and (_36120_, _36119_, _36092_);
  nor (_36121_, _10488_, _08751_);
  and (_36122_, _10488_, _08751_);
  nor (_36123_, _36122_, _36121_);
  not (_36124_, _36123_);
  and (_36125_, _08743_, _08747_);
  nor (_36126_, _08743_, _08747_);
  nor (_36128_, _36126_, _36125_);
  nor (_36129_, _36128_, _36124_);
  and (_36130_, _36128_, _36124_);
  nor (_36131_, _36130_, _36129_);
  and (_36132_, _36131_, _08740_);
  nor (_36133_, _36131_, _08740_);
  or (_36134_, _36133_, _36132_);
  and (_36135_, _36134_, _08738_);
  nor (_36136_, _36134_, _08738_);
  or (_36137_, _36136_, _36135_);
  and (_36139_, _36137_, _08735_);
  nor (_36140_, _36137_, _08735_);
  or (_36141_, _36140_, _36139_);
  and (_36142_, _36141_, _06556_);
  nor (_36143_, _36141_, _06556_);
  or (_36144_, _36143_, _36142_);
  and (_36145_, _36144_, _04013_);
  or (_36146_, _36145_, _08580_);
  or (_36147_, _36146_, _36120_);
  nor (_36148_, _10506_, _08791_);
  and (_36150_, _10506_, _08791_);
  nor (_36151_, _36150_, _36148_);
  not (_36152_, _08785_);
  and (_36153_, _36152_, _08787_);
  nor (_36154_, _36152_, _08787_);
  nor (_36155_, _36154_, _36153_);
  and (_36156_, _36155_, _36151_);
  nor (_36157_, _36155_, _36151_);
  nor (_36158_, _36157_, _36156_);
  not (_36159_, _08782_);
  nor (_36161_, _08778_, _08775_);
  and (_36162_, _08778_, _08775_);
  nor (_36163_, _36162_, _36161_);
  nor (_36164_, _36163_, _36159_);
  and (_36165_, _36163_, _36159_);
  nor (_36166_, _36165_, _36164_);
  and (_36167_, _36166_, _36158_);
  nor (_36168_, _36166_, _36158_);
  or (_36169_, _36168_, _36167_);
  and (_36170_, _36169_, _08535_);
  nor (_36172_, _36169_, _08535_);
  or (_36173_, _36172_, _36170_);
  or (_36174_, _36173_, _08583_);
  and (_36175_, _36174_, _06567_);
  and (_36176_, _36175_, _36147_);
  nor (_36177_, _15436_, _15005_);
  and (_36178_, _15436_, _15005_);
  or (_36179_, _36178_, _36177_);
  nor (_36180_, _15832_, _15749_);
  and (_36181_, _15832_, _15749_);
  nor (_36183_, _36181_, _36180_);
  nor (_36184_, _36183_, _36179_);
  and (_36185_, _36183_, _36179_);
  nor (_36186_, _36185_, _36184_);
  and (_36187_, _36186_, _16396_);
  nor (_36188_, _36186_, _16396_);
  or (_36189_, _36188_, _36187_);
  and (_36190_, _36189_, _16745_);
  nor (_36191_, _36189_, _16745_);
  or (_36192_, _36191_, _36190_);
  and (_36194_, _36192_, _17076_);
  nor (_36195_, _36192_, _17076_);
  or (_36196_, _36195_, _36194_);
  and (_36197_, _36196_, _08592_);
  nor (_36198_, _36196_, _08592_);
  or (_36199_, _36198_, _36197_);
  and (_36200_, _36199_, _03914_);
  or (_36201_, _36200_, _36176_);
  and (_36202_, _36201_, _35081_);
  not (_36203_, _35081_);
  nand (_36205_, _35051_, _36203_);
  nand (_36206_, _36205_, _08119_);
  or (_36207_, _36206_, _36202_);
  not (_36208_, _16486_);
  not (_36209_, _16065_);
  nor (_36210_, _15441_, _15020_);
  and (_36211_, _15441_, _15020_);
  or (_36212_, _36211_, _36210_);
  nor (_36213_, _36212_, _15754_);
  and (_36214_, _36212_, _15754_);
  nor (_36216_, _36214_, _36213_);
  and (_36217_, _36216_, _36209_);
  nor (_36218_, _36216_, _36209_);
  nor (_36219_, _36218_, _36217_);
  nor (_36220_, _36219_, _16401_);
  and (_36221_, _36219_, _16401_);
  or (_36222_, _36221_, _36220_);
  nor (_36223_, _36222_, _36208_);
  and (_36224_, _36222_, _36208_);
  nor (_36225_, _36224_, _36223_);
  nor (_36227_, _36225_, _17081_);
  and (_36228_, _36225_, _17081_);
  or (_36229_, _36228_, _36227_);
  nand (_36230_, _36229_, _08111_);
  or (_36231_, _36229_, _08111_);
  and (_36232_, _36231_, _36230_);
  or (_36233_, _36232_, _08119_);
  and (_36234_, _36233_, _08599_);
  and (_36235_, _36234_, _36207_);
  not (_36236_, _16070_);
  nor (_36238_, _15446_, _15077_);
  and (_36239_, _15446_, _15077_);
  or (_36240_, _36239_, _36238_);
  nor (_36241_, _36240_, _15759_);
  and (_36242_, _36240_, _15759_);
  nor (_36243_, _36242_, _36241_);
  and (_36244_, _36243_, _36236_);
  nor (_36245_, _36243_, _36236_);
  nor (_36246_, _36245_, _36244_);
  and (_36247_, _36246_, _16147_);
  nor (_36249_, _36246_, _16147_);
  nor (_36250_, _36249_, _36247_);
  nor (_36251_, _36250_, _16752_);
  and (_36252_, _36250_, _16752_);
  or (_36253_, _36252_, _36251_);
  nor (_36254_, _36253_, _16828_);
  and (_36255_, _36253_, _16828_);
  or (_36256_, _36255_, _36254_);
  nor (_36257_, _36256_, _08623_);
  and (_36258_, _36256_, _08623_);
  or (_36260_, _36258_, _36257_);
  and (_36261_, _36260_, _08597_);
  or (_36262_, _36261_, _04022_);
  or (_36263_, _36262_, _36235_);
  and (_36264_, _36263_, _35080_);
  nor (_36265_, _15237_, _15085_);
  and (_36266_, _15237_, _15085_);
  or (_36267_, _36266_, _36265_);
  nor (_36268_, _36267_, _15765_);
  and (_36269_, _36267_, _15765_);
  nor (_36271_, _36269_, _36268_);
  and (_36272_, _36271_, _16080_);
  nor (_36273_, _36271_, _16080_);
  nor (_36274_, _36273_, _36272_);
  nor (_36275_, _36274_, _16415_);
  and (_36276_, _36274_, _16415_);
  or (_36277_, _36276_, _36275_);
  nor (_36278_, _36277_, _16763_);
  and (_36279_, _36277_, _16763_);
  or (_36280_, _36279_, _36278_);
  and (_36282_, _36280_, _17094_);
  nor (_36283_, _36280_, _17094_);
  nor (_36284_, _36283_, _36282_);
  nand (_36285_, _36284_, _08683_);
  or (_36286_, _36284_, _08683_);
  and (_36287_, _36286_, _36285_);
  and (_36288_, _36287_, _08627_);
  or (_36289_, _36288_, _08657_);
  or (_36290_, _36289_, _36264_);
  and (_36291_, _29228_, _10704_);
  nor (_36293_, _15247_, _15246_);
  nor (_36294_, _15535_, \oc8051_golden_model_1.ACC [3]);
  and (_36295_, _15535_, \oc8051_golden_model_1.ACC [3]);
  nor (_36296_, _36295_, _36294_);
  and (_36297_, _36296_, _35206_);
  nor (_36298_, _36296_, _35206_);
  nor (_36299_, _36298_, _36297_);
  nor (_36300_, _36299_, _36293_);
  and (_36301_, _36299_, _36293_);
  nor (_36302_, _36301_, _36300_);
  nand (_36304_, _36302_, _08657_);
  and (_36305_, _36304_, _36291_);
  and (_36306_, _36305_, _36290_);
  not (_36307_, _36291_);
  nand (_36308_, _36307_, _35051_);
  nand (_36309_, _36308_, _11984_);
  or (_36310_, _36309_, _36306_);
  nor (_36311_, _15462_, _15122_);
  nor (_36312_, _36311_, _35813_);
  nor (_36313_, _36312_, _15773_);
  and (_36315_, _36312_, _15773_);
  or (_36316_, _36315_, _36313_);
  nor (_36317_, _36316_, _15828_);
  and (_36318_, _36316_, _15828_);
  nor (_36319_, _36318_, _36317_);
  and (_36320_, _36319_, _16423_);
  nor (_36321_, _36319_, _16423_);
  nor (_36322_, _36321_, _36320_);
  and (_36323_, _36322_, _16483_);
  nor (_36324_, _36322_, _16483_);
  or (_36326_, _36324_, _36323_);
  nor (_36327_, _36326_, _17103_);
  and (_36328_, _36326_, _17103_);
  or (_36329_, _36328_, _36327_);
  or (_36330_, _36329_, _08037_);
  nand (_36331_, _36329_, _08037_);
  and (_36332_, _36331_, _36330_);
  or (_36333_, _36332_, _11984_);
  and (_36334_, _36333_, _11987_);
  and (_36335_, _36334_, _36310_);
  and (_36337_, _36332_, _04456_);
  or (_36338_, _36337_, _08691_);
  or (_36339_, _36338_, _36335_);
  nor (_36340_, _14995_, _08713_);
  and (_36341_, _14995_, _08713_);
  nor (_36342_, _36341_, _36340_);
  and (_36343_, _36342_, _15778_);
  nor (_36344_, _36342_, _15778_);
  nor (_36345_, _36344_, _36343_);
  and (_36346_, _36345_, _16092_);
  nor (_36348_, _36345_, _16092_);
  nor (_36349_, _36348_, _36346_);
  and (_36350_, _36349_, _16429_);
  nor (_36351_, _36349_, _16429_);
  nor (_36352_, _36351_, _36350_);
  nor (_36353_, _36352_, _16774_);
  and (_36354_, _36352_, _16774_);
  or (_36355_, _36354_, _36353_);
  and (_36356_, _36355_, _17109_);
  nor (_36357_, _36355_, _17109_);
  nor (_36359_, _36357_, _36356_);
  or (_36360_, _36359_, _08729_);
  nand (_36361_, _36359_, _08729_);
  and (_36362_, _36361_, _36360_);
  or (_36363_, _36362_, _10058_);
  and (_36364_, _36363_, _10056_);
  and (_36365_, _36364_, _36339_);
  nor (_36366_, _15469_, _35837_);
  nor (_36367_, _36366_, _35838_);
  nor (_36368_, _36367_, _15783_);
  and (_36370_, _36367_, _15783_);
  or (_36371_, _36370_, _36368_);
  nor (_36372_, _36371_, _16099_);
  and (_36373_, _36371_, _16099_);
  nor (_36374_, _36373_, _36372_);
  nor (_36375_, _36374_, _16434_);
  and (_36376_, _36374_, _16434_);
  or (_36377_, _36376_, _36375_);
  nor (_36378_, _36377_, _16781_);
  and (_36379_, _36377_, _16781_);
  nor (_36381_, _36379_, _36378_);
  and (_36382_, _36381_, _17114_);
  nor (_36383_, _36381_, _17114_);
  nor (_36384_, _36383_, _36382_);
  and (_36385_, _36384_, _08768_);
  nor (_36386_, _36384_, _08768_);
  or (_36387_, _36386_, _36385_);
  and (_36388_, _36387_, _03779_);
  and (_36389_, _29249_, _08773_);
  nor (_36390_, _04200_, _03777_);
  and (_36392_, _36390_, _36389_);
  not (_36393_, _10506_);
  and (_36394_, _36393_, _08792_);
  nor (_36395_, _36393_, _08792_);
  nor (_36396_, _36395_, _36394_);
  and (_36397_, _36396_, _15788_);
  nor (_36398_, _36396_, _15788_);
  nor (_36399_, _36398_, _36397_);
  and (_36400_, _36399_, _16105_);
  nor (_36401_, _36399_, _16105_);
  nor (_36403_, _36401_, _36400_);
  and (_36404_, _36403_, _16440_);
  nor (_36405_, _36403_, _16440_);
  nor (_36406_, _36405_, _36404_);
  and (_36407_, _36406_, _16786_);
  nor (_36408_, _36406_, _16786_);
  nor (_36409_, _36408_, _36407_);
  and (_36410_, _36409_, _17120_);
  nor (_36411_, _36409_, _17120_);
  nor (_36412_, _36411_, _36410_);
  or (_36414_, _36412_, _08808_);
  nand (_36415_, _36412_, _08808_);
  and (_36416_, _36415_, _08733_);
  nand (_36417_, _36416_, _36414_);
  nand (_36418_, _36417_, _36392_);
  or (_36419_, _36418_, _36388_);
  or (_36420_, _36419_, _36365_);
  and (_36421_, _04196_, _03420_);
  nor (_36422_, _36392_, _35051_);
  nor (_36423_, _36422_, _36421_);
  and (_36425_, _36423_, _36420_);
  or (_36426_, _05053_, _04812_);
  nor (_36427_, _06583_, _36426_);
  nand (_36428_, _35051_, _36421_);
  nand (_36429_, _36428_, _36427_);
  or (_36430_, _36429_, _36425_);
  or (_36431_, _36427_, _35051_);
  and (_36432_, _36431_, _03774_);
  and (_36433_, _36432_, _36430_);
  and (_36434_, _35240_, _03773_);
  or (_36436_, _36434_, _08815_);
  or (_36437_, _36436_, _36433_);
  not (_36438_, _08821_);
  and (_36439_, _15535_, _36438_);
  and (_36440_, _36439_, \oc8051_golden_model_1.ACC [3]);
  nor (_36441_, _36439_, \oc8051_golden_model_1.ACC [3]);
  nor (_36442_, _36441_, _36440_);
  and (_36443_, _36442_, _16453_);
  nor (_36444_, _36442_, _16453_);
  nor (_36445_, _36444_, _36443_);
  and (_36447_, _16797_, _07036_);
  nor (_36448_, _16797_, _07036_);
  nor (_36449_, _36448_, _36447_);
  nor (_36450_, _36449_, _36445_);
  and (_36451_, _36449_, _36445_);
  or (_36452_, _36451_, _36450_);
  nor (_36453_, _36452_, _08827_);
  and (_36454_, _36452_, _08827_);
  nor (_36455_, _36454_, _36453_);
  nand (_36456_, _36455_, _08815_);
  and (_36458_, _36456_, _12016_);
  and (_36459_, _36458_, _36437_);
  and (_36460_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_36461_, _36460_, _08200_);
  nand (_36462_, _36461_, _36299_);
  or (_36463_, _36461_, _36299_);
  and (_36464_, _36463_, _36462_);
  nand (_36465_, _36464_, _08820_);
  nand (_36466_, _36465_, _04819_);
  or (_36467_, _36466_, _36459_);
  and (_36469_, _36467_, _35053_);
  or (_36470_, _36469_, _03374_);
  nor (_36471_, _35371_, _03375_);
  nor (_36472_, _36471_, _04197_);
  and (_36473_, _36472_, _36470_);
  nor (_36474_, _36473_, _35052_);
  nor (_36475_, _36474_, _35036_);
  or (_36476_, _04629_, _04488_);
  and (_36477_, _35051_, _35036_);
  or (_36478_, _36477_, _36476_);
  or (_36480_, _36478_, _36475_);
  not (_36481_, _36476_);
  nor (_36482_, _35051_, _36481_);
  nor (_36483_, _36482_, _05018_);
  and (_36484_, _36483_, _36480_);
  and (_36485_, _35051_, _05018_);
  or (_36486_, _36485_, _26459_);
  or (_36487_, _36486_, _36484_);
  or (_36488_, _35051_, _05038_);
  and (_36489_, _36488_, _04060_);
  and (_36491_, _36489_, _36487_);
  not (_36492_, _16129_);
  nor (_36493_, _15493_, _15038_);
  and (_36494_, _15493_, _15038_);
  nor (_36495_, _36494_, _36493_);
  and (_36496_, _36495_, _15810_);
  nor (_36497_, _36495_, _15810_);
  nor (_36498_, _36497_, _36496_);
  nor (_36499_, _36498_, _36492_);
  and (_36500_, _36498_, _36492_);
  or (_36502_, _36500_, _36499_);
  and (_36503_, _36502_, _16466_);
  nor (_36504_, _36502_, _16466_);
  or (_36505_, _36504_, _36503_);
  and (_36506_, _36505_, _16811_);
  nor (_36507_, _36505_, _16811_);
  or (_36508_, _36507_, _36506_);
  and (_36509_, _36508_, _17143_);
  nor (_36510_, _36508_, _17143_);
  or (_36511_, _36510_, _36509_);
  and (_36513_, _36511_, _08840_);
  nor (_36514_, _36511_, _08840_);
  or (_36515_, _36514_, _36513_);
  and (_36516_, _36515_, _03772_);
  or (_36517_, _36516_, _08837_);
  or (_36518_, _36517_, _36491_);
  not (_36519_, _08845_);
  and (_36520_, _15535_, _36519_);
  and (_36521_, _36520_, \oc8051_golden_model_1.ACC [3]);
  nor (_36522_, _36520_, \oc8051_golden_model_1.ACC [3]);
  nor (_36524_, _36522_, _36521_);
  or (_36525_, _17148_, _16472_);
  nand (_36526_, _17148_, _16472_);
  and (_36527_, _36526_, _36525_);
  or (_36528_, _36527_, _36524_);
  nand (_36529_, _36527_, _36524_);
  and (_36530_, _36529_, _36528_);
  nor (_36531_, _16816_, _08852_);
  and (_36532_, _16816_, _08852_);
  nor (_36533_, _36532_, _36531_);
  nor (_36535_, _36533_, _36530_);
  nand (_36536_, _36533_, _36530_);
  nand (_36537_, _36536_, _08837_);
  or (_36538_, _36537_, _36535_);
  and (_36539_, _36538_, _36518_);
  or (_36540_, _36539_, _08844_);
  not (_36541_, _08844_);
  or (_36542_, _35051_, _36541_);
  and (_36543_, _36542_, _10969_);
  and (_36544_, _36543_, _36540_);
  nand (_36546_, _35051_, _03901_);
  nand (_36547_, _36546_, _28948_);
  or (_36548_, _36547_, _36544_);
  or (_36549_, _35051_, _28948_);
  and (_36550_, _36549_, _43152_);
  and (_36551_, _36550_, _36548_);
  or (_36552_, _36551_, _35035_);
  and (_43571_, _36552_, _41894_);
  not (_36553_, \oc8051_golden_model_1.PSW [1]);
  nor (_36554_, _43152_, _36553_);
  nor (_36556_, _05424_, _36553_);
  nor (_36557_, _08751_, _11709_);
  or (_36558_, _36557_, _36556_);
  or (_36559_, _36558_, _06572_);
  and (_36560_, _05424_, _04900_);
  or (_36561_, _36560_, _36556_);
  or (_36562_, _36561_, _04733_);
  or (_36563_, _05424_, \oc8051_golden_model_1.PSW [1]);
  and (_36564_, _12262_, _05424_);
  not (_36565_, _36564_);
  and (_36567_, _36565_, _36563_);
  or (_36568_, _36567_, _04722_);
  and (_36569_, _05424_, \oc8051_golden_model_1.ACC [1]);
  or (_36570_, _36569_, _36556_);
  and (_36571_, _36570_, _04707_);
  nor (_36572_, _04707_, _36553_);
  or (_36573_, _36572_, _03850_);
  or (_36574_, _36573_, _36571_);
  and (_36575_, _36574_, _03764_);
  and (_36576_, _36575_, _36568_);
  nor (_36578_, _06094_, _36553_);
  and (_36579_, _12249_, _06094_);
  or (_36580_, _36579_, _36578_);
  and (_36581_, _36580_, _03763_);
  or (_36582_, _36581_, _03848_);
  or (_36583_, _36582_, _36576_);
  and (_36584_, _36583_, _36562_);
  or (_36585_, _36584_, _03854_);
  or (_36586_, _36570_, _03855_);
  and (_36587_, _36586_, _03760_);
  and (_36589_, _36587_, _36585_);
  and (_36590_, _12252_, _06094_);
  or (_36591_, _36590_, _36578_);
  and (_36592_, _36591_, _03759_);
  or (_36593_, _36592_, _03752_);
  or (_36594_, _36593_, _36589_);
  and (_36595_, _36579_, _12248_);
  or (_36596_, _36578_, _03753_);
  or (_36597_, _36596_, _36595_);
  and (_36598_, _36597_, _03747_);
  and (_36600_, _36598_, _36594_);
  not (_36601_, _06094_);
  nor (_36602_, _12293_, _36601_);
  or (_36603_, _36602_, _36578_);
  and (_36604_, _36603_, _03746_);
  or (_36605_, _36604_, _08474_);
  or (_36606_, _36605_, _36600_);
  or (_36607_, _36561_, _07925_);
  and (_36608_, _36607_, _36606_);
  or (_36609_, _36608_, _03737_);
  and (_36611_, _06961_, _05424_);
  or (_36612_, _36556_, _03738_);
  or (_36613_, _36612_, _36611_);
  and (_36614_, _36613_, _03820_);
  and (_36615_, _36614_, _36609_);
  nor (_36616_, _12352_, _11709_);
  or (_36617_, _36616_, _36556_);
  and (_36618_, _36617_, _03455_);
  or (_36619_, _36618_, _36615_);
  and (_36620_, _36619_, _04778_);
  nand (_36622_, _05424_, _04595_);
  and (_36623_, _36563_, _03903_);
  and (_36624_, _36623_, _36622_);
  or (_36625_, _36624_, _36620_);
  and (_36626_, _36625_, _04790_);
  or (_36627_, _12366_, _11709_);
  and (_36628_, _36563_, _03897_);
  and (_36629_, _36628_, _36627_);
  or (_36630_, _36629_, _04018_);
  or (_36631_, _36630_, _36626_);
  nand (_36633_, _08750_, _05424_);
  and (_36634_, _36633_, _36558_);
  or (_36635_, _36634_, _04792_);
  and (_36636_, _36635_, _03909_);
  and (_36637_, _36636_, _36631_);
  or (_36638_, _12244_, _11709_);
  and (_36639_, _36563_, _03908_);
  and (_36640_, _36639_, _36638_);
  or (_36641_, _36640_, _04027_);
  or (_36642_, _36641_, _36637_);
  nor (_36644_, _36556_, _04785_);
  nand (_36645_, _36644_, _36633_);
  and (_36646_, _36645_, _06567_);
  and (_36647_, _36646_, _36642_);
  or (_36648_, _36622_, _08366_);
  and (_36649_, _36563_, _03914_);
  and (_36650_, _36649_, _36648_);
  or (_36651_, _36650_, _04011_);
  or (_36652_, _36651_, _36647_);
  and (_36653_, _36652_, _36559_);
  or (_36655_, _36653_, _03773_);
  or (_36656_, _36567_, _03774_);
  and (_36657_, _36656_, _03375_);
  and (_36658_, _36657_, _36655_);
  and (_36659_, _36591_, _03374_);
  or (_36660_, _36659_, _03772_);
  or (_36661_, _36660_, _36658_);
  or (_36662_, _36556_, _04060_);
  or (_36663_, _36662_, _36564_);
  and (_36664_, _36663_, _43152_);
  and (_36666_, _36664_, _36661_);
  or (_36667_, _36666_, _36554_);
  and (_43572_, _36667_, _41894_);
  and (_36668_, _43156_, \oc8051_golden_model_1.PSW [2]);
  nor (_36669_, _08726_, _36093_);
  and (_36670_, _08726_, _08525_);
  or (_36671_, _36670_, _36669_);
  and (_36672_, _36671_, _08691_);
  not (_36673_, _04435_);
  nor (_36674_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  nand (_36676_, _36674_, _07035_);
  nand (_36677_, _36676_, _07010_);
  nor (_36678_, _08250_, \oc8051_golden_model_1.ACC [7]);
  and (_36679_, _08250_, \oc8051_golden_model_1.ACC [7]);
  nor (_36680_, _36679_, _36678_);
  not (_36681_, _36680_);
  or (_36682_, _36681_, _11726_);
  nand (_36683_, _36681_, _11726_);
  and (_36684_, _36683_, _36682_);
  and (_36685_, _36684_, _08316_);
  nor (_36687_, _36684_, _08316_);
  or (_36688_, _36687_, _36685_);
  and (_36689_, _36688_, _04330_);
  and (_36690_, _36601_, \oc8051_golden_model_1.PSW [2]);
  and (_36691_, _12464_, _06094_);
  and (_36692_, _36691_, _12463_);
  or (_36693_, _36692_, _36690_);
  and (_36694_, _36693_, _03752_);
  and (_36695_, _12467_, _06094_);
  or (_36696_, _36695_, _36690_);
  and (_36698_, _36696_, _03759_);
  and (_36699_, _11709_, \oc8051_golden_model_1.PSW [2]);
  and (_36700_, _05424_, _05307_);
  or (_36701_, _36700_, _36699_);
  or (_36702_, _36701_, _04733_);
  nor (_36703_, _12471_, _11709_);
  or (_36704_, _36703_, _36699_);
  or (_36705_, _36704_, _04722_);
  and (_36706_, _05424_, \oc8051_golden_model_1.ACC [2]);
  or (_36707_, _36706_, _36699_);
  and (_36709_, _36707_, _04707_);
  and (_36710_, _04708_, \oc8051_golden_model_1.PSW [2]);
  or (_36711_, _36710_, _03850_);
  or (_36712_, _36711_, _36709_);
  and (_36713_, _36712_, _03764_);
  and (_36714_, _36713_, _36705_);
  or (_36715_, _36691_, _36690_);
  and (_36716_, _36715_, _03763_);
  or (_36717_, _36716_, _03848_);
  or (_36718_, _36717_, _36714_);
  and (_36720_, _36718_, _36702_);
  or (_36721_, _36720_, _03854_);
  or (_36722_, _36707_, _03855_);
  and (_36723_, _36722_, _03760_);
  and (_36724_, _36723_, _36721_);
  or (_36725_, _36724_, _36698_);
  and (_36726_, _36725_, _03753_);
  or (_36727_, _36726_, _36694_);
  and (_36728_, _36727_, _07405_);
  or (_36729_, _14343_, _14233_);
  or (_36731_, _36729_, _14455_);
  or (_36732_, _36731_, _14571_);
  or (_36733_, _36732_, _14686_);
  or (_36734_, _36733_, _14799_);
  or (_36735_, _36734_, _07911_);
  or (_36736_, _36735_, _14920_);
  and (_36737_, _36736_, _07399_);
  or (_36738_, _36737_, _15513_);
  or (_36739_, _36738_, _36728_);
  nor (_36740_, _08042_, _11988_);
  not (_36742_, _05568_);
  or (_36743_, _08042_, _36742_);
  and (_36744_, _36743_, _06554_);
  or (_36745_, _36744_, _36740_);
  nand (_36746_, _36745_, _11889_);
  or (_36747_, _36745_, _11889_);
  and (_36748_, _36747_, _36746_);
  nor (_36749_, _36748_, _35497_);
  and (_36750_, _36748_, _35497_);
  or (_36751_, _36750_, _36749_);
  or (_36753_, _36751_, _08153_);
  and (_36754_, _36753_, _08248_);
  and (_36755_, _36754_, _36739_);
  or (_36756_, _36755_, _36689_);
  and (_36757_, _36756_, _03888_);
  and (_36758_, _08325_, \oc8051_golden_model_1.ACC [7]);
  nor (_36759_, _08325_, \oc8051_golden_model_1.ACC [7]);
  or (_36760_, _36759_, _36758_);
  or (_36761_, _36760_, _11719_);
  nand (_36762_, _36760_, _11719_);
  and (_36764_, _36762_, _36761_);
  and (_36765_, _36764_, _08390_);
  nor (_36766_, _36764_, _08390_);
  or (_36767_, _36766_, _36765_);
  and (_36768_, _36767_, _03883_);
  or (_36769_, _36768_, _08320_);
  or (_36770_, _36769_, _36757_);
  not (_36771_, _11907_);
  not (_36772_, _08401_);
  and (_36773_, _08455_, _36772_);
  nand (_36775_, _36773_, _36771_);
  or (_36776_, _36773_, _36771_);
  and (_36777_, _36776_, _36775_);
  or (_36778_, _36777_, _08321_);
  and (_36779_, _36778_, _03747_);
  and (_36780_, _36779_, _36770_);
  nor (_36781_, _12514_, _36601_);
  or (_36782_, _36781_, _36690_);
  and (_36783_, _36782_, _03746_);
  or (_36784_, _36783_, _07927_);
  or (_36786_, _36784_, _36780_);
  and (_36787_, _06965_, _05424_);
  or (_36788_, _36699_, _03738_);
  or (_36789_, _36788_, _36787_);
  or (_36790_, _36701_, _07925_);
  and (_36791_, _36790_, _03820_);
  and (_36792_, _36791_, _36789_);
  and (_36793_, _36792_, _36786_);
  nor (_36794_, _12572_, _11709_);
  or (_36795_, _36794_, _36699_);
  and (_36797_, _36795_, _03455_);
  or (_36798_, _36797_, _07010_);
  or (_36799_, _36798_, _36793_);
  and (_36800_, _36799_, _36677_);
  or (_36801_, _36800_, _03903_);
  and (_36802_, _05424_, _06495_);
  or (_36803_, _36802_, _36699_);
  or (_36804_, _36803_, _04778_);
  and (_36805_, _36804_, _04790_);
  and (_36806_, _36805_, _36801_);
  and (_36808_, _12586_, _05424_);
  or (_36809_, _36808_, _36699_);
  and (_36810_, _36809_, _03897_);
  or (_36811_, _36810_, _36806_);
  and (_36812_, _36811_, _04792_);
  and (_36813_, _08748_, _05424_);
  or (_36814_, _36813_, _36699_);
  and (_36815_, _36814_, _04018_);
  or (_36816_, _36815_, _36812_);
  and (_36817_, _36816_, _03909_);
  or (_36819_, _36699_, _05765_);
  and (_36820_, _36803_, _03908_);
  and (_36821_, _36820_, _36819_);
  or (_36822_, _36821_, _36817_);
  and (_36823_, _36822_, _04785_);
  and (_36824_, _36707_, _04027_);
  and (_36825_, _36824_, _36819_);
  or (_36826_, _36825_, _03914_);
  or (_36827_, _36826_, _36823_);
  nor (_36828_, _12585_, _11709_);
  or (_36830_, _36699_, _06567_);
  or (_36831_, _36830_, _36828_);
  and (_36832_, _36831_, _06572_);
  and (_36833_, _36832_, _36827_);
  nor (_36834_, _08747_, _11709_);
  or (_36835_, _36834_, _36699_);
  and (_36836_, _36835_, _04011_);
  or (_36837_, _36836_, _08590_);
  or (_36838_, _36837_, _36833_);
  nand (_36839_, _08597_, _03420_);
  and (_36841_, _36740_, _08108_);
  nor (_36842_, _36745_, _11702_);
  nor (_36843_, _36842_, _36740_);
  and (_36844_, _36843_, _08111_);
  or (_36845_, _36844_, _36841_);
  or (_36846_, _36845_, _08119_);
  and (_36847_, _36846_, _36839_);
  and (_36848_, _36847_, _36838_);
  and (_36849_, _04760_, _03382_);
  and (_36850_, _36679_, _08620_);
  nor (_36852_, _36681_, _11965_);
  nor (_36853_, _36852_, _36679_);
  and (_36854_, _36853_, _08623_);
  or (_36855_, _36854_, _36850_);
  and (_36856_, _36855_, _36849_);
  or (_36857_, _36856_, _36848_);
  and (_36858_, _36857_, _36673_);
  and (_36859_, _36855_, _04435_);
  or (_36860_, _36859_, _04022_);
  or (_36861_, _36860_, _36858_);
  and (_36863_, _36758_, _08650_);
  nor (_36864_, _36760_, _11970_);
  nor (_36865_, _36864_, _36758_);
  and (_36866_, _36865_, _08653_);
  or (_36867_, _36866_, _36863_);
  or (_36868_, _36867_, _04023_);
  and (_36869_, _36868_, _08659_);
  and (_36870_, _36869_, _36861_);
  nand (_36871_, _08398_, \oc8051_golden_model_1.ACC [7]);
  nor (_36872_, _08398_, \oc8051_golden_model_1.ACC [7]);
  or (_36874_, _36872_, _11976_);
  and (_36875_, _36874_, _36871_);
  and (_36876_, _36875_, _08683_);
  nor (_36877_, _36875_, _08683_);
  or (_36878_, _36877_, _36876_);
  nand (_36879_, _36878_, _08627_);
  nand (_36880_, _36879_, _11984_);
  or (_36881_, _36880_, _36870_);
  nand (_36882_, _08034_, _11988_);
  and (_36883_, _11989_, _36882_);
  or (_36885_, _36883_, _11984_);
  and (_36886_, _36885_, _36881_);
  or (_36887_, _36886_, _04456_);
  or (_36888_, _36883_, _11987_);
  and (_36889_, _36888_, _10058_);
  and (_36890_, _36889_, _36887_);
  or (_36891_, _36890_, _36672_);
  and (_36892_, _36891_, _10056_);
  or (_36893_, _08765_, _06556_);
  and (_36894_, _12007_, _36893_);
  not (_36896_, _36040_);
  or (_36897_, _36896_, _08804_);
  and (_36898_, _36897_, _08733_);
  and (_36899_, _36898_, _12011_);
  or (_36900_, _36899_, _03773_);
  or (_36901_, _36900_, _36894_);
  or (_36902_, _36901_, _36892_);
  or (_36903_, _36704_, _03774_);
  and (_36904_, _36903_, _03375_);
  and (_36905_, _36904_, _36902_);
  and (_36907_, _36696_, _03374_);
  or (_36908_, _36907_, _03772_);
  or (_36909_, _36908_, _36905_);
  and (_36910_, _12642_, _05424_);
  or (_36911_, _36699_, _04060_);
  or (_36912_, _36911_, _36910_);
  and (_36913_, _36912_, _43152_);
  and (_36914_, _36913_, _36909_);
  or (_36915_, _36914_, _36668_);
  and (_43573_, _36915_, _41894_);
  nor (_36917_, _43152_, _05135_);
  nor (_36918_, _05424_, _05135_);
  nor (_36919_, _12681_, _11709_);
  or (_36920_, _36919_, _36918_);
  or (_36921_, _36920_, _04722_);
  and (_36922_, _05424_, \oc8051_golden_model_1.ACC [3]);
  or (_36923_, _36922_, _36918_);
  and (_36924_, _36923_, _04707_);
  nor (_36925_, _04707_, _05135_);
  or (_36926_, _36925_, _03850_);
  or (_36928_, _36926_, _36924_);
  and (_36929_, _36928_, _03764_);
  and (_36930_, _36929_, _36921_);
  nor (_36931_, _06094_, _05135_);
  and (_36932_, _12674_, _06094_);
  or (_36933_, _36932_, _36931_);
  and (_36934_, _36933_, _03763_);
  or (_36935_, _36934_, _03848_);
  or (_36936_, _36935_, _36930_);
  and (_36937_, _05424_, _05119_);
  or (_36939_, _36937_, _36918_);
  or (_36940_, _36939_, _04733_);
  and (_36941_, _36940_, _36936_);
  or (_36942_, _36941_, _03854_);
  or (_36943_, _36923_, _03855_);
  and (_36944_, _36943_, _03760_);
  and (_36945_, _36944_, _36942_);
  and (_36946_, _12667_, _06094_);
  or (_36947_, _36946_, _36931_);
  and (_36948_, _36947_, _03759_);
  or (_36950_, _36948_, _03752_);
  or (_36951_, _36950_, _36945_);
  or (_36952_, _36931_, _12673_);
  and (_36953_, _36952_, _36933_);
  or (_36954_, _36953_, _03753_);
  and (_36955_, _36954_, _03747_);
  and (_36956_, _36955_, _36951_);
  nor (_36957_, _12668_, _36601_);
  or (_36958_, _36957_, _36931_);
  and (_36959_, _36958_, _03746_);
  or (_36961_, _36959_, _07927_);
  or (_36962_, _36961_, _36956_);
  or (_36963_, _36939_, _07925_);
  and (_36964_, _06964_, _05424_);
  or (_36965_, _36918_, _03738_);
  or (_36966_, _36965_, _36964_);
  and (_36967_, _36966_, _36963_);
  and (_36968_, _36967_, _36962_);
  or (_36969_, _36968_, _03455_);
  nor (_36970_, _12775_, _11709_);
  or (_36972_, _36918_, _03820_);
  or (_36973_, _36972_, _36970_);
  and (_36974_, _36973_, _04778_);
  and (_36975_, _36974_, _36969_);
  and (_36976_, _05424_, _06345_);
  or (_36977_, _36976_, _36918_);
  and (_36978_, _36977_, _03903_);
  or (_36979_, _36978_, _03897_);
  or (_36980_, _36979_, _36975_);
  and (_36981_, _12789_, _05424_);
  or (_36983_, _36918_, _04790_);
  or (_36984_, _36983_, _36981_);
  and (_36985_, _36984_, _04792_);
  and (_36986_, _36985_, _36980_);
  and (_36987_, _10491_, _05424_);
  or (_36988_, _36987_, _36918_);
  and (_36989_, _36988_, _04018_);
  or (_36990_, _36989_, _36986_);
  and (_36991_, _36990_, _03909_);
  or (_36992_, _36918_, _05622_);
  and (_36994_, _36977_, _03908_);
  and (_36995_, _36994_, _36992_);
  or (_36996_, _36995_, _36991_);
  and (_36997_, _36996_, _04785_);
  and (_36998_, _36923_, _04027_);
  and (_36999_, _36998_, _36992_);
  or (_37000_, _36999_, _03914_);
  or (_37001_, _37000_, _36997_);
  nor (_37002_, _12788_, _11709_);
  or (_37003_, _36918_, _06567_);
  or (_37005_, _37003_, _37002_);
  and (_37006_, _37005_, _06572_);
  and (_37007_, _37006_, _37001_);
  nor (_37008_, _08742_, _11709_);
  or (_37009_, _37008_, _36918_);
  and (_37010_, _37009_, _04011_);
  or (_37011_, _37010_, _03773_);
  or (_37012_, _37011_, _37007_);
  or (_37013_, _36920_, _03774_);
  and (_37014_, _37013_, _03375_);
  and (_37016_, _37014_, _37012_);
  and (_37017_, _36947_, _03374_);
  or (_37018_, _37017_, _03772_);
  or (_37019_, _37018_, _37016_);
  and (_37020_, _12848_, _05424_);
  or (_37021_, _36918_, _04060_);
  or (_37022_, _37021_, _37020_);
  and (_37023_, _37022_, _43152_);
  and (_37024_, _37023_, _37019_);
  or (_37025_, _37024_, _36917_);
  and (_43574_, _37025_, _41894_);
  and (_37027_, _43156_, \oc8051_golden_model_1.PSW [4]);
  and (_37028_, _11709_, \oc8051_golden_model_1.PSW [4]);
  and (_37029_, _12997_, _05424_);
  or (_37030_, _37029_, _37028_);
  and (_37031_, _37030_, _03897_);
  and (_37032_, _06969_, _05424_);
  or (_37033_, _37028_, _03738_);
  or (_37034_, _37033_, _37032_);
  and (_37035_, _05950_, _05424_);
  or (_37037_, _37035_, _37028_);
  or (_37038_, _37037_, _07925_);
  nor (_37039_, _12891_, _11709_);
  or (_37040_, _37039_, _37028_);
  or (_37041_, _37040_, _04722_);
  and (_37042_, _05424_, \oc8051_golden_model_1.ACC [4]);
  or (_37043_, _37042_, _37028_);
  and (_37044_, _37043_, _04707_);
  and (_37045_, _04708_, \oc8051_golden_model_1.PSW [4]);
  or (_37046_, _37045_, _03850_);
  or (_37048_, _37046_, _37044_);
  and (_37049_, _37048_, _03764_);
  and (_37050_, _37049_, _37041_);
  and (_37051_, _36601_, \oc8051_golden_model_1.PSW [4]);
  and (_37052_, _12875_, _06094_);
  or (_37053_, _37052_, _37051_);
  and (_37054_, _37053_, _03763_);
  or (_37055_, _37054_, _03848_);
  or (_37056_, _37055_, _37050_);
  or (_37057_, _37037_, _04733_);
  and (_37059_, _37057_, _37056_);
  or (_37060_, _37059_, _03854_);
  or (_37061_, _37043_, _03855_);
  and (_37062_, _37061_, _03760_);
  and (_37063_, _37062_, _37060_);
  and (_37064_, _12870_, _06094_);
  or (_37065_, _37064_, _37051_);
  and (_37066_, _37065_, _03759_);
  or (_37067_, _37066_, _03752_);
  or (_37068_, _37067_, _37063_);
  or (_37070_, _37051_, _12874_);
  and (_37071_, _37070_, _37053_);
  or (_37072_, _37071_, _03753_);
  and (_37073_, _37072_, _03747_);
  and (_37074_, _37073_, _37068_);
  nor (_37075_, _12872_, _36601_);
  or (_37076_, _37075_, _37051_);
  and (_37077_, _37076_, _03746_);
  or (_37078_, _37077_, _08474_);
  or (_37079_, _37078_, _37074_);
  and (_37081_, _37079_, _37038_);
  or (_37082_, _37081_, _03737_);
  and (_37083_, _37082_, _37034_);
  or (_37084_, _37083_, _03455_);
  nor (_37085_, _12982_, _11709_);
  or (_37086_, _37085_, _37028_);
  or (_37087_, _37086_, _03820_);
  and (_37088_, _37087_, _37084_);
  or (_37089_, _37088_, _03903_);
  and (_37090_, _06456_, _05424_);
  or (_37092_, _37090_, _37028_);
  or (_37093_, _37092_, _04778_);
  and (_37094_, _37093_, _04790_);
  and (_37095_, _37094_, _37089_);
  or (_37096_, _37095_, _37031_);
  and (_37097_, _37096_, _04792_);
  and (_37098_, _08741_, _05424_);
  or (_37099_, _37098_, _37028_);
  and (_37100_, _37099_, _04018_);
  or (_37101_, _37100_, _37097_);
  and (_37103_, _37101_, _03909_);
  or (_37104_, _37028_, _08336_);
  and (_37105_, _37092_, _03908_);
  and (_37106_, _37105_, _37104_);
  or (_37107_, _37106_, _37103_);
  and (_37108_, _37107_, _04785_);
  and (_37109_, _37043_, _04027_);
  and (_37110_, _37109_, _37104_);
  or (_37111_, _37110_, _03914_);
  or (_37112_, _37111_, _37108_);
  nor (_37114_, _12996_, _11709_);
  or (_37115_, _37028_, _06567_);
  or (_37116_, _37115_, _37114_);
  and (_37117_, _37116_, _06572_);
  and (_37118_, _37117_, _37112_);
  nor (_37119_, _08740_, _11709_);
  or (_37120_, _37119_, _37028_);
  and (_37121_, _37120_, _04011_);
  or (_37122_, _37121_, _03773_);
  or (_37123_, _37122_, _37118_);
  or (_37125_, _37040_, _03774_);
  and (_37126_, _37125_, _03375_);
  and (_37127_, _37126_, _37123_);
  and (_37128_, _37065_, _03374_);
  or (_37129_, _37128_, _03772_);
  or (_37130_, _37129_, _37127_);
  and (_37131_, _13056_, _05424_);
  or (_37132_, _37028_, _04060_);
  or (_37133_, _37132_, _37131_);
  and (_37134_, _37133_, _43152_);
  and (_37136_, _37134_, _37130_);
  or (_37137_, _37136_, _37027_);
  and (_43575_, _37137_, _41894_);
  and (_37138_, _43156_, \oc8051_golden_model_1.PSW [5]);
  and (_37139_, _11709_, \oc8051_golden_model_1.PSW [5]);
  and (_37140_, _06447_, _05424_);
  or (_37141_, _37140_, _37139_);
  or (_37142_, _37141_, _04778_);
  nor (_37143_, _13090_, _11709_);
  or (_37144_, _37143_, _37139_);
  and (_37146_, _37144_, _03850_);
  and (_37147_, _04708_, \oc8051_golden_model_1.PSW [5]);
  and (_37148_, _05424_, \oc8051_golden_model_1.ACC [5]);
  or (_37149_, _37148_, _37139_);
  and (_37150_, _37149_, _04707_);
  or (_37151_, _37150_, _37147_);
  and (_37152_, _37151_, _04722_);
  or (_37153_, _37152_, _03857_);
  or (_37154_, _37153_, _37146_);
  and (_37155_, _36601_, \oc8051_golden_model_1.PSW [5]);
  and (_37157_, _13094_, _06094_);
  or (_37158_, _37157_, _37155_);
  or (_37159_, _37158_, _03764_);
  and (_37160_, _05857_, _05424_);
  or (_37161_, _37160_, _37139_);
  or (_37162_, _37161_, _04733_);
  and (_37163_, _37162_, _37159_);
  and (_37164_, _37163_, _37154_);
  or (_37165_, _37164_, _03854_);
  or (_37166_, _37149_, _03855_);
  and (_37168_, _37166_, _03760_);
  and (_37169_, _37168_, _37165_);
  and (_37170_, _13071_, _06094_);
  or (_37171_, _37170_, _37155_);
  and (_37172_, _37171_, _03759_);
  or (_37173_, _37172_, _03752_);
  or (_37174_, _37173_, _37169_);
  or (_37175_, _37155_, _13109_);
  and (_37176_, _37175_, _37158_);
  or (_37177_, _37176_, _03753_);
  and (_37179_, _37177_, _03747_);
  and (_37180_, _37179_, _37174_);
  nor (_37181_, _13073_, _36601_);
  or (_37182_, _37181_, _37155_);
  and (_37183_, _37182_, _03746_);
  or (_37184_, _37183_, _07927_);
  or (_37185_, _37184_, _37180_);
  and (_37186_, _06968_, _05424_);
  or (_37187_, _37139_, _03738_);
  or (_37188_, _37187_, _37186_);
  or (_37190_, _37161_, _07925_);
  and (_37191_, _37190_, _03820_);
  and (_37192_, _37191_, _37188_);
  and (_37193_, _37192_, _37185_);
  nor (_37194_, _13182_, _11709_);
  or (_37195_, _37194_, _37139_);
  and (_37196_, _37195_, _03455_);
  or (_37197_, _37196_, _03903_);
  or (_37198_, _37197_, _37193_);
  and (_37199_, _37198_, _37142_);
  or (_37201_, _37199_, _03897_);
  and (_37202_, _13196_, _05424_);
  or (_37203_, _37139_, _04790_);
  or (_37204_, _37203_, _37202_);
  and (_37205_, _37204_, _04792_);
  and (_37206_, _37205_, _37201_);
  and (_37207_, _10493_, _05424_);
  or (_37208_, _37207_, _37139_);
  and (_37209_, _37208_, _04018_);
  or (_37210_, _37209_, _37206_);
  and (_37212_, _37210_, _03909_);
  or (_37213_, _37139_, _08335_);
  and (_37214_, _37141_, _03908_);
  and (_37215_, _37214_, _37213_);
  or (_37216_, _37215_, _37212_);
  and (_37217_, _37216_, _04785_);
  and (_37218_, _37149_, _04027_);
  and (_37219_, _37218_, _37213_);
  or (_37220_, _37219_, _03914_);
  or (_37221_, _37220_, _37217_);
  nor (_37223_, _13195_, _11709_);
  or (_37224_, _37139_, _06567_);
  or (_37225_, _37224_, _37223_);
  and (_37226_, _37225_, _06572_);
  and (_37227_, _37226_, _37221_);
  nor (_37228_, _08738_, _11709_);
  or (_37229_, _37228_, _37139_);
  and (_37230_, _37229_, _04011_);
  or (_37231_, _37230_, _03773_);
  or (_37232_, _37231_, _37227_);
  or (_37234_, _37144_, _03774_);
  and (_37235_, _37234_, _03375_);
  and (_37236_, _37235_, _37232_);
  and (_37237_, _37171_, _03374_);
  or (_37238_, _37237_, _03772_);
  or (_37239_, _37238_, _37236_);
  and (_37240_, _13255_, _05424_);
  or (_37241_, _37139_, _04060_);
  or (_37242_, _37241_, _37240_);
  and (_37243_, _37242_, _43152_);
  and (_37245_, _37243_, _37239_);
  or (_37246_, _37245_, _37138_);
  and (_43576_, _37246_, _41894_);
  nor (_37247_, _43152_, _15880_);
  or (_37248_, _08028_, _07999_);
  not (_37249_, _08113_);
  or (_37250_, _08102_, _08064_);
  and (_37251_, _37250_, _37249_);
  nor (_37252_, _13401_, _11709_);
  nor (_37253_, _05424_, _15880_);
  or (_37255_, _37253_, _06567_);
  or (_37256_, _37255_, _37252_);
  and (_37257_, _13394_, _05424_);
  or (_37258_, _37257_, _37253_);
  or (_37259_, _37258_, _04778_);
  or (_37260_, _08064_, _04330_);
  or (_37261_, _37260_, _08140_);
  and (_37262_, _37261_, _15018_);
  nor (_37263_, _13293_, _11709_);
  or (_37264_, _37263_, _37253_);
  or (_37266_, _37264_, _04722_);
  and (_37267_, _05424_, \oc8051_golden_model_1.ACC [6]);
  or (_37268_, _37267_, _37253_);
  and (_37269_, _37268_, _04707_);
  nor (_37270_, _04707_, _15880_);
  or (_37271_, _37270_, _03850_);
  or (_37272_, _37271_, _37269_);
  and (_37273_, _37272_, _03764_);
  and (_37274_, _37273_, _37266_);
  nor (_37275_, _06094_, _15880_);
  and (_37277_, _13297_, _06094_);
  or (_37278_, _37277_, _37275_);
  and (_37279_, _37278_, _03763_);
  or (_37280_, _37279_, _03848_);
  or (_37281_, _37280_, _37274_);
  and (_37282_, _06065_, _05424_);
  or (_37283_, _37282_, _37253_);
  or (_37284_, _37283_, _04733_);
  and (_37285_, _37284_, _37281_);
  or (_37286_, _37285_, _03854_);
  or (_37288_, _37268_, _03855_);
  and (_37289_, _37288_, _03760_);
  and (_37290_, _37289_, _37286_);
  and (_37291_, _13277_, _06094_);
  or (_37292_, _37291_, _37275_);
  and (_37293_, _37292_, _03759_);
  or (_37294_, _37293_, _03752_);
  or (_37295_, _37294_, _37290_);
  or (_37296_, _37275_, _13312_);
  and (_37297_, _37296_, _37278_);
  or (_37299_, _37297_, _03753_);
  and (_37300_, _37299_, _08153_);
  and (_37301_, _37300_, _37295_);
  or (_37302_, _37301_, _37262_);
  or (_37303_, _08268_, _08248_);
  or (_37304_, _37303_, _08306_);
  and (_37305_, _37304_, _37302_);
  or (_37306_, _37305_, _10086_);
  or (_37307_, _08395_, _08321_);
  or (_37308_, _37307_, _08448_);
  and (_37310_, _37308_, _03747_);
  or (_37311_, _08337_, _03888_);
  or (_37312_, _37311_, _08380_);
  and (_37313_, _37312_, _37310_);
  and (_37314_, _37313_, _37306_);
  nor (_37315_, _13279_, _36601_);
  or (_37316_, _37315_, _37275_);
  and (_37317_, _37316_, _03746_);
  or (_37318_, _37317_, _07927_);
  or (_37319_, _37318_, _37314_);
  and (_37321_, _06641_, _05424_);
  or (_37322_, _37253_, _03738_);
  or (_37323_, _37322_, _37321_);
  or (_37324_, _37283_, _07925_);
  and (_37325_, _37324_, _03820_);
  and (_37326_, _37325_, _37323_);
  and (_37327_, _37326_, _37319_);
  nor (_37328_, _13387_, _11709_);
  or (_37329_, _37328_, _37253_);
  and (_37330_, _37329_, _03455_);
  or (_37332_, _37330_, _03903_);
  or (_37333_, _37332_, _37327_);
  and (_37334_, _37333_, _37259_);
  or (_37335_, _37334_, _03897_);
  and (_37336_, _13402_, _05424_);
  or (_37337_, _37336_, _37253_);
  or (_37338_, _37337_, _04790_);
  and (_37339_, _37338_, _04792_);
  and (_37340_, _37339_, _37335_);
  and (_37341_, _08736_, _05424_);
  or (_37343_, _37341_, _37253_);
  and (_37344_, _37343_, _04018_);
  or (_37345_, _37344_, _37340_);
  and (_37346_, _37345_, _03909_);
  or (_37347_, _37253_, _08322_);
  and (_37348_, _37258_, _03908_);
  and (_37349_, _37348_, _37347_);
  or (_37350_, _37349_, _37346_);
  and (_37351_, _37350_, _04785_);
  and (_37352_, _37268_, _04027_);
  and (_37354_, _37352_, _37347_);
  or (_37355_, _37354_, _03914_);
  or (_37356_, _37355_, _37351_);
  and (_37357_, _37356_, _37256_);
  or (_37358_, _37357_, _04011_);
  nor (_37359_, _08735_, _11709_);
  or (_37360_, _37359_, _37253_);
  or (_37361_, _37360_, _06572_);
  and (_37362_, _37361_, _08113_);
  and (_37363_, _37362_, _37358_);
  or (_37365_, _37363_, _37251_);
  and (_37366_, _37365_, _04221_);
  and (_37367_, _37250_, _04220_);
  or (_37368_, _37367_, _04616_);
  or (_37369_, _37368_, _37366_);
  or (_37370_, _37250_, _04617_);
  and (_37371_, _37370_, _37369_);
  or (_37372_, _37371_, _04432_);
  nor (_37373_, _37250_, _04433_);
  and (_37374_, _03719_, _03382_);
  nor (_37376_, _37374_, _37373_);
  nand (_37377_, _37376_, _37372_);
  nand (_37378_, _37374_, _37250_);
  and (_37379_, _37378_, _36839_);
  nand (_37380_, _37379_, _37377_);
  or (_37381_, _08614_, _08268_);
  or (_37382_, _37381_, _36839_);
  and (_37383_, _37382_, _36673_);
  and (_37384_, _37383_, _37380_);
  and (_37385_, _37381_, _04435_);
  or (_37387_, _37385_, _04022_);
  or (_37388_, _37387_, _37384_);
  or (_37389_, _08337_, _04023_);
  or (_37390_, _37389_, _08644_);
  and (_37391_, _37390_, _08659_);
  and (_37392_, _37391_, _37388_);
  or (_37393_, _08674_, _08395_);
  and (_37394_, _37393_, _08627_);
  or (_37395_, _37394_, _15460_);
  or (_37396_, _37395_, _37392_);
  and (_37398_, _37396_, _37248_);
  or (_37399_, _37398_, _08691_);
  or (_37400_, _08720_, _10058_);
  and (_37401_, _37400_, _04140_);
  and (_37402_, _37401_, _37399_);
  or (_37403_, _08759_, _08733_);
  and (_37404_, _37403_, _10057_);
  or (_37405_, _37404_, _37402_);
  or (_37406_, _08799_, _15201_);
  and (_37407_, _37406_, _37405_);
  or (_37409_, _37407_, _03773_);
  or (_37410_, _37264_, _03774_);
  and (_37411_, _37410_, _03375_);
  and (_37412_, _37411_, _37409_);
  and (_37413_, _37292_, _03374_);
  or (_37414_, _37413_, _03772_);
  or (_37415_, _37414_, _37412_);
  nor (_37416_, _13460_, _11709_);
  or (_37417_, _37253_, _04060_);
  or (_37418_, _37417_, _37416_);
  and (_37420_, _37418_, _43152_);
  and (_37421_, _37420_, _37415_);
  or (_37422_, _37421_, _37247_);
  and (_43577_, _37422_, _41894_);
  and (_37423_, _43156_, \oc8051_golden_model_1.P0INREG [0]);
  or (_37424_, _37423_, _01115_);
  and (_43580_, _37424_, _41894_);
  and (_37425_, _43156_, \oc8051_golden_model_1.P0INREG [1]);
  or (_37426_, _37425_, _01130_);
  and (_43581_, _37426_, _41894_);
  and (_37428_, _43156_, \oc8051_golden_model_1.P0INREG [2]);
  or (_37429_, _37428_, _01138_);
  and (_43582_, _37429_, _41894_);
  and (_37430_, _43156_, \oc8051_golden_model_1.P0INREG [3]);
  or (_37431_, _37430_, _01123_);
  and (_43583_, _37431_, _41894_);
  and (_37432_, _43156_, \oc8051_golden_model_1.P0INREG [4]);
  or (_37433_, _37432_, _01150_);
  and (_43584_, _37433_, _41894_);
  and (_37434_, _43156_, \oc8051_golden_model_1.P0INREG [5]);
  or (_37436_, _37434_, _01165_);
  and (_43587_, _37436_, _41894_);
  and (_37437_, _43156_, \oc8051_golden_model_1.P0INREG [6]);
  or (_37438_, _37437_, _01172_);
  and (_43588_, _37438_, _41894_);
  and (_37439_, _43156_, \oc8051_golden_model_1.P1INREG [0]);
  or (_37440_, _37439_, _01294_);
  and (_43589_, _37440_, _41894_);
  and (_37441_, _43156_, \oc8051_golden_model_1.P1INREG [1]);
  or (_37442_, _37441_, _01272_);
  and (_43591_, _37442_, _41894_);
  and (_37444_, _43156_, \oc8051_golden_model_1.P1INREG [2]);
  or (_37445_, _37444_, _01287_);
  and (_43592_, _37445_, _41894_);
  and (_37446_, _43156_, \oc8051_golden_model_1.P1INREG [3]);
  or (_37447_, _37446_, _01280_);
  and (_43593_, _37447_, _41894_);
  and (_37448_, _43156_, \oc8051_golden_model_1.P1INREG [4]);
  or (_37449_, _37448_, _01327_);
  and (_43594_, _37449_, _41894_);
  and (_37451_, _43156_, \oc8051_golden_model_1.P1INREG [5]);
  or (_37452_, _37451_, _01305_);
  and (_43595_, _37452_, _41894_);
  and (_37453_, _43156_, \oc8051_golden_model_1.P1INREG [6]);
  or (_37454_, _37453_, _01320_);
  and (_43596_, _37454_, _41894_);
  and (_37455_, _43156_, \oc8051_golden_model_1.P2INREG [0]);
  or (_37456_, _37455_, _01184_);
  and (_43599_, _37456_, _41894_);
  and (_37457_, _43156_, \oc8051_golden_model_1.P2INREG [1]);
  or (_37459_, _37457_, _01206_);
  and (_43600_, _37459_, _41894_);
  and (_37460_, _43156_, \oc8051_golden_model_1.P2INREG [2]);
  or (_37461_, _37460_, _01199_);
  and (_43601_, _37461_, _41894_);
  and (_37462_, _43156_, \oc8051_golden_model_1.P2INREG [3]);
  or (_37463_, _37462_, _01192_);
  and (_43602_, _37463_, _41894_);
  and (_37464_, _43156_, \oc8051_golden_model_1.P2INREG [4]);
  or (_37465_, _37464_, _01217_);
  and (_43603_, _37465_, _41894_);
  and (_37467_, _43156_, \oc8051_golden_model_1.P2INREG [5]);
  or (_37468_, _37467_, _01239_);
  and (_43604_, _37468_, _41894_);
  and (_37469_, _43156_, \oc8051_golden_model_1.P2INREG [6]);
  or (_37470_, _37469_, _01232_);
  and (_43605_, _37470_, _41894_);
  and (_37471_, _43156_, \oc8051_golden_model_1.P3INREG [0]);
  or (_37472_, _37471_, _01428_);
  and (_43607_, _37472_, _41894_);
  and (_37474_, _43156_, \oc8051_golden_model_1.P3INREG [1]);
  or (_37475_, _37474_, _01421_);
  and (_43608_, _37475_, _41894_);
  and (_37476_, _43156_, \oc8051_golden_model_1.P3INREG [2]);
  or (_37477_, _37476_, _01403_);
  and (_43609_, _37477_, _41894_);
  and (_37478_, _43156_, \oc8051_golden_model_1.P3INREG [3]);
  or (_37479_, _37478_, _01414_);
  and (_43610_, _37479_, _41894_);
  and (_37480_, _43156_, \oc8051_golden_model_1.P3INREG [4]);
  or (_37482_, _37480_, _01390_);
  and (_43611_, _37482_, _41894_);
  and (_37483_, _43156_, \oc8051_golden_model_1.P3INREG [5]);
  or (_37484_, _37483_, _01380_);
  and (_43612_, _37484_, _41894_);
  and (_37485_, _43156_, \oc8051_golden_model_1.P3INREG [6]);
  or (_37486_, _37485_, _01358_);
  and (_43613_, _37486_, _41894_);
  and (_00005_[6], _01359_, _41894_);
  and (_00005_[5], _01381_, _41894_);
  and (_00005_[4], _01391_, _41894_);
  and (_00005_[3], _01415_, _41894_);
  and (_00005_[2], _01404_, _41894_);
  and (_00005_[1], _01422_, _41894_);
  and (_00005_[0], _01429_, _41894_);
  and (_00004_[6], _01233_, _41894_);
  and (_00004_[5], _01240_, _41894_);
  and (_00004_[4], _01218_, _41894_);
  and (_00004_[3], _01193_, _41894_);
  and (_00004_[2], _01200_, _41894_);
  and (_00004_[1], _01207_, _41894_);
  and (_00004_[0], _01185_, _41894_);
  and (_00003_[6], _01321_, _41894_);
  and (_00003_[5], _01306_, _41894_);
  and (_00003_[4], _01328_, _41894_);
  and (_00003_[3], _01281_, _41894_);
  and (_00003_[2], _01288_, _41894_);
  and (_00003_[1], _01273_, _41894_);
  and (_00003_[0], _01295_, _41894_);
  and (_00002_[6], _01173_, _41894_);
  and (_00002_[5], _01166_, _41894_);
  and (_00002_[4], _01151_, _41894_);
  and (_00002_[3], _01124_, _41894_);
  and (_00002_[2], _01139_, _41894_);
  and (_00002_[1], _01131_, _41894_);
  and (_00002_[0], _01116_, _41894_);
  nor (_37490_, _21490_, _21146_);
  nor (_37491_, _21749_, _21576_);
  and (_37492_, _37491_, _37490_);
  nor (_37493_, _21061_, _20978_);
  nor (_37495_, _20894_, _20554_);
  and (_37496_, _37495_, _37493_);
  and (_37497_, _37496_, _37492_);
  nor (_37498_, _22882_, _22794_);
  not (_37499_, _22969_);
  and (_37500_, _23858_, _37499_);
  and (_37501_, _37500_, _37498_);
  nor (_37502_, _22185_, _22097_);
  nor (_37503_, _22707_, _22361_);
  and (_37504_, _37503_, _37502_);
  and (_37506_, _37504_, _37501_);
  and (_37507_, _37506_, _37497_);
  and (_37508_, _09556_, _09474_);
  not (_37509_, _17501_);
  and (_37510_, _37509_, _09636_);
  and (_37511_, _37510_, _37508_);
  and (_37512_, _09128_, _08942_);
  and (_37513_, _09393_, _09313_);
  and (_37514_, _37513_, _37512_);
  and (_37515_, _37514_, _37511_);
  not (_37517_, _19161_);
  and (_37518_, _19268_, _37517_);
  nor (_37519_, _20381_, _20294_);
  and (_37520_, _37519_, _37518_);
  nor (_37521_, _17763_, _17588_);
  nor (_37522_, _18986_, _18899_);
  and (_37523_, _37522_, _37521_);
  and (_37524_, _37523_, _37520_);
  and (_37525_, _37524_, _37515_);
  and (_37526_, _37525_, _37507_);
  nor (_37528_, _19495_, _18096_);
  nor (_37529_, _24083_, _23304_);
  nand (_37530_, _37529_, _37528_);
  nor (_37531_, _37530_, _18324_);
  and (_37532_, _37531_, _37526_);
  nor (_37533_, _19608_, _18210_);
  nor (_37534_, _24201_, _23417_);
  and (_37535_, _37534_, _37533_);
  not (_37536_, _17676_);
  and (_37537_, _17870_, _37536_);
  nor (_37539_, _19073_, _17983_);
  and (_37540_, _37539_, _37537_);
  nor (_37541_, _18812_, _18725_);
  nor (_37542_, _20208_, _20120_);
  and (_37543_, _37542_, _37541_);
  nor (_37544_, _21227_, _20636_);
  nor (_37545_, _22445_, _21833_);
  and (_37546_, _37545_, _37544_);
  or (_37547_, _04600_, _03178_);
  or (_37548_, _37547_, _10643_);
  nor (_37550_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor (_37551_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor (_37552_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and (_37553_, _37552_, _37551_);
  and (_37554_, _37553_, _37550_);
  nor (_37555_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_37556_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and (_37557_, _37556_, _37555_);
  nor (_37558_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor (_37559_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and (_37561_, _37559_, _37558_);
  and (_37562_, _37561_, _37557_);
  and (_37563_, _37562_, _37554_);
  nor (_37564_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor (_37565_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and (_37566_, _37565_, _37564_);
  nor (_37567_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor (_37568_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and (_37569_, _37568_, _37567_);
  and (_37570_, _37569_, _37566_);
  nor (_37572_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_37573_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and (_37574_, _37573_, _37572_);
  nor (_37575_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor (_37576_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and (_37577_, _37576_, _37575_);
  and (_37578_, _37577_, _37574_);
  and (_37579_, _37578_, _37570_);
  and (_37580_, _37579_, _37563_);
  nor (_37581_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor (_37583_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and (_37584_, _37583_, _37581_);
  nor (_37585_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_37586_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and (_37587_, _37586_, _37585_);
  and (_37588_, _37587_, _37584_);
  nor (_37589_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  nor (_37590_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  and (_37591_, _37590_, _37589_);
  nor (_37592_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor (_37594_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and (_37595_, _37594_, _37592_);
  and (_37596_, _37595_, _37591_);
  and (_37597_, _37596_, _37588_);
  nor (_37598_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_37599_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and (_37600_, _37599_, _37598_);
  nor (_37601_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  nor (_37602_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  and (_37603_, _37602_, _37601_);
  and (_37605_, _37603_, _37600_);
  nor (_37606_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor (_37607_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and (_37608_, _37607_, _37606_);
  nor (_37609_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor (_37610_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and (_37611_, _37610_, _37609_);
  and (_37612_, _37611_, _37608_);
  and (_37613_, _37612_, _37605_);
  and (_37614_, _37613_, _37597_);
  nor (_37616_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and (_37617_, _37616_, op0_cnst);
  nor (_37618_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor (_37619_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and (_37620_, _37619_, _37618_);
  nor (_37621_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor (_37622_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and (_37623_, _37622_, _37621_);
  and (_37624_, _37623_, _37620_);
  and (_37625_, _37624_, _37617_);
  nor (_37627_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_37628_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and (_37629_, _37628_, _37627_);
  nor (_37630_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor (_37631_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and (_37632_, _37631_, _37630_);
  and (_37633_, _37632_, _37629_);
  and (_37634_, \oc8051_golden_model_1.TCON [1], _19166_);
  nor (_37635_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and (_37636_, _37635_, _37634_);
  nor (_37638_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor (_37639_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and (_37640_, _37639_, _37638_);
  and (_37641_, _37640_, _37636_);
  and (_37642_, _37641_, _37633_);
  and (_37643_, _37642_, _37625_);
  and (_37644_, _37643_, _37614_);
  and (_37645_, _37644_, _37580_);
  nand (_37646_, _37645_, _37548_);
  nor (_37647_, _37646_, _17238_);
  nor (_37649_, _20033_, _18636_);
  and (_37650_, _37649_, _37647_);
  and (_37651_, _37650_, _37546_);
  nor (_37652_, _17414_, _17326_);
  and (_37653_, _37652_, _37651_);
  and (_37654_, _37653_, _37543_);
  nor (_37655_, _22620_, _22533_);
  nor (_37656_, _22010_, _21922_);
  and (_37657_, _37656_, _37655_);
  nor (_37658_, _20809_, _20723_);
  nor (_37660_, _21399_, _21312_);
  and (_37661_, _37660_, _37658_);
  and (_37662_, _37661_, _37657_);
  and (_37663_, _37662_, _37654_);
  and (_37664_, _37663_, _37540_);
  not (_37665_, _23076_);
  or (_37666_, _23191_, _37665_);
  nor (_37667_, _37666_, _23970_);
  not (_37668_, _20467_);
  and (_37669_, _37668_, _19381_);
  nor (_37671_, _22273_, _21662_);
  and (_37672_, _37671_, _37669_);
  and (_37673_, _37672_, _37667_);
  and (_37674_, _37673_, _37664_);
  and (_37675_, _37674_, _37535_);
  and (_37676_, _37675_, _37532_);
  nor (_37677_, _24313_, _23758_);
  nor (_37678_, _24539_, _24424_);
  and (_37679_, _37678_, _37677_);
  nor (_37680_, _19722_, _18552_);
  nor (_37682_, _23531_, _19950_);
  and (_37683_, _37682_, _37680_);
  and (_37684_, _37683_, _37679_);
  and (_37685_, _37684_, _37676_);
  or (_37686_, _19835_, _18439_);
  nor (_37687_, _37686_, _23644_);
  nor (_37688_, _09233_, _09048_);
  nor (_37689_, _09847_, _09741_);
  and (_37690_, _37689_, _37688_);
  and (_37691_, _37690_, _37687_);
  and (_37693_, _37691_, _37685_);
  or (_00001_, _37693_, rst);
  and (_00005_[7], _01373_, _41894_);
  and (_00004_[7], _01226_, _41894_);
  and (_00003_[7], _01314_, _41894_);
  and (_00002_[7], _01159_, _41894_);
  and (_37694_, _37693_, inst_finished_r);
  nor (_37695_, word_in[3], word_in[2]);
  not (_37696_, _37695_);
  not (_37697_, word_in[1]);
  and (_37699_, _37697_, word_in[0]);
  and (_37700_, _37699_, \oc8051_golden_model_1.IRAM[1] [0]);
  nor (_37701_, _37697_, word_in[0]);
  and (_37702_, _37701_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor (_37703_, _37702_, _37700_);
  nor (_37704_, word_in[1], word_in[0]);
  and (_37705_, _37704_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_37706_, word_in[1], word_in[0]);
  and (_37707_, _37706_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor (_37708_, _37707_, _37705_);
  and (_37710_, _37708_, _37703_);
  nor (_37711_, _37710_, _37696_);
  not (_37712_, word_in[3]);
  nor (_37713_, _37712_, word_in[2]);
  not (_37714_, _37713_);
  and (_37715_, _37699_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_37716_, _37701_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor (_37717_, _37716_, _37715_);
  and (_37718_, _37704_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_37719_, _37706_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor (_37721_, _37719_, _37718_);
  and (_37722_, _37721_, _37717_);
  nor (_37723_, _37722_, _37714_);
  nor (_37724_, _37723_, _37711_);
  and (_37725_, _37712_, word_in[2]);
  not (_37726_, _37725_);
  and (_37727_, _37699_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_37728_, _37701_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_37729_, _37728_, _37727_);
  and (_37730_, _37704_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_37732_, _37706_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_37733_, _37732_, _37730_);
  and (_37734_, _37733_, _37729_);
  nor (_37735_, _37734_, _37726_);
  and (_37736_, word_in[3], word_in[2]);
  not (_37737_, _37736_);
  and (_37738_, _37699_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_37739_, _37701_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor (_37740_, _37739_, _37738_);
  and (_37741_, _37704_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_37743_, _37706_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor (_37744_, _37743_, _37741_);
  and (_37745_, _37744_, _37740_);
  nor (_37746_, _37745_, _37737_);
  nor (_37747_, _37746_, _37735_);
  and (_37748_, _37747_, _37724_);
  and (_37749_, _37706_, _37725_);
  and (_37750_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_37751_, _37695_, _37706_);
  and (_37752_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_37754_, _37752_, _37750_);
  and (_37755_, _37736_, _37701_);
  and (_37756_, _37755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_37757_, _37713_, _37699_);
  and (_37758_, _37757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_37759_, _37758_, _37756_);
  and (_37760_, _37759_, _37754_);
  and (_37761_, _37701_, _37725_);
  and (_37762_, _37761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_37763_, _37699_, _37725_);
  and (_37765_, _37763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_37766_, _37765_, _37762_);
  and (_37767_, _37704_, _37725_);
  and (_37768_, _37767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_37769_, _37695_, _37699_);
  and (_37770_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_37771_, _37770_, _37768_);
  and (_37772_, _37771_, _37766_);
  and (_37773_, _37772_, _37760_);
  and (_37774_, _37736_, _37699_);
  and (_37776_, _37774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_37777_, _37713_, _37706_);
  and (_37778_, _37777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_37779_, _37778_, _37776_);
  and (_37780_, _37736_, _37706_);
  and (_37781_, _37780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_37782_, _37736_, _37704_);
  and (_37783_, _37782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_37784_, _37783_, _37781_);
  and (_37785_, _37784_, _37779_);
  and (_37787_, _37695_, _37704_);
  and (_37788_, _37787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_37789_, _37695_, _37701_);
  and (_37790_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_37791_, _37790_, _37788_);
  and (_37792_, _37713_, _37701_);
  and (_37793_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_37794_, _37713_, _37704_);
  and (_37795_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_37796_, _37795_, _37793_);
  and (_37798_, _37796_, _37791_);
  and (_37799_, _37798_, _37785_);
  and (_37800_, _37799_, _37773_);
  nand (_37801_, _37800_, _37748_);
  or (_37802_, _37800_, _37748_);
  and (_37803_, _37802_, _37801_);
  and (_37804_, _37699_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_37805_, _37701_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor (_37806_, _37805_, _37804_);
  and (_37807_, _37704_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_37809_, _37706_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor (_37810_, _37809_, _37807_);
  and (_37811_, _37810_, _37806_);
  nor (_37812_, _37811_, _37696_);
  and (_37813_, _37699_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_37814_, _37701_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor (_37815_, _37814_, _37813_);
  and (_37816_, _37704_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_37817_, _37706_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor (_37818_, _37817_, _37816_);
  and (_37820_, _37818_, _37815_);
  nor (_37821_, _37820_, _37737_);
  nor (_37822_, _37821_, _37812_);
  and (_37823_, _37699_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_37824_, _37701_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor (_37825_, _37824_, _37823_);
  and (_37826_, _37704_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_37827_, _37706_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_37828_, _37827_, _37826_);
  and (_37829_, _37828_, _37825_);
  nor (_37831_, _37829_, _37726_);
  and (_37832_, _37699_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_37833_, _37701_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor (_37834_, _37833_, _37832_);
  and (_37835_, _37704_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_37836_, _37706_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor (_37837_, _37836_, _37835_);
  and (_37838_, _37837_, _37834_);
  nor (_37839_, _37838_, _37714_);
  nor (_37840_, _37839_, _37831_);
  and (_37842_, _37840_, _37822_);
  and (_37843_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37844_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_37845_, _37844_, _37843_);
  and (_37846_, _37774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_37847_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_37848_, _37847_, _37846_);
  and (_37849_, _37848_, _37845_);
  and (_37850_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_37851_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_37853_, _37851_, _37850_);
  and (_37854_, _37763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_37855_, _37767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_37856_, _37855_, _37854_);
  and (_37857_, _37856_, _37853_);
  and (_37858_, _37857_, _37849_);
  and (_37859_, _37777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_37860_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_37861_, _37860_, _37859_);
  and (_37862_, _37755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_37864_, _37757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_37865_, _37864_, _37862_);
  and (_37866_, _37865_, _37861_);
  and (_37867_, _37761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_37868_, _37787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_37869_, _37868_, _37867_);
  and (_37870_, _37780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_37871_, _37782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_37872_, _37871_, _37870_);
  and (_37873_, _37872_, _37869_);
  and (_37875_, _37873_, _37866_);
  and (_37876_, _37875_, _37858_);
  nand (_37877_, _37876_, _37842_);
  or (_37878_, _37876_, _37842_);
  and (_37879_, _37878_, _37877_);
  or (_37880_, _37879_, _37803_);
  and (_37881_, _37699_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_37882_, _37701_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_37883_, _37882_, _37881_);
  and (_37884_, _37704_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_37886_, _37706_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor (_37887_, _37886_, _37884_);
  and (_37888_, _37887_, _37883_);
  nor (_37889_, _37888_, _37726_);
  and (_37890_, _37699_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_37891_, _37701_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor (_37892_, _37891_, _37890_);
  and (_37893_, _37704_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_37894_, _37706_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor (_37895_, _37894_, _37893_);
  and (_37897_, _37895_, _37892_);
  nor (_37898_, _37897_, _37737_);
  nor (_37899_, _37898_, _37889_);
  and (_37900_, _37699_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_37901_, _37701_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor (_37902_, _37901_, _37900_);
  and (_37903_, _37704_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_37904_, _37706_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor (_37905_, _37904_, _37903_);
  and (_37906_, _37905_, _37902_);
  nor (_37908_, _37906_, _37696_);
  and (_37909_, _37699_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_37910_, _37701_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor (_37911_, _37910_, _37909_);
  and (_37912_, _37704_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_37913_, _37706_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor (_37914_, _37913_, _37912_);
  and (_37915_, _37914_, _37911_);
  nor (_37916_, _37915_, _37714_);
  nor (_37917_, _37916_, _37908_);
  and (_37919_, _37917_, _37899_);
  and (_37920_, _37761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_37921_, _37763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_37922_, _37921_, _37920_);
  and (_37923_, _37780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_37924_, _37777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_37925_, _37924_, _37923_);
  and (_37926_, _37925_, _37922_);
  and (_37927_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_37928_, _37757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_37930_, _37928_, _37927_);
  and (_37931_, _37774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_37932_, _37782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_37933_, _37932_, _37931_);
  and (_37934_, _37933_, _37930_);
  and (_37935_, _37934_, _37926_);
  and (_37936_, _37787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_37937_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_37938_, _37937_, _37936_);
  and (_37939_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_37941_, _37767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_37942_, _37941_, _37939_);
  and (_37943_, _37942_, _37938_);
  and (_37944_, _37755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_37945_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_37946_, _37945_, _37944_);
  and (_37947_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_37948_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_37949_, _37948_, _37947_);
  and (_37950_, _37949_, _37946_);
  and (_37952_, _37950_, _37943_);
  and (_37953_, _37952_, _37935_);
  nand (_37954_, _37953_, _37919_);
  or (_37955_, _37953_, _37919_);
  and (_37956_, _37955_, _37954_);
  and (_37957_, _37699_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_37958_, _37701_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor (_37959_, _37958_, _37957_);
  and (_37960_, _37704_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_37961_, _37706_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor (_37963_, _37961_, _37960_);
  and (_37964_, _37963_, _37959_);
  nor (_37965_, _37964_, _37726_);
  and (_37966_, _37699_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_37967_, _37701_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor (_37968_, _37967_, _37966_);
  and (_37969_, _37704_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_37970_, _37706_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor (_37971_, _37970_, _37969_);
  and (_37972_, _37971_, _37968_);
  nor (_37974_, _37972_, _37714_);
  nor (_37975_, _37974_, _37965_);
  and (_37976_, _37699_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_37977_, _37701_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor (_37978_, _37977_, _37976_);
  and (_37979_, _37704_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_37980_, _37706_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor (_37981_, _37980_, _37979_);
  and (_37982_, _37981_, _37978_);
  nor (_37983_, _37982_, _37696_);
  and (_37985_, _37699_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_37986_, _37701_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor (_37987_, _37986_, _37985_);
  and (_37988_, _37704_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_37989_, _37706_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor (_37990_, _37989_, _37988_);
  and (_37991_, _37990_, _37987_);
  nor (_37992_, _37991_, _37737_);
  nor (_37993_, _37992_, _37983_);
  and (_37994_, _37993_, _37975_);
  not (_37996_, _37994_);
  and (_37997_, _37767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_37998_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_37999_, _37998_, _37997_);
  and (_38000_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_38001_, _37761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_38002_, _38001_, _38000_);
  and (_38003_, _38002_, _37999_);
  and (_38004_, _37774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_38005_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_38007_, _38005_, _38004_);
  and (_38008_, _37780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_38009_, _37782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_38010_, _38009_, _38008_);
  and (_38011_, _38010_, _38007_);
  and (_38012_, _38011_, _38003_);
  and (_38013_, _37757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_38014_, _37787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_38015_, _38014_, _38013_);
  and (_38016_, _37777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_38018_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_38019_, _38018_, _38016_);
  and (_38020_, _38019_, _38015_);
  and (_38021_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_38022_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_38023_, _38022_, _38021_);
  and (_38024_, _37755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_38025_, _37763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_38026_, _38025_, _38024_);
  and (_38027_, _38026_, _38023_);
  and (_38029_, _38027_, _38020_);
  and (_38030_, _38029_, _38012_);
  nor (_38031_, _38030_, _37996_);
  and (_38032_, _38030_, _37996_);
  or (_38033_, _38032_, _38031_);
  or (_38034_, _38033_, _37956_);
  or (_38035_, _38034_, _37880_);
  and (_38036_, _37699_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_38037_, _37701_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor (_38038_, _38037_, _38036_);
  and (_38040_, _37704_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_38041_, _37706_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor (_38042_, _38041_, _38040_);
  and (_38043_, _38042_, _38038_);
  nor (_38044_, _38043_, _37726_);
  and (_38045_, _37699_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_38046_, _37701_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor (_38047_, _38046_, _38045_);
  and (_38048_, _37704_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_38049_, _37706_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor (_38051_, _38049_, _38048_);
  and (_38052_, _38051_, _38047_);
  nor (_38053_, _38052_, _37737_);
  nor (_38054_, _38053_, _38044_);
  and (_38055_, _37699_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_38056_, _37701_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor (_38057_, _38056_, _38055_);
  and (_38058_, _37704_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_38059_, _37706_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor (_38060_, _38059_, _38058_);
  and (_38062_, _38060_, _38057_);
  nor (_38063_, _38062_, _37696_);
  and (_38064_, _37699_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_38065_, _37701_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor (_38066_, _38065_, _38064_);
  and (_38067_, _37704_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_38068_, _37706_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor (_38069_, _38068_, _38067_);
  and (_38070_, _38069_, _38066_);
  nor (_38071_, _38070_, _37714_);
  nor (_38073_, _38071_, _38063_);
  and (_38074_, _38073_, _38054_);
  and (_38075_, _37774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_38076_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_38077_, _38076_, _38075_);
  and (_38078_, _37763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_38079_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_38080_, _38079_, _38078_);
  and (_38081_, _38080_, _38077_);
  and (_38082_, _37777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_38084_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_38085_, _38084_, _38082_);
  and (_38086_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_38087_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_38088_, _38087_, _38086_);
  and (_38089_, _38088_, _38085_);
  and (_38090_, _38089_, _38081_);
  and (_38091_, _37761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_38092_, _37767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_38093_, _38092_, _38091_);
  and (_38095_, _37780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_38096_, _37787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_38097_, _38096_, _38095_);
  and (_38098_, _38097_, _38093_);
  and (_38099_, _37755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_38100_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_38101_, _38100_, _38099_);
  and (_38102_, _37782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_38103_, _37757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_38104_, _38103_, _38102_);
  and (_38106_, _38104_, _38101_);
  and (_38107_, _38106_, _38098_);
  and (_38108_, _38107_, _38090_);
  nand (_38109_, _38108_, _38074_);
  or (_38110_, _38108_, _38074_);
  and (_38111_, _38110_, _38109_);
  and (_38112_, _37699_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_38113_, _37701_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor (_38114_, _38113_, _38112_);
  and (_38115_, _37704_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_38117_, _37706_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor (_38118_, _38117_, _38115_);
  and (_38119_, _38118_, _38114_);
  nor (_38120_, _38119_, _37726_);
  and (_38121_, _37699_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_38122_, _37701_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor (_38123_, _38122_, _38121_);
  and (_38124_, _37704_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_38125_, _37706_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor (_38126_, _38125_, _38124_);
  and (_38128_, _38126_, _38123_);
  nor (_38129_, _38128_, _37737_);
  nor (_38130_, _38129_, _38120_);
  and (_38131_, _37699_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_38132_, _37701_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor (_38133_, _38132_, _38131_);
  and (_38134_, _37704_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_38135_, _37706_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor (_38136_, _38135_, _38134_);
  and (_38137_, _38136_, _38133_);
  nor (_38139_, _38137_, _37696_);
  and (_38140_, _37699_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_38141_, _37701_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor (_38142_, _38141_, _38140_);
  and (_38143_, _37704_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_38144_, _37706_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor (_38145_, _38144_, _38143_);
  and (_38146_, _38145_, _38142_);
  nor (_38147_, _38146_, _37714_);
  nor (_38148_, _38147_, _38139_);
  and (_38150_, _38148_, _38130_);
  and (_38151_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_38152_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_38153_, _38152_, _38151_);
  and (_38154_, _37780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_38155_, _37757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_38156_, _38155_, _38154_);
  and (_38157_, _38156_, _38153_);
  and (_38158_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_38159_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_38161_, _38159_, _38158_);
  and (_38162_, _37763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_38163_, _37767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_38164_, _38163_, _38162_);
  and (_38165_, _38164_, _38161_);
  and (_38166_, _38165_, _38157_);
  and (_38167_, _37782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_38168_, _37777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_38169_, _38168_, _38167_);
  and (_38170_, _37755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_38172_, _37774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_38173_, _38172_, _38170_);
  and (_38174_, _38173_, _38169_);
  and (_38175_, _37761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_38176_, _37787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_38177_, _38176_, _38175_);
  and (_38178_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_38179_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_38180_, _38179_, _38178_);
  and (_38181_, _38180_, _38177_);
  and (_38183_, _38181_, _38174_);
  and (_38184_, _38183_, _38166_);
  nand (_38185_, _38184_, _38150_);
  or (_38186_, _38184_, _38150_);
  and (_38187_, _38186_, _38185_);
  or (_38188_, _38187_, _38111_);
  and (_38189_, _37699_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_38190_, _37701_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor (_38191_, _38190_, _38189_);
  and (_38192_, _37704_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_38194_, _37706_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor (_38195_, _38194_, _38192_);
  and (_38196_, _38195_, _38191_);
  nor (_38197_, _38196_, _37726_);
  and (_38198_, _37699_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_38199_, _37701_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_38200_, _38199_, _38198_);
  and (_38201_, _37704_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_38202_, _37706_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor (_38203_, _38202_, _38201_);
  and (_38205_, _38203_, _38200_);
  nor (_38206_, _38205_, _37737_);
  nor (_38207_, _38206_, _38197_);
  and (_38208_, _37699_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_38209_, _37701_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor (_38210_, _38209_, _38208_);
  and (_38211_, _37704_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_38212_, _37706_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor (_38213_, _38212_, _38211_);
  and (_38214_, _38213_, _38210_);
  nor (_38216_, _38214_, _37696_);
  and (_38217_, _37699_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_38218_, _37701_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor (_38219_, _38218_, _38217_);
  and (_38220_, _37704_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_38221_, _37706_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_38222_, _38221_, _38220_);
  and (_38223_, _38222_, _38219_);
  nor (_38224_, _38223_, _37714_);
  nor (_38225_, _38224_, _38216_);
  and (_38227_, _38225_, _38207_);
  and (_38228_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_38229_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_38230_, _38229_, _38228_);
  and (_38231_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_38232_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_38233_, _38232_, _38231_);
  and (_38234_, _38233_, _38230_);
  and (_38235_, _37774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_38236_, _37782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor (_38238_, _38236_, _38235_);
  and (_38239_, _37763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_38240_, _37767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_38241_, _38240_, _38239_);
  and (_38242_, _38241_, _38238_);
  and (_38243_, _38242_, _38234_);
  and (_38244_, _37755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_38245_, _37777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_38246_, _38245_, _38244_);
  and (_38247_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_38249_, _37787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_38250_, _38249_, _38247_);
  and (_38251_, _38250_, _38246_);
  and (_38252_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_38253_, _37757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_38254_, _38253_, _38252_);
  and (_38255_, _37780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_38256_, _37761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_38257_, _38256_, _38255_);
  and (_38258_, _38257_, _38254_);
  and (_38260_, _38258_, _38251_);
  and (_38261_, _38260_, _38243_);
  or (_38262_, _38261_, _38227_);
  nand (_38263_, _38261_, _38227_);
  and (_38264_, _38263_, _38262_);
  and (_38265_, _37699_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_38266_, _37701_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor (_38267_, _38266_, _38265_);
  and (_38268_, _37704_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_38269_, _37706_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor (_38271_, _38269_, _38268_);
  and (_38272_, _38271_, _38267_);
  nor (_38273_, _38272_, _37696_);
  and (_38274_, _37699_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_38275_, _37701_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor (_38276_, _38275_, _38274_);
  and (_38277_, _37704_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_38278_, _37706_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor (_38279_, _38278_, _38277_);
  and (_38280_, _38279_, _38276_);
  nor (_38282_, _38280_, _37714_);
  nor (_38283_, _38282_, _38273_);
  and (_38284_, _37699_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_38285_, _37701_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor (_38286_, _38285_, _38284_);
  and (_38287_, _37704_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_38288_, _37706_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor (_38289_, _38288_, _38287_);
  and (_38290_, _38289_, _38286_);
  nor (_38291_, _38290_, _37726_);
  and (_38293_, _37699_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_38294_, _37701_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_38295_, _38294_, _38293_);
  and (_38296_, _37704_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_38297_, _37706_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_38298_, _38297_, _38296_);
  and (_38299_, _38298_, _38295_);
  nor (_38300_, _38299_, _37737_);
  nor (_38301_, _38300_, _38291_);
  and (_38302_, _38301_, _38283_);
  and (_38304_, _37782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_38305_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_38306_, _38305_, _38304_);
  and (_38307_, _37774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_38308_, _37749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_38309_, _38308_, _38307_);
  and (_38310_, _38309_, _38306_);
  and (_38311_, _37755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_38312_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_38313_, _38312_, _38311_);
  and (_38315_, _37787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_38316_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_38317_, _38316_, _38315_);
  and (_38318_, _38317_, _38313_);
  and (_38319_, _38318_, _38310_);
  and (_38320_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_38321_, _37767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_38322_, _38321_, _38320_);
  and (_38323_, _37780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_38324_, _37777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_38326_, _38324_, _38323_);
  and (_38327_, _38326_, _38322_);
  and (_38328_, _37757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_38329_, _37761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_38330_, _38329_, _38328_);
  and (_38331_, _37763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_38332_, _37751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_38333_, _38332_, _38331_);
  and (_38334_, _38333_, _38330_);
  and (_38335_, _38334_, _38327_);
  and (_38337_, _38335_, _38319_);
  not (_38338_, _38337_);
  nor (_38339_, _38338_, _38302_);
  and (_38340_, _38338_, _38302_);
  or (_38341_, _38340_, _38339_);
  or (_38342_, _38341_, _38264_);
  or (_38343_, _38342_, _38188_);
  or (_38344_, _38343_, _38035_);
  and (property_invalid_iram, _38344_, _37694_);
  nand (_38345_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38347_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38348_, _38347_, _38345_);
  and (_38349_, _07190_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_38350_, _07190_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_38351_, _38350_, _38349_);
  or (_38352_, _38351_, _38348_);
  nor (_38353_, _03474_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38354_, _03474_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_38355_, _38354_, _38353_);
  and (_38356_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38358_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_38359_, _38358_, _38356_);
  or (_38360_, _38359_, _38355_);
  or (_38361_, _38360_, _38352_);
  or (_38362_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38363_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38364_, _38363_, _38362_);
  or (_38365_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_38366_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38367_, _38366_, _38365_);
  or (_38369_, _38367_, _38364_);
  and (_38370_, _07036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_38371_, _07036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_38372_, _38371_, _38370_);
  nand (_38373_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38374_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_38375_, _38374_, _38373_);
  or (_38376_, _38375_, _38372_);
  or (_38377_, _38376_, _38369_);
  or (_38378_, _38377_, _38361_);
  and (property_invalid_acc, _38378_, _37694_);
  nor (_38380_, _28262_, _44086_);
  nor (_38381_, _26849_, _44070_);
  and (_38382_, _28262_, _44086_);
  or (_38383_, _38382_, _38381_);
  or (_38384_, _38383_, _38380_);
  and (_38385_, _27555_, _44078_);
  nor (_38386_, _28622_, _44090_);
  nor (_38387_, _27204_, _44074_);
  and (_38388_, _27204_, _44074_);
  or (_38390_, _38388_, _38387_);
  or (_38391_, _38390_, _38386_);
  and (_38392_, _27917_, _44082_);
  and (_38393_, _29289_, _38645_);
  nor (_38394_, _29289_, _38645_);
  nand (_38395_, _28951_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_38396_, _28951_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38397_, _38396_, _38395_);
  nor (_38398_, _29929_, _38635_);
  or (_38399_, _26100_, _44062_);
  nand (_38401_, _26100_, _44062_);
  and (_38402_, _38401_, _38399_);
  and (_38403_, _29929_, _38635_);
  or (_38404_, _38403_, _38402_);
  or (_38405_, _38404_, _38398_);
  and (_38406_, _30581_, _38631_);
  nor (_38407_, _30581_, _38631_);
  or (_38408_, _38407_, _38406_);
  or (_38409_, _38408_, _38405_);
  nor (_38410_, _10981_, _38667_);
  and (_38412_, _10981_, _38667_);
  or (_38413_, _38412_, _38410_);
  or (_38414_, _38413_, _38409_);
  and (_38415_, _30243_, _38656_);
  nor (_38416_, _30243_, _38656_);
  or (_38417_, _38416_, _38415_);
  or (_38418_, _38417_, _38414_);
  and (_38419_, _30882_, _38662_);
  nor (_38420_, _30882_, _38662_);
  or (_38421_, _38420_, _38419_);
  or (_38422_, _38421_, _38418_);
  and (_38423_, _29600_, _38650_);
  nor (_38424_, _29600_, _38650_);
  or (_38425_, _38424_, _38423_);
  or (_38426_, _38425_, _38422_);
  or (_38427_, _38426_, _38397_);
  or (_38428_, _38427_, _38394_);
  or (_38429_, _38428_, _38393_);
  or (_38430_, _38429_, _38392_);
  nor (_38431_, _27917_, _44082_);
  and (_38433_, _28622_, _44090_);
  or (_38434_, _38433_, _38431_);
  or (_38435_, _38434_, _38430_);
  or (_38436_, _38435_, _38391_);
  or (_38437_, _38436_, _38385_);
  nor (_38438_, _27555_, _44078_);
  and (_38439_, _26849_, _44070_);
  or (_38440_, _38439_, _38438_);
  or (_38441_, _38440_, _38437_);
  or (_38442_, _38441_, _38384_);
  and (_38444_, _26475_, _44066_);
  nor (_38445_, _26475_, _44066_);
  or (_38446_, _38445_, _38444_);
  or (_38447_, _38446_, _38442_);
  and (_38448_, _37693_, _43152_);
  and (property_invalid_pc, _38448_, _38447_);
  buf (_01385_, _41894_);
  buf (_01438_, _41894_);
  buf (_01491_, _41894_);
  buf (_01543_, _41894_);
  buf (_01595_, _41894_);
  buf (_01647_, _41894_);
  buf (_01698_, _41894_);
  buf (_01750_, _41894_);
  buf (_01802_, _41894_);
  buf (_01853_, _41894_);
  buf (_01892_, _41894_);
  buf (_01945_, _41894_);
  buf (_01998_, _41894_);
  buf (_02049_, _41894_);
  buf (_02101_, _41894_);
  buf (_02153_, _41894_);
  buf (_38964_, _38866_);
  buf (_38965_, _38867_);
  buf (_38978_, _38866_);
  buf (_38979_, _38867_);
  buf (_39292_, _38886_);
  buf (_39293_, _38888_);
  buf (_39294_, _38889_);
  buf (_39295_, _38890_);
  buf (_39296_, _38891_);
  buf (_39297_, _38892_);
  buf (_39298_, _38894_);
  buf (_39300_, _38895_);
  buf (_39301_, _38896_);
  buf (_39302_, _38897_);
  buf (_39303_, _38898_);
  buf (_39304_, _38900_);
  buf (_39305_, _38901_);
  buf (_39306_, _38902_);
  buf (_39357_, _38886_);
  buf (_39358_, _38888_);
  buf (_39359_, _38889_);
  buf (_39360_, _38890_);
  buf (_39361_, _38891_);
  buf (_39362_, _38892_);
  buf (_39363_, _38894_);
  buf (_39365_, _38895_);
  buf (_39366_, _38896_);
  buf (_39367_, _38897_);
  buf (_39368_, _38898_);
  buf (_39369_, _38900_);
  buf (_39370_, _38901_);
  buf (_39371_, _38902_);
  buf (_39764_, _39668_);
  buf (_39879_, _39668_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _01389_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _01393_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _01397_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _01401_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _01405_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _01409_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _01413_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _01382_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _01385_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _01442_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _01446_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _01450_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _01454_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _01458_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _01462_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _01466_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _01435_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _01438_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _01896_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _01900_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _01904_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _01908_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _01912_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _01916_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _01920_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _01889_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _01892_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _01949_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _01953_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _01957_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _01961_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _01965_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _01969_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _01973_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _01942_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _01945_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _02001_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _02005_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _02009_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _02013_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _02017_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _02021_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _02025_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _01995_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _01998_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _02053_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _02057_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _02061_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _02065_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _02069_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _02073_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _02076_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _02046_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _02049_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _02105_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _02109_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _02112_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _02116_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _02120_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _02124_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _02128_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _02098_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _02101_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _02157_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _02161_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _02164_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _02168_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _02172_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _02176_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _02180_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _02150_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _02153_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _01495_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _01499_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _01503_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _01507_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _01511_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _01515_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _01519_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _01488_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _01491_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _01547_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _01551_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _01555_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _01559_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _01562_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _01566_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _01570_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _01540_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _01543_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _01599_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _01603_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _01607_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _01611_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _01615_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _01619_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _01622_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _01592_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _01595_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _01651_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _01655_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _01659_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _01662_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _01666_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _01670_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _01674_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _01644_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _01647_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _01702_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _01706_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _01710_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _01714_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _01718_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _01722_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _01726_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _01696_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _01698_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _01754_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _01758_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _01762_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _01766_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _01770_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _01774_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _01777_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _01747_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _01750_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _01806_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _01810_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _01813_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _01817_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _01821_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _01825_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _01829_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _01799_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _01802_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _01857_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _01861_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _01865_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _01869_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _01873_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _01877_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _01881_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _01850_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _01853_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _40911_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _40912_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _40914_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _40915_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _40916_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _40917_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _40918_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40679_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _40899_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _40900_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _40902_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _40903_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _40904_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _40905_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _40906_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _40908_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _40887_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _40888_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _40890_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _40891_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _40892_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _40893_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _40894_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _40896_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40875_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40876_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40877_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40879_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40880_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40881_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40882_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40883_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40863_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40864_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40865_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40866_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40868_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40869_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40870_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40871_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40851_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40852_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40853_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40854_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40855_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40857_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40858_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40859_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40839_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40840_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40841_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40842_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40843_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40845_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40846_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40847_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40826_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40828_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40829_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40830_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40831_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40832_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40834_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40835_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40814_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40815_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40816_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40817_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40819_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40820_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40821_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40822_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40802_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40803_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40804_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40805_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40806_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40808_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40809_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40810_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40790_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40791_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40792_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40793_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40794_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40796_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40797_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40798_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40777_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40779_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40780_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40781_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40782_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40783_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40785_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40786_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40765_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40766_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40767_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40768_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40770_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40771_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40772_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40773_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40752_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40754_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40755_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40756_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40757_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40758_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40760_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40761_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40740_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40741_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40742_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40743_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40745_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40746_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40747_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40748_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40726_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40727_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40729_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40730_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40731_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40733_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40734_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40735_);
  dff (\oc8051_golden_model_1.B [0], _43376_);
  dff (\oc8051_golden_model_1.B [1], _43377_);
  dff (\oc8051_golden_model_1.B [2], _43378_);
  dff (\oc8051_golden_model_1.B [3], _43379_);
  dff (\oc8051_golden_model_1.B [4], _43380_);
  dff (\oc8051_golden_model_1.B [5], _43381_);
  dff (\oc8051_golden_model_1.B [6], _43382_);
  dff (\oc8051_golden_model_1.B [7], _40680_);
  dff (\oc8051_golden_model_1.ACC [0], _43383_);
  dff (\oc8051_golden_model_1.ACC [1], _43384_);
  dff (\oc8051_golden_model_1.ACC [2], _43385_);
  dff (\oc8051_golden_model_1.ACC [3], _43386_);
  dff (\oc8051_golden_model_1.ACC [4], _43387_);
  dff (\oc8051_golden_model_1.ACC [5], _43390_);
  dff (\oc8051_golden_model_1.ACC [6], _43391_);
  dff (\oc8051_golden_model_1.ACC [7], _40681_);
  dff (\oc8051_golden_model_1.SBUF [0], _43392_);
  dff (\oc8051_golden_model_1.SBUF [1], _43395_);
  dff (\oc8051_golden_model_1.SBUF [2], _43396_);
  dff (\oc8051_golden_model_1.SBUF [3], _43397_);
  dff (\oc8051_golden_model_1.SBUF [4], _43398_);
  dff (\oc8051_golden_model_1.SBUF [5], _43399_);
  dff (\oc8051_golden_model_1.SBUF [6], _43400_);
  dff (\oc8051_golden_model_1.SBUF [7], _40683_);
  dff (\oc8051_golden_model_1.SCON [0], _43401_);
  dff (\oc8051_golden_model_1.SCON [1], _43402_);
  dff (\oc8051_golden_model_1.SCON [2], _43403_);
  dff (\oc8051_golden_model_1.SCON [3], _43404_);
  dff (\oc8051_golden_model_1.SCON [4], _43405_);
  dff (\oc8051_golden_model_1.SCON [5], _43406_);
  dff (\oc8051_golden_model_1.SCON [6], _43407_);
  dff (\oc8051_golden_model_1.SCON [7], _40684_);
  dff (\oc8051_golden_model_1.PCON [0], _43410_);
  dff (\oc8051_golden_model_1.PCON [1], _43411_);
  dff (\oc8051_golden_model_1.PCON [2], _43412_);
  dff (\oc8051_golden_model_1.PCON [3], _43415_);
  dff (\oc8051_golden_model_1.PCON [4], _43416_);
  dff (\oc8051_golden_model_1.PCON [5], _43417_);
  dff (\oc8051_golden_model_1.PCON [6], _43418_);
  dff (\oc8051_golden_model_1.PCON [7], _40685_);
  dff (\oc8051_golden_model_1.TCON [0], _43419_);
  dff (\oc8051_golden_model_1.TCON [1], _43420_);
  dff (\oc8051_golden_model_1.TCON [2], _43421_);
  dff (\oc8051_golden_model_1.TCON [3], _43422_);
  dff (\oc8051_golden_model_1.TCON [4], _43423_);
  dff (\oc8051_golden_model_1.TCON [5], _43424_);
  dff (\oc8051_golden_model_1.TCON [6], _43425_);
  dff (\oc8051_golden_model_1.TCON [7], _40686_);
  dff (\oc8051_golden_model_1.TL0 [0], _43428_);
  dff (\oc8051_golden_model_1.TL0 [1], _43429_);
  dff (\oc8051_golden_model_1.TL0 [2], _43430_);
  dff (\oc8051_golden_model_1.TL0 [3], _43431_);
  dff (\oc8051_golden_model_1.TL0 [4], _43432_);
  dff (\oc8051_golden_model_1.TL0 [5], _43435_);
  dff (\oc8051_golden_model_1.TL0 [6], _43436_);
  dff (\oc8051_golden_model_1.TL0 [7], _40687_);
  dff (\oc8051_golden_model_1.TL1 [0], _43437_);
  dff (\oc8051_golden_model_1.TL1 [1], _43439_);
  dff (\oc8051_golden_model_1.TL1 [2], _43440_);
  dff (\oc8051_golden_model_1.TL1 [3], _43441_);
  dff (\oc8051_golden_model_1.TL1 [4], _43442_);
  dff (\oc8051_golden_model_1.TL1 [5], _43443_);
  dff (\oc8051_golden_model_1.TL1 [6], _43444_);
  dff (\oc8051_golden_model_1.TL1 [7], _40689_);
  dff (\oc8051_golden_model_1.TH0 [0], _43447_);
  dff (\oc8051_golden_model_1.TH0 [1], _43448_);
  dff (\oc8051_golden_model_1.TH0 [2], _43449_);
  dff (\oc8051_golden_model_1.TH0 [3], _43450_);
  dff (\oc8051_golden_model_1.TH0 [4], _43451_);
  dff (\oc8051_golden_model_1.TH0 [5], _43452_);
  dff (\oc8051_golden_model_1.TH0 [6], _43453_);
  dff (\oc8051_golden_model_1.TH0 [7], _40690_);
  dff (\oc8051_golden_model_1.TH1 [0], _43455_);
  dff (\oc8051_golden_model_1.TH1 [1], _43456_);
  dff (\oc8051_golden_model_1.TH1 [2], _43457_);
  dff (\oc8051_golden_model_1.TH1 [3], _43458_);
  dff (\oc8051_golden_model_1.TH1 [4], _43459_);
  dff (\oc8051_golden_model_1.TH1 [5], _43460_);
  dff (\oc8051_golden_model_1.TH1 [6], _43461_);
  dff (\oc8051_golden_model_1.TH1 [7], _40691_);
  dff (\oc8051_golden_model_1.TMOD [0], _43464_);
  dff (\oc8051_golden_model_1.TMOD [1], _43465_);
  dff (\oc8051_golden_model_1.TMOD [2], _43466_);
  dff (\oc8051_golden_model_1.TMOD [3], _43467_);
  dff (\oc8051_golden_model_1.TMOD [4], _43468_);
  dff (\oc8051_golden_model_1.TMOD [5], _43469_);
  dff (\oc8051_golden_model_1.TMOD [6], _43470_);
  dff (\oc8051_golden_model_1.TMOD [7], _40692_);
  dff (\oc8051_golden_model_1.IE [0], _43473_);
  dff (\oc8051_golden_model_1.IE [1], _43474_);
  dff (\oc8051_golden_model_1.IE [2], _43475_);
  dff (\oc8051_golden_model_1.IE [3], _43476_);
  dff (\oc8051_golden_model_1.IE [4], _43477_);
  dff (\oc8051_golden_model_1.IE [5], _43478_);
  dff (\oc8051_golden_model_1.IE [6], _43479_);
  dff (\oc8051_golden_model_1.IE [7], _40693_);
  dff (\oc8051_golden_model_1.IP [0], _43480_);
  dff (\oc8051_golden_model_1.IP [1], _43483_);
  dff (\oc8051_golden_model_1.IP [2], _43484_);
  dff (\oc8051_golden_model_1.IP [3], _43485_);
  dff (\oc8051_golden_model_1.IP [4], _43486_);
  dff (\oc8051_golden_model_1.IP [5], _43487_);
  dff (\oc8051_golden_model_1.IP [6], _43488_);
  dff (\oc8051_golden_model_1.IP [7], _40695_);
  dff (\oc8051_golden_model_1.DPL [0], _43491_);
  dff (\oc8051_golden_model_1.DPL [1], _43492_);
  dff (\oc8051_golden_model_1.DPL [2], _43493_);
  dff (\oc8051_golden_model_1.DPL [3], _43494_);
  dff (\oc8051_golden_model_1.DPL [4], _43495_);
  dff (\oc8051_golden_model_1.DPL [5], _43496_);
  dff (\oc8051_golden_model_1.DPL [6], _43497_);
  dff (\oc8051_golden_model_1.DPL [7], _40696_);
  dff (\oc8051_golden_model_1.DPH [0], _43498_);
  dff (\oc8051_golden_model_1.DPH [1], _43499_);
  dff (\oc8051_golden_model_1.DPH [2], _43500_);
  dff (\oc8051_golden_model_1.DPH [3], _43503_);
  dff (\oc8051_golden_model_1.DPH [4], _43504_);
  dff (\oc8051_golden_model_1.DPH [5], _43505_);
  dff (\oc8051_golden_model_1.DPH [6], _43506_);
  dff (\oc8051_golden_model_1.DPH [7], _40697_);
  dff (\oc8051_golden_model_1.PC [0], _43509_);
  dff (\oc8051_golden_model_1.PC [1], _43510_);
  dff (\oc8051_golden_model_1.PC [2], _43511_);
  dff (\oc8051_golden_model_1.PC [3], _43512_);
  dff (\oc8051_golden_model_1.PC [4], _43513_);
  dff (\oc8051_golden_model_1.PC [5], _43514_);
  dff (\oc8051_golden_model_1.PC [6], _43515_);
  dff (\oc8051_golden_model_1.PC [7], _43516_);
  dff (\oc8051_golden_model_1.PC [8], _43517_);
  dff (\oc8051_golden_model_1.PC [9], _43518_);
  dff (\oc8051_golden_model_1.PC [10], _43519_);
  dff (\oc8051_golden_model_1.PC [11], _43522_);
  dff (\oc8051_golden_model_1.PC [12], _43523_);
  dff (\oc8051_golden_model_1.PC [13], _43524_);
  dff (\oc8051_golden_model_1.PC [14], _43525_);
  dff (\oc8051_golden_model_1.PC [15], _40698_);
  dff (\oc8051_golden_model_1.P2 [0], _43528_);
  dff (\oc8051_golden_model_1.P2 [1], _43529_);
  dff (\oc8051_golden_model_1.P2 [2], _43530_);
  dff (\oc8051_golden_model_1.P2 [3], _43531_);
  dff (\oc8051_golden_model_1.P2 [4], _43532_);
  dff (\oc8051_golden_model_1.P2 [5], _43533_);
  dff (\oc8051_golden_model_1.P2 [6], _43534_);
  dff (\oc8051_golden_model_1.P2 [7], _40699_);
  dff (\oc8051_golden_model_1.P3 [0], _43535_);
  dff (\oc8051_golden_model_1.P3 [1], _43536_);
  dff (\oc8051_golden_model_1.P3 [2], _43537_);
  dff (\oc8051_golden_model_1.P3 [3], _43538_);
  dff (\oc8051_golden_model_1.P3 [4], _43539_);
  dff (\oc8051_golden_model_1.P3 [5], _43542_);
  dff (\oc8051_golden_model_1.P3 [6], _43543_);
  dff (\oc8051_golden_model_1.P3 [7], _40701_);
  dff (\oc8051_golden_model_1.P0 [0], _43544_);
  dff (\oc8051_golden_model_1.P0 [1], _43547_);
  dff (\oc8051_golden_model_1.P0 [2], _43548_);
  dff (\oc8051_golden_model_1.P0 [3], _43549_);
  dff (\oc8051_golden_model_1.P0 [4], _43550_);
  dff (\oc8051_golden_model_1.P0 [5], _43551_);
  dff (\oc8051_golden_model_1.P0 [6], _43552_);
  dff (\oc8051_golden_model_1.P0 [7], _40702_);
  dff (\oc8051_golden_model_1.P1 [0], _43553_);
  dff (\oc8051_golden_model_1.P1 [1], _43554_);
  dff (\oc8051_golden_model_1.P1 [2], _43555_);
  dff (\oc8051_golden_model_1.P1 [3], _43556_);
  dff (\oc8051_golden_model_1.P1 [4], _43557_);
  dff (\oc8051_golden_model_1.P1 [5], _43558_);
  dff (\oc8051_golden_model_1.P1 [6], _43559_);
  dff (\oc8051_golden_model_1.P1 [7], _40703_);
  dff (\oc8051_golden_model_1.SP [0], _43562_);
  dff (\oc8051_golden_model_1.SP [1], _43563_);
  dff (\oc8051_golden_model_1.SP [2], _43564_);
  dff (\oc8051_golden_model_1.SP [3], _43567_);
  dff (\oc8051_golden_model_1.SP [4], _43568_);
  dff (\oc8051_golden_model_1.SP [5], _43569_);
  dff (\oc8051_golden_model_1.SP [6], _43570_);
  dff (\oc8051_golden_model_1.SP [7], _40704_);
  dff (\oc8051_golden_model_1.PSW [0], _43571_);
  dff (\oc8051_golden_model_1.PSW [1], _43572_);
  dff (\oc8051_golden_model_1.PSW [2], _43573_);
  dff (\oc8051_golden_model_1.PSW [3], _43574_);
  dff (\oc8051_golden_model_1.PSW [4], _43575_);
  dff (\oc8051_golden_model_1.PSW [5], _43576_);
  dff (\oc8051_golden_model_1.PSW [6], _43577_);
  dff (\oc8051_golden_model_1.PSW [7], _40705_);
  dff (\oc8051_golden_model_1.P0INREG [0], _43580_);
  dff (\oc8051_golden_model_1.P0INREG [1], _43581_);
  dff (\oc8051_golden_model_1.P0INREG [2], _43582_);
  dff (\oc8051_golden_model_1.P0INREG [3], _43583_);
  dff (\oc8051_golden_model_1.P0INREG [4], _43584_);
  dff (\oc8051_golden_model_1.P0INREG [5], _43587_);
  dff (\oc8051_golden_model_1.P0INREG [6], _43588_);
  dff (\oc8051_golden_model_1.P0INREG [7], _40707_);
  dff (\oc8051_golden_model_1.P1INREG [0], _43589_);
  dff (\oc8051_golden_model_1.P1INREG [1], _43591_);
  dff (\oc8051_golden_model_1.P1INREG [2], _43592_);
  dff (\oc8051_golden_model_1.P1INREG [3], _43593_);
  dff (\oc8051_golden_model_1.P1INREG [4], _43594_);
  dff (\oc8051_golden_model_1.P1INREG [5], _43595_);
  dff (\oc8051_golden_model_1.P1INREG [6], _43596_);
  dff (\oc8051_golden_model_1.P1INREG [7], _40708_);
  dff (\oc8051_golden_model_1.P2INREG [0], _43599_);
  dff (\oc8051_golden_model_1.P2INREG [1], _43600_);
  dff (\oc8051_golden_model_1.P2INREG [2], _43601_);
  dff (\oc8051_golden_model_1.P2INREG [3], _43602_);
  dff (\oc8051_golden_model_1.P2INREG [4], _43603_);
  dff (\oc8051_golden_model_1.P2INREG [5], _43604_);
  dff (\oc8051_golden_model_1.P2INREG [6], _43605_);
  dff (\oc8051_golden_model_1.P2INREG [7], _40709_);
  dff (\oc8051_golden_model_1.P3INREG [0], _43607_);
  dff (\oc8051_golden_model_1.P3INREG [1], _43608_);
  dff (\oc8051_golden_model_1.P3INREG [2], _43609_);
  dff (\oc8051_golden_model_1.P3INREG [3], _43610_);
  dff (\oc8051_golden_model_1.P3INREG [4], _43611_);
  dff (\oc8051_golden_model_1.P3INREG [5], _43612_);
  dff (\oc8051_golden_model_1.P3INREG [6], _43613_);
  dff (\oc8051_golden_model_1.P3INREG [7], _40710_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02970_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02981_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03001_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03022_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03043_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00864_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03053_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00839_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03064_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03075_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03085_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03096_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03107_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03118_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03129_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00882_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02425_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22329_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02620_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02814_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03012_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03220_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03421_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03622_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03823_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04024_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04125_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04226_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04327_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04428_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04529_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04630_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04731_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24502_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38879_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38880_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38881_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38882_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38883_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38884_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38885_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38864_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38886_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38888_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38889_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38890_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38891_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38892_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38894_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38866_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38895_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38896_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38897_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38898_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38900_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38901_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38902_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38867_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _30379_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05963_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _30382_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05966_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _30384_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _30386_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05969_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _30388_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _30390_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05972_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _30392_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05975_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _30394_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _30396_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _30398_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _05978_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _30400_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05981_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _05984_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _06043_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _06045_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _05948_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _06048_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _06051_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _05951_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _06054_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _05954_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _06057_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _06060_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _06063_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _06066_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _06069_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _06072_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _06075_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _05957_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _05960_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39668_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _39701_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _39702_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _39703_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _39704_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _39705_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _39707_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _39708_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39669_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _39709_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _39710_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _39711_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _39712_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _39713_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _39714_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _39715_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39670_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _39716_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _39718_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _39719_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _39720_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _39721_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _39722_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _39723_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39672_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _39724_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _39725_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _39726_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _39727_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _39729_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _39730_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _39731_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39673_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39245_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39246_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39247_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39248_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38961_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39034_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39035_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39036_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39038_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39039_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39040_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39041_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39042_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39043_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39044_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39045_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39046_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39047_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39049_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39050_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38923_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39054_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39057_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39059_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39060_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39061_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39063_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39064_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39065_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39066_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39068_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39069_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38924_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39249_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39250_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39252_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39253_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39254_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39255_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39256_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39257_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39258_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39259_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39260_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39261_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39263_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39264_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39265_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39266_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39267_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39268_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39269_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39270_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39271_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39272_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39274_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39275_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39276_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39277_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39278_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39279_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39280_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39281_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39282_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38986_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38959_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39284_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39285_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39286_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39287_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39288_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39290_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39291_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39292_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39293_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39294_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39295_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39296_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39297_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39298_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38964_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39300_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39301_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39302_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39303_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39304_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39305_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39306_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38966_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38967_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39307_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39308_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39309_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39311_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39312_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39313_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39314_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38968_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39315_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39316_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39317_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39318_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39319_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39320_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39322_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39323_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39324_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39325_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39326_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39327_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39328_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39329_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39330_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38970_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39331_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39333_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39334_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39335_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39336_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39337_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39338_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39339_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39340_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39341_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39342_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39343_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39344_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39345_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39346_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38971_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38972_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38975_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38973_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39347_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39348_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39349_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39350_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39351_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39352_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39354_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38976_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38977_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39358_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39359_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39360_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39361_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39362_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39363_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38978_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39365_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39366_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39367_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39368_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39369_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39370_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39371_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38979_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _38980_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39372_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39373_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39374_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39376_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39377_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39378_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39379_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38982_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _38983_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38984_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39381_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39382_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38985_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39383_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39384_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39385_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39387_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39388_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39389_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39390_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39391_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39392_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39393_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39394_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39395_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39396_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39398_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39399_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39400_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39401_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39402_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39403_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39404_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39405_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39406_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39407_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39410_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39411_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39412_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39413_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39414_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39415_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39416_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38987_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39417_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39418_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39420_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39421_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39422_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39423_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39424_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38989_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38990_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38991_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39425_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39426_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39427_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39428_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39429_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39431_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39432_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39433_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39434_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39436_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39437_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39438_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39439_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39440_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38992_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38993_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38994_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38995_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39442_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39443_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39444_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39446_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39448_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39449_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39450_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39451_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39453_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39454_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39455_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39456_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39457_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38996_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38997_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39876_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39895_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39896_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39897_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39899_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39900_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39901_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39902_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39878_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39879_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39903_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39904_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _43906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _43910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _43914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _43918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _43922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _43926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _43930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _42959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _43874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _43878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _43882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _43886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _43890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _43894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _43898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _43901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _43842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _43846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _43850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _43854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _43858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _43862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _43866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _43869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _43214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _43220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _43226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _43232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _43238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _43244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _43250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _43253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _43261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _43265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _43269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _43273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _43277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _43279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _43282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _43285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _43293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _43297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _43301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _43305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _43309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _43313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _43317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _43320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _43361_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _43365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _43369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _43373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _43389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _43409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _43427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _43438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _43326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _43330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _43334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _43338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _43342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _43346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _43350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _43353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _43713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _43717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _43721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _43725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _43729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _43733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _43737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _43740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _43682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _43686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _43689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _43693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _43697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _43701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _43705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _43708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _43647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _43651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _43655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _43659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _43663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _43667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _43671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _43674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _43615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _43619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _43623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _43627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _43631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _43635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _43639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _43642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _43463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _43482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _43502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _43521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _43541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _43561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _43579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _43590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _43745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _43749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _43753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _43757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _43761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _43765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _43769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _43772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _43810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _43814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _43818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _43822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _43826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _43830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _43834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _43837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _43777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _43781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _43785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _43789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _43793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _43797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _43801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _43804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _01362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _01364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _01366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _01368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _01370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _01372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _01374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _42947_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39761_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39762_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39825_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39826_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39828_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39829_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39830_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39831_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39832_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39763_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24110_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22208_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08885_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08896_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08907_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08918_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13577_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13625_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13674_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12675_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _41894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _42811_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _42813_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _42817_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _42818_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _42820_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41892_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _42824_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _41890_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _41888_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _42826_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _42827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _41886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _42829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _42831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _41885_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _42833_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _42835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _41849_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _41847_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _41845_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _41844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _42837_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _42839_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _42841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _41841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _42843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _42844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _42846_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _42848_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _42850_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _42852_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _42854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _41839_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _42856_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _42858_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _42860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _42862_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _42864_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _42866_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _42868_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _41836_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35386_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41310_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41312_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41319_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41321_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41333_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35432_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41335_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41338_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41340_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35455_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21381_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21392_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21404_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21438_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16447_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09495_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10663_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10674_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10685_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09516_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [0], \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [1], \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [2], \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [3], \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [4], \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [5], \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [6], \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [7], \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [0], \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [1], \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [2], \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [3], \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [4], \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [5], \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [6], \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [7], \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [0], \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [1], \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [2], \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [3], \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [4], \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [5], \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [6], \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [7], \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [0], \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [1], \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [2], \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [3], \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [4], \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [5], \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [6], \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [7], \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1283 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1300 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1439 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1439 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1489 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1475 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1489 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1489 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1569 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1605 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1605 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1638 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1638 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1671 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1671 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1732 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1732 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1732 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1732 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1732 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1732 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1732 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1789 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1806 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1823 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1823 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1866 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1866 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1866 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1866 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1866 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1866 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1866 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1923 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1940 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1957 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1957 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2074 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2091 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2108 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2108 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2132 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2148 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2190 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2148 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2216 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2216 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2148 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2457 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2457 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2457 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2457 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2487 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2487 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2487 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2487 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2517 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2517 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2552 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2555 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2583 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2583 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2589 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2629 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2682 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2735 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2735 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2823 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2823 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2845 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2845 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2864 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2735 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2881 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.n2882 [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.n2882 [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.n2882 [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.n2882 [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.n2882 [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.n2882 [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.n2882 [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0988 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n0988 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n0988 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0988 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0988 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n0988 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n0988 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0989 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0990 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0991 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0992 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0993 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0995 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0996 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1003 , \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1011 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1011 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1011 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1011 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1011 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1011 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1011 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1017 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1018 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1019 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1026 , \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.n1027 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1027 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1027 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1027 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1027 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1043 , \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.n1044 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1044 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1044 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1044 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1044 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1044 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1044 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1156 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1156 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1156 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1156 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1158 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1158 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1158 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1158 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1160 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1160 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1160 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1160 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1161 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1161 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1162 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1163 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1164 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1165 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1165 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1166 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1213 , \oc8051_golden_model_1.n2555 [7]);
  buf(\oc8051_golden_model_1.n1258 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1259 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1259 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1259 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1259 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1259 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1259 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1259 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1259 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1259 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1260 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1261 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1261 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1261 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1261 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1261 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1262 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1263 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1263 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1263 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1264 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1265 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1265 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1266 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1266 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1266 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1266 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1266 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1266 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1266 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1267 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1267 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1267 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1267 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1267 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1267 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1268 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1269 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1270 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1271 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1272 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1273 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1274 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1282 , \oc8051_golden_model_1.n1283 [0]);
  buf(\oc8051_golden_model_1.n1283 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1283 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1283 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1283 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1283 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1283 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1283 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1299 , \oc8051_golden_model_1.n1300 [0]);
  buf(\oc8051_golden_model_1.n1300 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1300 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1300 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1300 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1300 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1300 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1300 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1343 [9], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1343 [10], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1343 [11], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1343 [12], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.n1343 [13], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.n1343 [14], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.n1343 [15], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n1345 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1345 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1345 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1345 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1345 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1345 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1345 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1345 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1346 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1352 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1360 , \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.n1361 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1361 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1361 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1361 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1361 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1361 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1361 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1363 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1363 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1363 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1363 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1363 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1363 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1363 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1363 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1363 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1367 [8], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1368 , \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1369 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1369 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1370 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1370 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1370 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1374 [4], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1375 , \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1376 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1376 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1376 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1376 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1376 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1384 , \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1385 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1385 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1385 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1385 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1385 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1385 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1386 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1386 [1], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1386 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1386 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1386 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1386 [5], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1386 [6], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1401 , \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.n1402 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1402 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1402 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1402 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1406 [8], \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.n1407 , \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.n1412 [4], \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.n1413 , \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.n1421 , \oc8051_golden_model_1.n1439 [2]);
  buf(\oc8051_golden_model_1.n1422 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1422 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1422 [2], \oc8051_golden_model_1.n1439 [2]);
  buf(\oc8051_golden_model_1.n1422 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1422 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1422 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1422 [6], \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.n1422 [7], \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.n1423 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1423 [1], \oc8051_golden_model_1.n1439 [2]);
  buf(\oc8051_golden_model_1.n1423 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1423 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1423 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1423 [5], \oc8051_golden_model_1.n1439 [6]);
  buf(\oc8051_golden_model_1.n1423 [6], \oc8051_golden_model_1.n1439 [7]);
  buf(\oc8051_golden_model_1.n1438 , \oc8051_golden_model_1.n1439 [0]);
  buf(\oc8051_golden_model_1.n1439 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1439 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1439 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1439 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1441 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1441 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1441 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1441 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1441 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n1441 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n1441 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n1441 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n1441 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1443 [8], \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.n1444 , \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.n1445 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1445 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1445 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1445 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1446 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1446 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1446 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1446 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1446 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1448 [4], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1449 , \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1450 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n1450 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n1450 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n1450 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n1450 [4], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n1450 [5], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n1450 [6], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n1450 [7], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n1450 [8], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n1457 , \oc8051_golden_model_1.n1475 [2]);
  buf(\oc8051_golden_model_1.n1458 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1458 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1458 [2], \oc8051_golden_model_1.n1475 [2]);
  buf(\oc8051_golden_model_1.n1458 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1458 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1458 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1458 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1458 [7], \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.n1459 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1459 [1], \oc8051_golden_model_1.n1475 [2]);
  buf(\oc8051_golden_model_1.n1459 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1459 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1459 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1459 [5], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1459 [6], \oc8051_golden_model_1.n1475 [7]);
  buf(\oc8051_golden_model_1.n1474 , \oc8051_golden_model_1.n1489 [0]);
  buf(\oc8051_golden_model_1.n1475 [0], \oc8051_golden_model_1.n1489 [0]);
  buf(\oc8051_golden_model_1.n1475 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1475 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1475 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1475 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1475 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1478 [8], \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.n1479 , \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.n1486 , \oc8051_golden_model_1.n1489 [2]);
  buf(\oc8051_golden_model_1.n1487 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1487 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1487 [2], \oc8051_golden_model_1.n1489 [2]);
  buf(\oc8051_golden_model_1.n1487 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1487 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1487 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1487 [6], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1487 [7], \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.n1488 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1488 [1], \oc8051_golden_model_1.n1489 [2]);
  buf(\oc8051_golden_model_1.n1488 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1488 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1488 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1488 [5], \oc8051_golden_model_1.n1489 [6]);
  buf(\oc8051_golden_model_1.n1488 [6], \oc8051_golden_model_1.n1489 [7]);
  buf(\oc8051_golden_model_1.n1489 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1489 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1489 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1489 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1491 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1491 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1491 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1491 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1491 [4], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.n1491 [5], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.n1491 [6], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.n1491 [7], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n1491 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1493 [8], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1494 , \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1495 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1495 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1495 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1495 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1495 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1497 [4], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1498 , \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1499 [0], \oc8051_golden_model_1.n2743 );
  buf(\oc8051_golden_model_1.n1499 [1], \oc8051_golden_model_1.n2742 );
  buf(\oc8051_golden_model_1.n1499 [2], \oc8051_golden_model_1.n2741 );
  buf(\oc8051_golden_model_1.n1499 [3], \oc8051_golden_model_1.n2740 );
  buf(\oc8051_golden_model_1.n1499 [4], \oc8051_golden_model_1.n2739 );
  buf(\oc8051_golden_model_1.n1499 [5], \oc8051_golden_model_1.n2738 );
  buf(\oc8051_golden_model_1.n1499 [6], \oc8051_golden_model_1.n2737 );
  buf(\oc8051_golden_model_1.n1499 [7], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n1499 [8], \oc8051_golden_model_1.n2736 );
  buf(\oc8051_golden_model_1.n1506 , \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1507 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1507 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1507 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1507 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1508 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1508 [1], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1508 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1508 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1508 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1508 [5], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1508 [6], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1523 , \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.n1524 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.n1524 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1524 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1524 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1524 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1524 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1524 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1524 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1527 , \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1528 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1528 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1528 [2], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1528 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1528 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1528 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1528 [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1528 [7], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1529 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1529 [1], \oc8051_golden_model_1.n1530 [2]);
  buf(\oc8051_golden_model_1.n1529 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1529 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1529 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1529 [5], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1529 [6], \oc8051_golden_model_1.n1530 [7]);
  buf(\oc8051_golden_model_1.n1530 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.n1530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1530 [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1532 [8], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1533 , \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1540 , \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1541 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1541 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1541 [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1541 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1541 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1541 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1541 [6], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1541 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.n1543 [6]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1543 [0], \oc8051_golden_model_1.n1546 [0]);
  buf(\oc8051_golden_model_1.n1543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1543 [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1543 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1544 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1544 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1544 [2], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1544 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1544 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1544 [6], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1544 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1545 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1545 [1], \oc8051_golden_model_1.n1546 [2]);
  buf(\oc8051_golden_model_1.n1545 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1545 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1545 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1545 [5], \oc8051_golden_model_1.n1546 [6]);
  buf(\oc8051_golden_model_1.n1545 [6], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1549 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1549 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1549 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1549 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1549 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1549 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1549 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1549 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1549 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1550 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1550 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1550 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1550 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1550 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1550 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1550 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1550 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1550 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1551 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1551 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1551 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1551 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1551 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1551 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1551 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1551 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1552 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1552 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1552 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1552 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1552 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1552 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1552 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1552 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1553 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1553 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1553 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1553 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1553 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1553 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1553 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1555 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1557 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1559 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1560 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1561 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 , \oc8051_golden_model_1.n1569 [0]);
  buf(\oc8051_golden_model_1.n1569 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1569 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1569 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1569 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1569 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1569 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1569 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1570 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1570 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1573 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [8], \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.n1576 , \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.n1577 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1577 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1579 [4], \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.n1580 , \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.n1587 , \oc8051_golden_model_1.n1605 [2]);
  buf(\oc8051_golden_model_1.n1588 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1588 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1588 [2], \oc8051_golden_model_1.n1605 [2]);
  buf(\oc8051_golden_model_1.n1588 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1588 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1588 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1588 [6], \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.n1588 [7], \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.n1589 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1589 [1], \oc8051_golden_model_1.n1605 [2]);
  buf(\oc8051_golden_model_1.n1589 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1589 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1589 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1589 [5], \oc8051_golden_model_1.n1605 [6]);
  buf(\oc8051_golden_model_1.n1589 [6], \oc8051_golden_model_1.n1605 [7]);
  buf(\oc8051_golden_model_1.n1604 , \oc8051_golden_model_1.n1605 [0]);
  buf(\oc8051_golden_model_1.n1605 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1605 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1605 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1605 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1609 [8], \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.n1610 , \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.n1612 [4], \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.n1613 , \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.n1620 , \oc8051_golden_model_1.n1638 [2]);
  buf(\oc8051_golden_model_1.n1621 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1621 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1621 [2], \oc8051_golden_model_1.n1638 [2]);
  buf(\oc8051_golden_model_1.n1621 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1621 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1621 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1621 [6], \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.n1621 [7], \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.n1622 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1622 [1], \oc8051_golden_model_1.n1638 [2]);
  buf(\oc8051_golden_model_1.n1622 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1622 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1622 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1622 [5], \oc8051_golden_model_1.n1638 [6]);
  buf(\oc8051_golden_model_1.n1622 [6], \oc8051_golden_model_1.n1638 [7]);
  buf(\oc8051_golden_model_1.n1637 , \oc8051_golden_model_1.n1638 [0]);
  buf(\oc8051_golden_model_1.n1638 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1638 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1638 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1638 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1642 [8], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.n1643 , \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.n1645 [4], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.n1646 , \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.n1653 , \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.n1654 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1654 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1654 [2], \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.n1654 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1654 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1654 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1654 [6], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.n1654 [7], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.n1655 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1655 [1], \oc8051_golden_model_1.n1671 [2]);
  buf(\oc8051_golden_model_1.n1655 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1655 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1655 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1655 [5], \oc8051_golden_model_1.n1671 [6]);
  buf(\oc8051_golden_model_1.n1655 [6], \oc8051_golden_model_1.n1671 [7]);
  buf(\oc8051_golden_model_1.n1670 , \oc8051_golden_model_1.n1671 [0]);
  buf(\oc8051_golden_model_1.n1671 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1671 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1671 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1671 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1675 [8], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.n1676 , \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.n1678 [4], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.n1679 , \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.n1686 , \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.n1687 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1687 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1687 [2], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.n1687 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1687 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1687 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1687 [6], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.n1687 [7], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.n1688 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1688 [1], \oc8051_golden_model_1.n1704 [2]);
  buf(\oc8051_golden_model_1.n1688 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1688 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1688 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1688 [5], \oc8051_golden_model_1.n1704 [6]);
  buf(\oc8051_golden_model_1.n1688 [6], \oc8051_golden_model_1.n1704 [7]);
  buf(\oc8051_golden_model_1.n1703 , \oc8051_golden_model_1.n1704 [0]);
  buf(\oc8051_golden_model_1.n1704 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1704 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1704 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1704 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1730 [1], \oc8051_golden_model_1.n1732 [1]);
  buf(\oc8051_golden_model_1.n1730 [2], \oc8051_golden_model_1.n1732 [2]);
  buf(\oc8051_golden_model_1.n1730 [3], \oc8051_golden_model_1.n1732 [3]);
  buf(\oc8051_golden_model_1.n1730 [4], \oc8051_golden_model_1.n1732 [4]);
  buf(\oc8051_golden_model_1.n1730 [5], \oc8051_golden_model_1.n1732 [5]);
  buf(\oc8051_golden_model_1.n1730 [6], \oc8051_golden_model_1.n1732 [6]);
  buf(\oc8051_golden_model_1.n1730 [7], \oc8051_golden_model_1.n1732 [7]);
  buf(\oc8051_golden_model_1.n1731 [0], \oc8051_golden_model_1.n1732 [1]);
  buf(\oc8051_golden_model_1.n1731 [1], \oc8051_golden_model_1.n1732 [2]);
  buf(\oc8051_golden_model_1.n1731 [2], \oc8051_golden_model_1.n1732 [3]);
  buf(\oc8051_golden_model_1.n1731 [3], \oc8051_golden_model_1.n1732 [4]);
  buf(\oc8051_golden_model_1.n1731 [4], \oc8051_golden_model_1.n1732 [5]);
  buf(\oc8051_golden_model_1.n1731 [5], \oc8051_golden_model_1.n1732 [6]);
  buf(\oc8051_golden_model_1.n1731 [6], \oc8051_golden_model_1.n1732 [7]);
  buf(\oc8051_golden_model_1.n1732 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n1788 , \oc8051_golden_model_1.n1789 [0]);
  buf(\oc8051_golden_model_1.n1789 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1789 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1789 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1789 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1789 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1789 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1789 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1805 , \oc8051_golden_model_1.n1806 [0]);
  buf(\oc8051_golden_model_1.n1806 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1806 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1806 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1806 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1806 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1806 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1806 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1822 , \oc8051_golden_model_1.n1823 [0]);
  buf(\oc8051_golden_model_1.n1823 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1823 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1823 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1823 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1823 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1823 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1823 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1839 , \oc8051_golden_model_1.n1840 [0]);
  buf(\oc8051_golden_model_1.n1840 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1840 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1840 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1840 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1840 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1840 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1840 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1864 [1], \oc8051_golden_model_1.n1866 [1]);
  buf(\oc8051_golden_model_1.n1864 [2], \oc8051_golden_model_1.n1866 [2]);
  buf(\oc8051_golden_model_1.n1864 [3], \oc8051_golden_model_1.n1866 [3]);
  buf(\oc8051_golden_model_1.n1864 [4], \oc8051_golden_model_1.n1866 [4]);
  buf(\oc8051_golden_model_1.n1864 [5], \oc8051_golden_model_1.n1866 [5]);
  buf(\oc8051_golden_model_1.n1864 [6], \oc8051_golden_model_1.n1866 [6]);
  buf(\oc8051_golden_model_1.n1864 [7], \oc8051_golden_model_1.n1866 [7]);
  buf(\oc8051_golden_model_1.n1865 [0], \oc8051_golden_model_1.n1866 [1]);
  buf(\oc8051_golden_model_1.n1865 [1], \oc8051_golden_model_1.n1866 [2]);
  buf(\oc8051_golden_model_1.n1865 [2], \oc8051_golden_model_1.n1866 [3]);
  buf(\oc8051_golden_model_1.n1865 [3], \oc8051_golden_model_1.n1866 [4]);
  buf(\oc8051_golden_model_1.n1865 [4], \oc8051_golden_model_1.n1866 [5]);
  buf(\oc8051_golden_model_1.n1865 [5], \oc8051_golden_model_1.n1866 [6]);
  buf(\oc8051_golden_model_1.n1865 [6], \oc8051_golden_model_1.n1866 [7]);
  buf(\oc8051_golden_model_1.n1866 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n1922 , \oc8051_golden_model_1.n1923 [0]);
  buf(\oc8051_golden_model_1.n1923 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1923 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1923 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1923 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1923 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1923 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1923 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1939 , \oc8051_golden_model_1.n1940 [0]);
  buf(\oc8051_golden_model_1.n1940 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1940 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1940 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1940 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1940 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1940 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1940 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1956 , \oc8051_golden_model_1.n1957 [0]);
  buf(\oc8051_golden_model_1.n1957 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1957 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1957 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1957 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1957 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1957 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1957 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1973 , \oc8051_golden_model_1.n1974 [0]);
  buf(\oc8051_golden_model_1.n1974 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1974 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1974 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1974 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1974 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1974 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1974 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2073 , \oc8051_golden_model_1.n2074 [0]);
  buf(\oc8051_golden_model_1.n2074 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2074 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2074 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2074 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2074 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2074 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2074 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2090 , \oc8051_golden_model_1.n2091 [0]);
  buf(\oc8051_golden_model_1.n2091 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2091 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2091 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2091 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2091 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2091 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2091 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2107 , \oc8051_golden_model_1.n2108 [0]);
  buf(\oc8051_golden_model_1.n2108 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2108 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2108 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2108 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2108 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2108 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2108 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2124 , \oc8051_golden_model_1.n2125 [0]);
  buf(\oc8051_golden_model_1.n2125 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2125 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2125 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2125 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2125 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2125 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2125 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2128 , \oc8051_golden_model_1.n2132 [7]);
  buf(\oc8051_golden_model_1.n2129 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2129 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2129 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2129 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2129 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2129 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2129 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2130 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2130 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2130 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2130 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2130 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2130 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2130 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2130 [7], \oc8051_golden_model_1.n2132 [7]);
  buf(\oc8051_golden_model_1.n2131 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2131 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2131 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2131 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2131 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2131 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2131 [6], \oc8051_golden_model_1.n2132 [7]);
  buf(\oc8051_golden_model_1.n2132 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2132 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2132 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2132 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2132 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2132 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2132 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2147 , \oc8051_golden_model_1.n2148 [0]);
  buf(\oc8051_golden_model_1.n2148 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2148 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2148 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2148 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2148 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2148 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2148 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2187 , \oc8051_golden_model_1.n2190 [7]);
  buf(\oc8051_golden_model_1.n2188 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2188 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2188 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2188 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2188 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2188 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2188 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2188 [7], \oc8051_golden_model_1.n2190 [7]);
  buf(\oc8051_golden_model_1.n2189 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2189 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2189 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2189 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2189 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2189 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2189 [6], \oc8051_golden_model_1.n2190 [7]);
  buf(\oc8051_golden_model_1.n2190 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2190 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2190 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2190 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2190 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2190 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2190 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2197 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2197 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2197 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2197 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2198 , \oc8051_golden_model_1.n2216 [2]);
  buf(\oc8051_golden_model_1.n2199 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2199 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2199 [2], \oc8051_golden_model_1.n2216 [2]);
  buf(\oc8051_golden_model_1.n2199 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2199 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2199 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2199 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2199 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2200 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2200 [1], \oc8051_golden_model_1.n2216 [2]);
  buf(\oc8051_golden_model_1.n2200 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2200 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2200 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2200 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2200 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2215 , \oc8051_golden_model_1.n2216 [0]);
  buf(\oc8051_golden_model_1.n2216 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2216 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2216 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2216 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2216 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2216 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2428 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2428 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2431 , \oc8051_golden_model_1.n2457 [7]);
  buf(\oc8051_golden_model_1.n2433 , \oc8051_golden_model_1.n2457 [6]);
  buf(\oc8051_golden_model_1.n2439 , \oc8051_golden_model_1.n2457 [2]);
  buf(\oc8051_golden_model_1.n2440 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2440 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2440 [2], \oc8051_golden_model_1.n2457 [2]);
  buf(\oc8051_golden_model_1.n2440 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2440 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2440 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2440 [6], \oc8051_golden_model_1.n2457 [6]);
  buf(\oc8051_golden_model_1.n2440 [7], \oc8051_golden_model_1.n2457 [7]);
  buf(\oc8051_golden_model_1.n2441 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2441 [1], \oc8051_golden_model_1.n2457 [2]);
  buf(\oc8051_golden_model_1.n2441 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2441 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2441 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2441 [5], \oc8051_golden_model_1.n2457 [6]);
  buf(\oc8051_golden_model_1.n2441 [6], \oc8051_golden_model_1.n2457 [7]);
  buf(\oc8051_golden_model_1.n2456 , \oc8051_golden_model_1.n2457 [0]);
  buf(\oc8051_golden_model_1.n2457 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2457 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2457 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2457 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2461 , \oc8051_golden_model_1.n2487 [7]);
  buf(\oc8051_golden_model_1.n2463 , \oc8051_golden_model_1.n2487 [6]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2487 [2]);
  buf(\oc8051_golden_model_1.n2470 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [2], \oc8051_golden_model_1.n2487 [2]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2470 [6], \oc8051_golden_model_1.n2487 [6]);
  buf(\oc8051_golden_model_1.n2470 [7], \oc8051_golden_model_1.n2487 [7]);
  buf(\oc8051_golden_model_1.n2471 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2471 [1], \oc8051_golden_model_1.n2487 [2]);
  buf(\oc8051_golden_model_1.n2471 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2471 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2471 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2471 [5], \oc8051_golden_model_1.n2487 [6]);
  buf(\oc8051_golden_model_1.n2471 [6], \oc8051_golden_model_1.n2487 [7]);
  buf(\oc8051_golden_model_1.n2486 , \oc8051_golden_model_1.n2487 [0]);
  buf(\oc8051_golden_model_1.n2487 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2487 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2487 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2487 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2491 , \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2493 , \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.n2499 , \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.n2500 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [2], \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2500 [6], \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.n2500 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2501 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2501 [1], \oc8051_golden_model_1.n2517 [2]);
  buf(\oc8051_golden_model_1.n2501 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2501 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2501 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2501 [5], \oc8051_golden_model_1.n2517 [6]);
  buf(\oc8051_golden_model_1.n2501 [6], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2516 , \oc8051_golden_model_1.n2517 [0]);
  buf(\oc8051_golden_model_1.n2517 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2517 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2517 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2517 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2521 , \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.n2523 , \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.n2530 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2530 [2], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.n2530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2530 [6], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.n2530 [7], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.n2531 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2531 [1], \oc8051_golden_model_1.n2547 [2]);
  buf(\oc8051_golden_model_1.n2531 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2531 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2531 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2531 [5], \oc8051_golden_model_1.n2547 [6]);
  buf(\oc8051_golden_model_1.n2531 [6], \oc8051_golden_model_1.n2547 [7]);
  buf(\oc8051_golden_model_1.n2546 , \oc8051_golden_model_1.n2547 [0]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2549 , \oc8051_golden_model_1.n2552 [7]);
  buf(\oc8051_golden_model_1.n2550 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2550 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2550 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2550 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2550 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2550 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2550 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2550 [7], \oc8051_golden_model_1.n2552 [7]);
  buf(\oc8051_golden_model_1.n2551 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2551 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2551 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2551 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2551 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2551 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2551 [6], \oc8051_golden_model_1.n2552 [7]);
  buf(\oc8051_golden_model_1.n2552 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2552 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2552 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2552 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2552 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2552 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2552 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2553 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2553 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2553 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2553 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2553 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2553 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2553 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2553 [7], \oc8051_golden_model_1.n2555 [7]);
  buf(\oc8051_golden_model_1.n2554 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2554 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2554 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2554 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2554 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2554 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2554 [6], \oc8051_golden_model_1.n2555 [7]);
  buf(\oc8051_golden_model_1.n2555 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2555 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2555 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2555 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2555 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2555 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2555 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2559 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2559 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2559 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2559 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2559 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2559 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2559 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2559 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2559 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2559 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2565 , \oc8051_golden_model_1.n2583 [2]);
  buf(\oc8051_golden_model_1.n2566 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.n2583 [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2567 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2567 [1], \oc8051_golden_model_1.n2583 [2]);
  buf(\oc8051_golden_model_1.n2567 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2567 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2567 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2567 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2567 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2582 , \oc8051_golden_model_1.n2583 [0]);
  buf(\oc8051_golden_model_1.n2583 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2583 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2583 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2583 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2583 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2583 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2586 , \oc8051_golden_model_1.n2589 [7]);
  buf(\oc8051_golden_model_1.n2587 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2587 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2587 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2587 [7], \oc8051_golden_model_1.n2589 [7]);
  buf(\oc8051_golden_model_1.n2588 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2588 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2588 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2588 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2588 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2588 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2588 [6], \oc8051_golden_model_1.n2589 [7]);
  buf(\oc8051_golden_model_1.n2589 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2589 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2589 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2589 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2589 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2589 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2589 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2626 , \oc8051_golden_model_1.n2629 [7]);
  buf(\oc8051_golden_model_1.n2627 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2627 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2627 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2627 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2627 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2627 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2627 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2627 [7], \oc8051_golden_model_1.n2629 [7]);
  buf(\oc8051_golden_model_1.n2628 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2628 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2628 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2628 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2628 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2628 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2628 [6], \oc8051_golden_model_1.n2629 [7]);
  buf(\oc8051_golden_model_1.n2629 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2629 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2629 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2629 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2629 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2629 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2629 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2634 , \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2635 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2635 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2635 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2635 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2635 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2635 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2635 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2635 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2636 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2636 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2636 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2636 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2636 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2636 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2636 [6], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2637 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2637 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2637 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2637 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2637 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2637 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2637 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2642 , \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2643 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2643 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2643 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2643 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2643 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2643 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2643 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2644 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2644 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2644 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2644 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2644 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2644 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2644 [6], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2645 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2645 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2645 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2645 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2645 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2645 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2645 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2650 , \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2651 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2651 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2651 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2651 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2651 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2651 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2651 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2651 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2658 , \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2659 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2659 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2659 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2659 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2659 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2659 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2659 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2659 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2660 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2660 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2660 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2660 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2660 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2660 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2660 [6], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2661 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2661 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2661 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2661 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2661 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2661 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2661 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2662 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2662 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2662 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2662 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2662 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2662 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2662 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2662 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2663 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2663 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2663 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2663 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2663 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2663 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2663 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2664 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2664 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2664 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2664 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2664 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2664 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2664 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2664 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2665 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2665 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2665 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2665 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2666 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2666 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2666 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2666 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2666 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2666 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2666 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2666 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2667 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2668 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2669 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2670 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2671 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2672 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2673 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2674 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2681 , \oc8051_golden_model_1.n2682 [0]);
  buf(\oc8051_golden_model_1.n2682 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2682 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2682 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2682 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2682 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2682 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2682 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2702 [1], \oc8051_golden_model_1.n2882 [1]);
  buf(\oc8051_golden_model_1.n2702 [2], \oc8051_golden_model_1.n2882 [2]);
  buf(\oc8051_golden_model_1.n2702 [3], \oc8051_golden_model_1.n2882 [3]);
  buf(\oc8051_golden_model_1.n2702 [4], \oc8051_golden_model_1.n2882 [4]);
  buf(\oc8051_golden_model_1.n2702 [5], \oc8051_golden_model_1.n2882 [5]);
  buf(\oc8051_golden_model_1.n2702 [6], \oc8051_golden_model_1.n2882 [6]);
  buf(\oc8051_golden_model_1.n2702 [7], \oc8051_golden_model_1.n2882 [7]);
  buf(\oc8051_golden_model_1.n2703 [0], \oc8051_golden_model_1.n2882 [1]);
  buf(\oc8051_golden_model_1.n2703 [1], \oc8051_golden_model_1.n2882 [2]);
  buf(\oc8051_golden_model_1.n2703 [2], \oc8051_golden_model_1.n2882 [3]);
  buf(\oc8051_golden_model_1.n2703 [3], \oc8051_golden_model_1.n2882 [4]);
  buf(\oc8051_golden_model_1.n2703 [4], \oc8051_golden_model_1.n2882 [5]);
  buf(\oc8051_golden_model_1.n2703 [5], \oc8051_golden_model_1.n2882 [6]);
  buf(\oc8051_golden_model_1.n2703 [6], \oc8051_golden_model_1.n2882 [7]);
  buf(\oc8051_golden_model_1.n2719 [1], \oc8051_golden_model_1.n2882 [1]);
  buf(\oc8051_golden_model_1.n2719 [2], \oc8051_golden_model_1.n2882 [2]);
  buf(\oc8051_golden_model_1.n2719 [3], \oc8051_golden_model_1.n2882 [3]);
  buf(\oc8051_golden_model_1.n2719 [4], \oc8051_golden_model_1.n2882 [4]);
  buf(\oc8051_golden_model_1.n2719 [5], \oc8051_golden_model_1.n2882 [5]);
  buf(\oc8051_golden_model_1.n2719 [6], \oc8051_golden_model_1.n2882 [6]);
  buf(\oc8051_golden_model_1.n2719 [7], \oc8051_golden_model_1.n2882 [7]);
  buf(\oc8051_golden_model_1.n2720 , \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n2721 , \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n2722 , \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n2723 , \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n2724 , \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n2725 , \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n2726 , \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n2727 , \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n2734 , \oc8051_golden_model_1.n2735 [0]);
  buf(\oc8051_golden_model_1.n2735 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2735 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2735 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2735 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2735 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2735 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2735 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2750 , \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2751 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2751 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2751 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2751 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2751 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2751 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2751 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2784 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2784 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2784 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2784 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2784 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2784 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2784 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2784 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2785 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2785 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2785 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2785 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2785 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2785 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2785 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2786 [0], \oc8051_golden_model_1.n2882 [0]);
  buf(\oc8051_golden_model_1.n2786 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2786 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2786 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2786 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2786 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2786 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2786 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2805 , \oc8051_golden_model_1.n2823 [7]);
  buf(\oc8051_golden_model_1.n2806 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2806 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2806 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2806 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2806 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2806 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2806 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2806 [7], \oc8051_golden_model_1.n2823 [7]);
  buf(\oc8051_golden_model_1.n2807 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2807 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2807 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2807 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2807 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2807 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2807 [6], \oc8051_golden_model_1.n2823 [7]);
  buf(\oc8051_golden_model_1.n2822 , \oc8051_golden_model_1.n2823 [0]);
  buf(\oc8051_golden_model_1.n2823 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2823 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2823 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2823 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2823 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2823 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2827 [0], \oc8051_golden_model_1.n2837 );
  buf(\oc8051_golden_model_1.n2827 [1], \oc8051_golden_model_1.n2836 );
  buf(\oc8051_golden_model_1.n2827 [2], \oc8051_golden_model_1.n2835 );
  buf(\oc8051_golden_model_1.n2827 [3], \oc8051_golden_model_1.n2834 );
  buf(\oc8051_golden_model_1.n2827 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2827 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2827 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2827 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2828 [0], \oc8051_golden_model_1.n2829 [4]);
  buf(\oc8051_golden_model_1.n2828 [1], \oc8051_golden_model_1.n2829 [5]);
  buf(\oc8051_golden_model_1.n2828 [2], \oc8051_golden_model_1.n2829 [6]);
  buf(\oc8051_golden_model_1.n2828 [3], \oc8051_golden_model_1.n2829 [7]);
  buf(\oc8051_golden_model_1.n2829 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2829 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2829 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2829 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2830 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2831 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2832 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2833 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2844 , \oc8051_golden_model_1.n2845 [0]);
  buf(\oc8051_golden_model_1.n2845 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2845 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2845 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2845 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2845 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2845 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2845 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2863 , \oc8051_golden_model_1.n2864 [0]);
  buf(\oc8051_golden_model_1.n2864 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2864 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2864 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2864 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2864 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2864 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2864 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2880 , \oc8051_golden_model_1.n2881 [0]);
  buf(\oc8051_golden_model_1.n2881 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2881 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2881 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2881 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2881 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2881 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2881 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(ie_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(ie_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(ie_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(ie_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(ie_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(ie_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(ie_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(ie_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
