
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_sp);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire _44029_;
  wire _44030_;
  wire _44031_;
  wire _44032_;
  wire _44033_;
  wire _44034_;
  wire _44035_;
  wire _44036_;
  wire _44037_;
  wire _44038_;
  wire _44039_;
  wire _44040_;
  wire _44041_;
  wire _44042_;
  wire _44043_;
  wire _44044_;
  wire _44045_;
  wire _44046_;
  wire _44047_;
  wire _44048_;
  wire _44049_;
  wire _44050_;
  wire _44051_;
  wire _44052_;
  wire _44053_;
  wire _44054_;
  wire _44055_;
  wire _44056_;
  wire _44057_;
  wire _44058_;
  wire _44059_;
  wire _44060_;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [6:0] \oc8051_golden_model_1.n0988 ;
  wire \oc8051_golden_model_1.n0989 ;
  wire \oc8051_golden_model_1.n0990 ;
  wire \oc8051_golden_model_1.n0991 ;
  wire \oc8051_golden_model_1.n0992 ;
  wire \oc8051_golden_model_1.n0993 ;
  wire \oc8051_golden_model_1.n0994 ;
  wire \oc8051_golden_model_1.n0995 ;
  wire \oc8051_golden_model_1.n0996 ;
  wire \oc8051_golden_model_1.n1003 ;
  wire [7:0] \oc8051_golden_model_1.n1004 ;
  wire [7:0] \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1017 ;
  wire \oc8051_golden_model_1.n1018 ;
  wire \oc8051_golden_model_1.n1019 ;
  wire \oc8051_golden_model_1.n1026 ;
  wire [7:0] \oc8051_golden_model_1.n1027 ;
  wire \oc8051_golden_model_1.n1043 ;
  wire [7:0] \oc8051_golden_model_1.n1044 ;
  wire [3:0] \oc8051_golden_model_1.n1137 ;
  wire [3:0] \oc8051_golden_model_1.n1139 ;
  wire [3:0] \oc8051_golden_model_1.n1141 ;
  wire [3:0] \oc8051_golden_model_1.n1142 ;
  wire [3:0] \oc8051_golden_model_1.n1143 ;
  wire [3:0] \oc8051_golden_model_1.n1144 ;
  wire [3:0] \oc8051_golden_model_1.n1145 ;
  wire [3:0] \oc8051_golden_model_1.n1146 ;
  wire [3:0] \oc8051_golden_model_1.n1147 ;
  wire \oc8051_golden_model_1.n1194 ;
  wire \oc8051_golden_model_1.n1239 ;
  wire [8:0] \oc8051_golden_model_1.n1240 ;
  wire [8:0] \oc8051_golden_model_1.n1241 ;
  wire [7:0] \oc8051_golden_model_1.n1242 ;
  wire \oc8051_golden_model_1.n1243 ;
  wire [2:0] \oc8051_golden_model_1.n1244 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [1:0] \oc8051_golden_model_1.n1246 ;
  wire [7:0] \oc8051_golden_model_1.n1247 ;
  wire [6:0] \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1251 ;
  wire \oc8051_golden_model_1.n1252 ;
  wire \oc8051_golden_model_1.n1253 ;
  wire \oc8051_golden_model_1.n1254 ;
  wire \oc8051_golden_model_1.n1255 ;
  wire \oc8051_golden_model_1.n1256 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [7:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1280 ;
  wire [7:0] \oc8051_golden_model_1.n1281 ;
  wire [15:0] \oc8051_golden_model_1.n1323 ;
  wire [7:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1327 ;
  wire \oc8051_golden_model_1.n1328 ;
  wire \oc8051_golden_model_1.n1329 ;
  wire \oc8051_golden_model_1.n1330 ;
  wire \oc8051_golden_model_1.n1331 ;
  wire \oc8051_golden_model_1.n1332 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire \oc8051_golden_model_1.n1340 ;
  wire [7:0] \oc8051_golden_model_1.n1341 ;
  wire [8:0] \oc8051_golden_model_1.n1343 ;
  wire [8:0] \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire [3:0] \oc8051_golden_model_1.n1349 ;
  wire [4:0] \oc8051_golden_model_1.n1350 ;
  wire [4:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [8:0] \oc8051_golden_model_1.n1356 ;
  wire \oc8051_golden_model_1.n1364 ;
  wire [7:0] \oc8051_golden_model_1.n1365 ;
  wire [6:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1381 ;
  wire [7:0] \oc8051_golden_model_1.n1382 ;
  wire [8:0] \oc8051_golden_model_1.n1404 ;
  wire \oc8051_golden_model_1.n1405 ;
  wire [4:0] \oc8051_golden_model_1.n1410 ;
  wire \oc8051_golden_model_1.n1411 ;
  wire \oc8051_golden_model_1.n1419 ;
  wire [7:0] \oc8051_golden_model_1.n1420 ;
  wire [6:0] \oc8051_golden_model_1.n1421 ;
  wire \oc8051_golden_model_1.n1436 ;
  wire [7:0] \oc8051_golden_model_1.n1437 ;
  wire [8:0] \oc8051_golden_model_1.n1439 ;
  wire [8:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1442 ;
  wire [3:0] \oc8051_golden_model_1.n1443 ;
  wire [4:0] \oc8051_golden_model_1.n1444 ;
  wire [4:0] \oc8051_golden_model_1.n1446 ;
  wire \oc8051_golden_model_1.n1447 ;
  wire [8:0] \oc8051_golden_model_1.n1448 ;
  wire \oc8051_golden_model_1.n1455 ;
  wire [7:0] \oc8051_golden_model_1.n1456 ;
  wire [6:0] \oc8051_golden_model_1.n1457 ;
  wire \oc8051_golden_model_1.n1472 ;
  wire [7:0] \oc8051_golden_model_1.n1473 ;
  wire [8:0] \oc8051_golden_model_1.n1476 ;
  wire \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1484 ;
  wire [7:0] \oc8051_golden_model_1.n1485 ;
  wire [6:0] \oc8051_golden_model_1.n1486 ;
  wire [7:0] \oc8051_golden_model_1.n1487 ;
  wire [8:0] \oc8051_golden_model_1.n1489 ;
  wire [8:0] \oc8051_golden_model_1.n1491 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [4:0] \oc8051_golden_model_1.n1493 ;
  wire [4:0] \oc8051_golden_model_1.n1495 ;
  wire \oc8051_golden_model_1.n1496 ;
  wire [8:0] \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1504 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire [4:0] \oc8051_golden_model_1.n1524 ;
  wire \oc8051_golden_model_1.n1525 ;
  wire [7:0] \oc8051_golden_model_1.n1526 ;
  wire [6:0] \oc8051_golden_model_1.n1527 ;
  wire [7:0] \oc8051_golden_model_1.n1528 ;
  wire [8:0] \oc8051_golden_model_1.n1530 ;
  wire \oc8051_golden_model_1.n1531 ;
  wire \oc8051_golden_model_1.n1538 ;
  wire [7:0] \oc8051_golden_model_1.n1539 ;
  wire [6:0] \oc8051_golden_model_1.n1540 ;
  wire [7:0] \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [6:0] \oc8051_golden_model_1.n1543 ;
  wire [7:0] \oc8051_golden_model_1.n1544 ;
  wire [8:0] \oc8051_golden_model_1.n1547 ;
  wire [8:0] \oc8051_golden_model_1.n1548 ;
  wire [7:0] \oc8051_golden_model_1.n1549 ;
  wire [7:0] \oc8051_golden_model_1.n1550 ;
  wire [6:0] \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1552 ;
  wire \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire \oc8051_golden_model_1.n1555 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire \oc8051_golden_model_1.n1557 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1559 ;
  wire \oc8051_golden_model_1.n1566 ;
  wire [7:0] \oc8051_golden_model_1.n1567 ;
  wire [7:0] \oc8051_golden_model_1.n1568 ;
  wire [8:0] \oc8051_golden_model_1.n1571 ;
  wire [8:0] \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire [4:0] \oc8051_golden_model_1.n1575 ;
  wire [4:0] \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1585 ;
  wire [7:0] \oc8051_golden_model_1.n1586 ;
  wire [6:0] \oc8051_golden_model_1.n1587 ;
  wire \oc8051_golden_model_1.n1602 ;
  wire [7:0] \oc8051_golden_model_1.n1603 ;
  wire [8:0] \oc8051_golden_model_1.n1607 ;
  wire \oc8051_golden_model_1.n1608 ;
  wire [4:0] \oc8051_golden_model_1.n1610 ;
  wire \oc8051_golden_model_1.n1611 ;
  wire \oc8051_golden_model_1.n1618 ;
  wire [7:0] \oc8051_golden_model_1.n1619 ;
  wire [6:0] \oc8051_golden_model_1.n1620 ;
  wire \oc8051_golden_model_1.n1635 ;
  wire [7:0] \oc8051_golden_model_1.n1636 ;
  wire [8:0] \oc8051_golden_model_1.n1640 ;
  wire \oc8051_golden_model_1.n1641 ;
  wire [4:0] \oc8051_golden_model_1.n1643 ;
  wire \oc8051_golden_model_1.n1644 ;
  wire \oc8051_golden_model_1.n1651 ;
  wire [7:0] \oc8051_golden_model_1.n1652 ;
  wire [6:0] \oc8051_golden_model_1.n1653 ;
  wire \oc8051_golden_model_1.n1668 ;
  wire [7:0] \oc8051_golden_model_1.n1669 ;
  wire [8:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1674 ;
  wire [4:0] \oc8051_golden_model_1.n1676 ;
  wire \oc8051_golden_model_1.n1677 ;
  wire \oc8051_golden_model_1.n1684 ;
  wire [7:0] \oc8051_golden_model_1.n1685 ;
  wire [6:0] \oc8051_golden_model_1.n1686 ;
  wire \oc8051_golden_model_1.n1701 ;
  wire [7:0] \oc8051_golden_model_1.n1702 ;
  wire [7:0] \oc8051_golden_model_1.n1727 ;
  wire [6:0] \oc8051_golden_model_1.n1728 ;
  wire [7:0] \oc8051_golden_model_1.n1729 ;
  wire \oc8051_golden_model_1.n1784 ;
  wire [7:0] \oc8051_golden_model_1.n1785 ;
  wire \oc8051_golden_model_1.n1801 ;
  wire [7:0] \oc8051_golden_model_1.n1802 ;
  wire \oc8051_golden_model_1.n1818 ;
  wire [7:0] \oc8051_golden_model_1.n1819 ;
  wire \oc8051_golden_model_1.n1835 ;
  wire [7:0] \oc8051_golden_model_1.n1836 ;
  wire [7:0] \oc8051_golden_model_1.n1859 ;
  wire [6:0] \oc8051_golden_model_1.n1860 ;
  wire [7:0] \oc8051_golden_model_1.n1861 ;
  wire \oc8051_golden_model_1.n1916 ;
  wire [7:0] \oc8051_golden_model_1.n1917 ;
  wire \oc8051_golden_model_1.n1933 ;
  wire [7:0] \oc8051_golden_model_1.n1934 ;
  wire \oc8051_golden_model_1.n1950 ;
  wire [7:0] \oc8051_golden_model_1.n1951 ;
  wire \oc8051_golden_model_1.n1967 ;
  wire [7:0] \oc8051_golden_model_1.n1968 ;
  wire \oc8051_golden_model_1.n2065 ;
  wire [7:0] \oc8051_golden_model_1.n2066 ;
  wire \oc8051_golden_model_1.n2082 ;
  wire [7:0] \oc8051_golden_model_1.n2083 ;
  wire \oc8051_golden_model_1.n2099 ;
  wire [7:0] \oc8051_golden_model_1.n2100 ;
  wire \oc8051_golden_model_1.n2116 ;
  wire [7:0] \oc8051_golden_model_1.n2117 ;
  wire \oc8051_golden_model_1.n2121 ;
  wire [6:0] \oc8051_golden_model_1.n2122 ;
  wire [7:0] \oc8051_golden_model_1.n2123 ;
  wire [6:0] \oc8051_golden_model_1.n2124 ;
  wire [7:0] \oc8051_golden_model_1.n2125 ;
  wire \oc8051_golden_model_1.n2140 ;
  wire [7:0] \oc8051_golden_model_1.n2141 ;
  wire \oc8051_golden_model_1.n2180 ;
  wire [7:0] \oc8051_golden_model_1.n2181 ;
  wire [6:0] \oc8051_golden_model_1.n2182 ;
  wire [7:0] \oc8051_golden_model_1.n2183 ;
  wire [3:0] \oc8051_golden_model_1.n2190 ;
  wire \oc8051_golden_model_1.n2191 ;
  wire [7:0] \oc8051_golden_model_1.n2192 ;
  wire [6:0] \oc8051_golden_model_1.n2193 ;
  wire \oc8051_golden_model_1.n2208 ;
  wire [7:0] \oc8051_golden_model_1.n2209 ;
  wire [7:0] \oc8051_golden_model_1.n2421 ;
  wire \oc8051_golden_model_1.n2424 ;
  wire \oc8051_golden_model_1.n2426 ;
  wire \oc8051_golden_model_1.n2432 ;
  wire [7:0] \oc8051_golden_model_1.n2433 ;
  wire [6:0] \oc8051_golden_model_1.n2434 ;
  wire \oc8051_golden_model_1.n2449 ;
  wire [7:0] \oc8051_golden_model_1.n2450 ;
  wire \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2456 ;
  wire \oc8051_golden_model_1.n2462 ;
  wire [7:0] \oc8051_golden_model_1.n2463 ;
  wire [6:0] \oc8051_golden_model_1.n2464 ;
  wire \oc8051_golden_model_1.n2479 ;
  wire [7:0] \oc8051_golden_model_1.n2480 ;
  wire \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2486 ;
  wire \oc8051_golden_model_1.n2492 ;
  wire [7:0] \oc8051_golden_model_1.n2493 ;
  wire [6:0] \oc8051_golden_model_1.n2494 ;
  wire \oc8051_golden_model_1.n2509 ;
  wire [7:0] \oc8051_golden_model_1.n2510 ;
  wire \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2516 ;
  wire \oc8051_golden_model_1.n2522 ;
  wire [7:0] \oc8051_golden_model_1.n2523 ;
  wire [6:0] \oc8051_golden_model_1.n2524 ;
  wire \oc8051_golden_model_1.n2539 ;
  wire [7:0] \oc8051_golden_model_1.n2540 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire [7:0] \oc8051_golden_model_1.n2545 ;
  wire [7:0] \oc8051_golden_model_1.n2546 ;
  wire [6:0] \oc8051_golden_model_1.n2547 ;
  wire [7:0] \oc8051_golden_model_1.n2548 ;
  wire [15:0] \oc8051_golden_model_1.n2552 ;
  wire \oc8051_golden_model_1.n2558 ;
  wire [7:0] \oc8051_golden_model_1.n2559 ;
  wire [6:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2575 ;
  wire [7:0] \oc8051_golden_model_1.n2576 ;
  wire \oc8051_golden_model_1.n2579 ;
  wire [7:0] \oc8051_golden_model_1.n2580 ;
  wire [6:0] \oc8051_golden_model_1.n2581 ;
  wire [7:0] \oc8051_golden_model_1.n2582 ;
  wire \oc8051_golden_model_1.n2614 ;
  wire [7:0] \oc8051_golden_model_1.n2615 ;
  wire [6:0] \oc8051_golden_model_1.n2616 ;
  wire [7:0] \oc8051_golden_model_1.n2617 ;
  wire \oc8051_golden_model_1.n2622 ;
  wire [7:0] \oc8051_golden_model_1.n2623 ;
  wire [6:0] \oc8051_golden_model_1.n2624 ;
  wire [7:0] \oc8051_golden_model_1.n2625 ;
  wire \oc8051_golden_model_1.n2630 ;
  wire [7:0] \oc8051_golden_model_1.n2631 ;
  wire [6:0] \oc8051_golden_model_1.n2632 ;
  wire [7:0] \oc8051_golden_model_1.n2633 ;
  wire \oc8051_golden_model_1.n2638 ;
  wire [7:0] \oc8051_golden_model_1.n2639 ;
  wire [6:0] \oc8051_golden_model_1.n2640 ;
  wire [7:0] \oc8051_golden_model_1.n2641 ;
  wire \oc8051_golden_model_1.n2646 ;
  wire [7:0] \oc8051_golden_model_1.n2647 ;
  wire [6:0] \oc8051_golden_model_1.n2648 ;
  wire [7:0] \oc8051_golden_model_1.n2649 ;
  wire [7:0] \oc8051_golden_model_1.n2674 ;
  wire [6:0] \oc8051_golden_model_1.n2675 ;
  wire [7:0] \oc8051_golden_model_1.n2676 ;
  wire [3:0] \oc8051_golden_model_1.n2677 ;
  wire [7:0] \oc8051_golden_model_1.n2678 ;
  wire \oc8051_golden_model_1.n2679 ;
  wire \oc8051_golden_model_1.n2680 ;
  wire \oc8051_golden_model_1.n2681 ;
  wire \oc8051_golden_model_1.n2682 ;
  wire \oc8051_golden_model_1.n2683 ;
  wire \oc8051_golden_model_1.n2684 ;
  wire \oc8051_golden_model_1.n2685 ;
  wire \oc8051_golden_model_1.n2686 ;
  wire \oc8051_golden_model_1.n2693 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire [6:0] \oc8051_golden_model_1.n2715 ;
  wire [7:0] \oc8051_golden_model_1.n2731 ;
  wire \oc8051_golden_model_1.n2732 ;
  wire \oc8051_golden_model_1.n2733 ;
  wire \oc8051_golden_model_1.n2734 ;
  wire \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2736 ;
  wire \oc8051_golden_model_1.n2737 ;
  wire \oc8051_golden_model_1.n2738 ;
  wire \oc8051_golden_model_1.n2739 ;
  wire \oc8051_golden_model_1.n2746 ;
  wire [7:0] \oc8051_golden_model_1.n2747 ;
  wire \oc8051_golden_model_1.n2748 ;
  wire \oc8051_golden_model_1.n2749 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2762 ;
  wire [7:0] \oc8051_golden_model_1.n2763 ;
  wire [7:0] \oc8051_golden_model_1.n2795 ;
  wire [6:0] \oc8051_golden_model_1.n2796 ;
  wire [7:0] \oc8051_golden_model_1.n2797 ;
  wire \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire [6:0] \oc8051_golden_model_1.n2818 ;
  wire \oc8051_golden_model_1.n2833 ;
  wire [7:0] \oc8051_golden_model_1.n2834 ;
  wire [7:0] \oc8051_golden_model_1.n2838 ;
  wire [3:0] \oc8051_golden_model_1.n2839 ;
  wire [7:0] \oc8051_golden_model_1.n2840 ;
  wire \oc8051_golden_model_1.n2841 ;
  wire \oc8051_golden_model_1.n2842 ;
  wire \oc8051_golden_model_1.n2843 ;
  wire \oc8051_golden_model_1.n2844 ;
  wire \oc8051_golden_model_1.n2845 ;
  wire \oc8051_golden_model_1.n2846 ;
  wire \oc8051_golden_model_1.n2847 ;
  wire \oc8051_golden_model_1.n2848 ;
  wire \oc8051_golden_model_1.n2855 ;
  wire [7:0] \oc8051_golden_model_1.n2856 ;
  wire \oc8051_golden_model_1.n2874 ;
  wire [7:0] \oc8051_golden_model_1.n2875 ;
  wire \oc8051_golden_model_1.n2891 ;
  wire [7:0] \oc8051_golden_model_1.n2892 ;
  wire [7:0] \oc8051_golden_model_1.n2893 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  wire property_invalid_psw_1_r;
  output property_invalid_sp;
  wire property_invalid_sp_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_41806_, rst);
  not (_15625_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_15636_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15647_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15636_);
  and (_15658_, _15647_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_15669_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15636_);
  and (_15680_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _15636_);
  nor (_15691_, _15680_, _15669_);
  and (_15702_, _15691_, _15658_);
  nor (_15713_, _15702_, _15625_);
  and (_15724_, _15625_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15735_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_15746_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _15735_);
  nor (_15757_, _15746_, _15724_);
  not (_15768_, _15757_);
  and (_15779_, _15768_, _15702_);
  or (_15790_, _15779_, _15713_);
  and (_22434_, _15790_, _41806_);
  nor (_15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15821_, _15810_);
  and (_15832_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_15843_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_15854_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_15865_, _15854_);
  not (_15876_, _15746_);
  nor (_15887_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_15898_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_15909_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _15898_);
  nor (_15920_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_15931_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_15942_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _15931_);
  nor (_15953_, _15942_, _15920_);
  nor (_15964_, _15953_, _15909_);
  not (_15975_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_15986_, _15909_, _15975_);
  nor (_15997_, _15986_, _15964_);
  and (_16008_, _15997_, _15887_);
  not (_16019_, _16008_);
  and (_16030_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16041_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_16052_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16063_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _16052_);
  and (_16074_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_16085_, _16074_, _16041_);
  and (_16096_, _16085_, _16019_);
  nor (_16107_, _16096_, _15876_);
  not (_16118_, _15724_);
  nor (_16128_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_16139_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _15931_);
  nor (_16150_, _16139_, _16128_);
  nor (_16161_, _16150_, _15909_);
  not (_16172_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_16183_, _15909_, _16172_);
  nor (_16194_, _16183_, _16161_);
  and (_16205_, _16194_, _15887_);
  not (_16216_, _16205_);
  and (_16227_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_16238_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_16249_, _16238_, _16227_);
  and (_16260_, _16249_, _16216_);
  nor (_16271_, _16260_, _16118_);
  nor (_16282_, _16271_, _16107_);
  nor (_16293_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_16304_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _15931_);
  nor (_16315_, _16304_, _16293_);
  nor (_16326_, _16315_, _15909_);
  not (_16337_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_16348_, _15909_, _16337_);
  nor (_16359_, _16348_, _16326_);
  and (_16370_, _16359_, _15887_);
  not (_16381_, _16370_);
  and (_16392_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_16403_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_16414_, _16403_, _16392_);
  and (_16425_, _16414_, _16381_);
  nor (_16436_, _16425_, _15768_);
  nor (_16446_, _16436_, _15810_);
  and (_16457_, _16446_, _16282_);
  nor (_16468_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_16479_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _15931_);
  nor (_16490_, _16479_, _16468_);
  nor (_16501_, _16490_, _15909_);
  not (_16512_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_16523_, _15909_, _16512_);
  nor (_16534_, _16523_, _16501_);
  and (_16556_, _16534_, _15887_);
  not (_16557_, _16556_);
  and (_16568_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_16579_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_16590_, _16579_, _16568_);
  and (_16601_, _16590_, _16557_);
  and (_16612_, _16601_, _15810_);
  nor (_16623_, _16612_, _16457_);
  not (_16634_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16645_, _16634_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16656_, _16645_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16667_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_16678_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16689_, _16678_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16700_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_16711_, _16700_, _16667_);
  nor (_16722_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16733_, _16722_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16744_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_16755_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16766_, _16645_, _16755_);
  and (_16776_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_16787_, _16776_, _16744_);
  and (_16798_, _16787_, _16711_);
  and (_16809_, _16722_, _16634_);
  and (_16820_, _16809_, _16534_);
  and (_16831_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16842_, _16831_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16853_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_16864_, _16831_, _16755_);
  and (_16875_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_16886_, _16875_, _16853_);
  not (_16897_, _16886_);
  nor (_16908_, _16897_, _16820_);
  and (_16919_, _16908_, _16798_);
  not (_16930_, _16919_);
  and (_16941_, _16930_, _16623_);
  not (_16952_, _16941_);
  nor (_16963_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_16974_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _15931_);
  nor (_16985_, _16974_, _16963_);
  nor (_16996_, _16985_, _15909_);
  not (_17007_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_17018_, _15909_, _17007_);
  nor (_17029_, _17018_, _16996_);
  and (_17040_, _17029_, _15887_);
  not (_17051_, _17040_);
  and (_17062_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_17073_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_17084_, _17073_, _17062_);
  and (_17094_, _17084_, _17051_);
  nor (_17105_, _17094_, _15876_);
  nor (_17116_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_17127_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _15931_);
  nor (_17138_, _17127_, _17116_);
  nor (_17149_, _17138_, _15909_);
  not (_17160_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_17171_, _15909_, _17160_);
  nor (_17181_, _17171_, _17149_);
  and (_17192_, _17181_, _15887_);
  not (_17203_, _17192_);
  and (_17214_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_17225_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17236_, _17225_, _17214_);
  and (_17247_, _17236_, _17203_);
  nor (_17258_, _17247_, _16118_);
  nor (_17278_, _17258_, _17105_);
  nor (_17279_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_17300_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _15931_);
  nor (_17301_, _17300_, _17279_);
  nor (_17312_, _17301_, _15909_);
  not (_17323_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_17334_, _15909_, _17323_);
  nor (_17345_, _17334_, _17312_);
  and (_17356_, _17345_, _15887_);
  not (_17366_, _17356_);
  and (_17377_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_17388_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_17399_, _17388_, _17377_);
  and (_17410_, _17399_, _17366_);
  nor (_17421_, _17410_, _15768_);
  nor (_17432_, _17421_, _15810_);
  and (_17443_, _17432_, _17278_);
  nor (_17454_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_17464_, _15931_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_17475_, _17464_, _17454_);
  nor (_17486_, _17475_, _15909_);
  not (_17497_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_17508_, _15909_, _17497_);
  nor (_17519_, _17508_, _17486_);
  and (_17530_, _17519_, _15887_);
  not (_17541_, _17530_);
  and (_17552_, _16030_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_17562_, _16063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_17573_, _17562_, _17552_);
  and (_17584_, _17573_, _17541_);
  and (_17595_, _17584_, _15810_);
  or (_17606_, _17595_, _17443_);
  and (_17617_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_17628_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_17639_, _17628_, _17617_);
  and (_17649_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_17660_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_17671_, _17660_, _17649_);
  and (_17682_, _17671_, _17639_);
  and (_17693_, _17519_, _16809_);
  and (_17704_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_17715_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_17726_, _17715_, _17704_);
  not (_17737_, _17726_);
  nor (_17747_, _17737_, _17693_);
  and (_17758_, _17747_, _17682_);
  nor (_17769_, _17758_, _17606_);
  and (_17780_, _17769_, _16952_);
  not (_17791_, _17780_);
  and (_17802_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_17813_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_17824_, _17813_, _17802_);
  and (_17834_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_17845_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_17856_, _17845_, _17834_);
  and (_17867_, _17856_, _17824_);
  and (_17878_, _17181_, _16809_);
  and (_17889_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_17900_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17911_, _17900_, _17889_);
  not (_17922_, _17911_);
  nor (_17932_, _17922_, _17878_);
  and (_17943_, _17932_, _17867_);
  nor (_17954_, _17943_, _17606_);
  and (_17965_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_17976_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_17987_, _17976_, _17965_);
  and (_17998_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_18009_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_18019_, _18009_, _17998_);
  and (_18030_, _18019_, _17987_);
  and (_18041_, _16809_, _16194_);
  and (_18052_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_18063_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_18074_, _18063_, _18052_);
  not (_18085_, _18074_);
  nor (_18096_, _18085_, _18041_);
  and (_18107_, _18096_, _18030_);
  not (_18117_, _18107_);
  and (_18128_, _18117_, _16623_);
  and (_18139_, _17954_, _18128_);
  and (_18150_, _16930_, _18139_);
  nor (_18161_, _16941_, _18139_);
  nor (_18172_, _18161_, _18150_);
  and (_18183_, _18172_, _17954_);
  and (_18194_, _17769_, _16941_);
  nor (_18204_, _16919_, _17606_);
  not (_18215_, _17758_);
  and (_18226_, _18215_, _16623_);
  nor (_18237_, _18226_, _18204_);
  nor (_18248_, _18237_, _18194_);
  and (_18259_, _18248_, _18183_);
  nor (_18270_, _18248_, _18183_);
  nor (_18281_, _18270_, _18259_);
  and (_18292_, _18281_, _18150_);
  nor (_18302_, _18292_, _18259_);
  nor (_18313_, _18302_, _17791_);
  nor (_18324_, _17606_, _18107_);
  and (_18335_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_18346_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_18357_, _18346_, _18335_);
  and (_18368_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_18379_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_18390_, _18379_, _18368_);
  and (_18400_, _18390_, _18357_);
  and (_18411_, _17029_, _16809_);
  and (_18422_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_18433_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_18444_, _18433_, _18422_);
  not (_18455_, _18444_);
  nor (_18466_, _18455_, _18411_);
  and (_18477_, _18466_, _18400_);
  not (_18488_, _18477_);
  and (_18498_, _18488_, _16623_);
  and (_18509_, _18498_, _18324_);
  not (_18520_, _17943_);
  and (_18531_, _18520_, _16623_);
  nor (_18542_, _18531_, _18324_);
  nor (_18553_, _18542_, _18139_);
  and (_18564_, _18553_, _18509_);
  nor (_18575_, _16941_, _17954_);
  nor (_18586_, _18575_, _18183_);
  and (_18597_, _18586_, _18564_);
  nor (_18608_, _18281_, _18150_);
  nor (_18618_, _18608_, _18292_);
  and (_18629_, _18618_, _18597_);
  nor (_18640_, _18618_, _18597_);
  nor (_18651_, _18640_, _18629_);
  not (_18662_, _18651_);
  and (_18673_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_18684_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_18695_, _18684_, _18673_);
  and (_18706_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_18717_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_18727_, _18717_, _18706_);
  and (_18738_, _18727_, _18695_);
  and (_18749_, _17345_, _16809_);
  and (_18760_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_18771_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_18782_, _18771_, _18760_);
  not (_18793_, _18782_);
  nor (_18804_, _18793_, _18749_);
  and (_18815_, _18804_, _18738_);
  nor (_18826_, _18815_, _17606_);
  and (_18837_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_18847_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_18858_, _18847_, _18837_);
  and (_18869_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_18880_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_18891_, _18880_, _18869_);
  and (_18902_, _18891_, _18858_);
  and (_18913_, _16809_, _15997_);
  and (_18924_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_18935_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_18946_, _18935_, _18924_);
  not (_18957_, _18946_);
  nor (_18967_, _18957_, _18913_);
  and (_18978_, _18967_, _18902_);
  not (_18989_, _18978_);
  and (_19000_, _18989_, _16623_);
  and (_19011_, _19000_, _18826_);
  not (_19022_, _18815_);
  and (_19033_, _19022_, _16623_);
  not (_19044_, _19033_);
  nor (_19055_, _18978_, _17606_);
  and (_19066_, _19055_, _19044_);
  and (_19076_, _19066_, _18498_);
  nor (_19087_, _19076_, _19011_);
  nor (_19098_, _18477_, _17606_);
  nor (_19109_, _19098_, _18128_);
  nor (_19120_, _19109_, _18509_);
  not (_19131_, _19120_);
  nor (_19142_, _19131_, _19087_);
  nor (_19153_, _18553_, _18509_);
  nor (_19164_, _19153_, _18564_);
  and (_19175_, _19164_, _19142_);
  nor (_19186_, _18586_, _18564_);
  nor (_19196_, _19186_, _18597_);
  and (_19207_, _19196_, _19175_);
  and (_19218_, _16656_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_19229_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_19240_, _19229_, _19218_);
  and (_19251_, _16733_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_19262_, _16766_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_19273_, _19262_, _19251_);
  and (_19284_, _19273_, _19240_);
  and (_19294_, _16809_, _16359_);
  and (_19305_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_19316_, _16842_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_19327_, _19316_, _19305_);
  not (_19338_, _19327_);
  nor (_19349_, _19338_, _19294_);
  and (_19360_, _19349_, _19284_);
  nor (_19371_, _19360_, _17606_);
  and (_19382_, _19371_, _19033_);
  nor (_19393_, _19000_, _18826_);
  nor (_19404_, _19393_, _19011_);
  and (_19414_, _19404_, _19382_);
  nor (_19425_, _19066_, _18498_);
  nor (_19436_, _19425_, _19076_);
  and (_19447_, _19436_, _19414_);
  and (_19458_, _19131_, _19087_);
  nor (_19469_, _19458_, _19142_);
  and (_19480_, _19469_, _19447_);
  nor (_19491_, _19164_, _19142_);
  nor (_19502_, _19491_, _19175_);
  and (_19513_, _19502_, _19480_);
  nor (_19523_, _19196_, _19175_);
  nor (_19534_, _19523_, _19207_);
  and (_19545_, _19534_, _19513_);
  nor (_19556_, _19545_, _19207_);
  nor (_19567_, _19556_, _18662_);
  nor (_19578_, _19567_, _18629_);
  and (_19589_, _18302_, _17791_);
  nor (_19600_, _19589_, _18313_);
  not (_19611_, _19600_);
  nor (_19622_, _19611_, _19578_);
  or (_19633_, _19622_, _18194_);
  nor (_19643_, _19633_, _18313_);
  nor (_19654_, _19643_, _15865_);
  and (_19665_, _19643_, _15865_);
  nor (_19676_, _19665_, _19654_);
  not (_19687_, _19676_);
  and (_19698_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_19709_, _19611_, _19578_);
  nor (_19720_, _19709_, _19622_);
  and (_19731_, _19720_, _19698_);
  and (_19742_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_19753_, _19556_, _18662_);
  nor (_19763_, _19753_, _19567_);
  and (_19774_, _19763_, _19742_);
  nor (_19785_, _19763_, _19742_);
  nor (_19796_, _19785_, _19774_);
  not (_19807_, _19796_);
  and (_19818_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_19829_, _19534_, _19513_);
  nor (_19840_, _19829_, _19545_);
  and (_19851_, _19840_, _19818_);
  nor (_19862_, _19840_, _19818_);
  nor (_19872_, _19862_, _19851_);
  not (_19883_, _19872_);
  and (_19894_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_19905_, _19502_, _19480_);
  nor (_19916_, _19905_, _19513_);
  and (_19927_, _19916_, _19894_);
  nor (_19938_, _19916_, _19894_);
  nor (_19949_, _19938_, _19927_);
  not (_19960_, _19949_);
  and (_19971_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_19981_, _19469_, _19447_);
  nor (_19992_, _19981_, _19480_);
  and (_20003_, _19992_, _19971_);
  and (_20014_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_20025_, _19436_, _19414_);
  nor (_20036_, _20025_, _19447_);
  and (_20047_, _20036_, _20014_);
  and (_20058_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_20069_, _19404_, _19382_);
  nor (_20080_, _20069_, _19414_);
  and (_20091_, _20080_, _20058_);
  nor (_20101_, _20036_, _20014_);
  nor (_20112_, _20101_, _20047_);
  and (_20123_, _20112_, _20091_);
  nor (_20134_, _20123_, _20047_);
  not (_20145_, _20134_);
  nor (_20156_, _19992_, _19971_);
  nor (_20167_, _20156_, _20003_);
  and (_20178_, _20167_, _20145_);
  nor (_20189_, _20178_, _20003_);
  nor (_20200_, _20189_, _19960_);
  nor (_20211_, _20200_, _19927_);
  nor (_20222_, _20211_, _19883_);
  nor (_20232_, _20222_, _19851_);
  nor (_20243_, _20232_, _19807_);
  nor (_20254_, _20243_, _19774_);
  nor (_20265_, _19720_, _19698_);
  nor (_20276_, _20265_, _19731_);
  not (_20287_, _20276_);
  nor (_20298_, _20287_, _20254_);
  nor (_20309_, _20298_, _19731_);
  nor (_20320_, _20309_, _19687_);
  nor (_20331_, _20320_, _19654_);
  not (_20342_, _20331_);
  and (_20352_, _20342_, _15843_);
  and (_20363_, _20352_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_20374_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_20385_, _20374_, _20363_);
  and (_20396_, _20385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_20407_, _20396_, _15832_);
  and (_20418_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20429_, _20418_, _20407_);
  and (_20440_, _20407_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20451_, _20440_, _20429_);
  and (_24620_, _20451_, _41806_);
  nor (_20471_, _15702_, _15735_);
  and (_20482_, _15702_, _15735_);
  or (_20493_, _20482_, _20471_);
  and (_02465_, _20493_, _41806_);
  not (_20514_, _19360_);
  and (_20525_, _20514_, _16623_);
  and (_02660_, _20525_, _41806_);
  nor (_20546_, _19371_, _19033_);
  nor (_20557_, _20546_, _19382_);
  and (_02854_, _20557_, _41806_);
  nor (_20578_, _20080_, _20058_);
  nor (_20589_, _20578_, _20091_);
  and (_03057_, _20589_, _41806_);
  nor (_20609_, _20112_, _20091_);
  nor (_20620_, _20609_, _20123_);
  and (_03268_, _20620_, _41806_);
  nor (_20641_, _20167_, _20145_);
  nor (_20652_, _20641_, _20178_);
  and (_03469_, _20652_, _41806_);
  and (_20673_, _20189_, _19960_);
  nor (_20684_, _20673_, _20200_);
  and (_03670_, _20684_, _41806_);
  and (_20705_, _20211_, _19883_);
  nor (_20715_, _20705_, _20222_);
  and (_03871_, _20715_, _41806_);
  and (_20736_, _20232_, _19807_);
  nor (_20747_, _20736_, _20243_);
  and (_04072_, _20747_, _41806_);
  and (_20768_, _20287_, _20254_);
  nor (_20779_, _20768_, _20298_);
  and (_04173_, _20779_, _41806_);
  and (_20800_, _20309_, _19687_);
  nor (_20811_, _20800_, _20320_);
  and (_04274_, _20811_, _41806_);
  nor (_20832_, _20342_, _15843_);
  nor (_20842_, _20832_, _20352_);
  and (_04375_, _20842_, _41806_);
  and (_20863_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_20874_, _20863_, _20352_);
  nor (_20885_, _20874_, _20363_);
  and (_04476_, _20885_, _41806_);
  nor (_20906_, _20374_, _20363_);
  nor (_20917_, _20906_, _20385_);
  and (_04577_, _20917_, _41806_);
  and (_20937_, _15821_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_20948_, _20937_, _20385_);
  nor (_20959_, _20948_, _20396_);
  and (_04678_, _20959_, _41806_);
  nor (_20980_, _20396_, _15832_);
  nor (_20991_, _20980_, _20407_);
  and (_04779_, _20991_, _41806_);
  and (_21012_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15636_);
  nor (_21023_, _21012_, _15647_);
  not (_21034_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_21044_, _15669_, _21034_);
  and (_21055_, _21044_, _21023_);
  and (_21066_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_21077_, _21066_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21088_, _21066_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21099_, _21088_, _21077_);
  and (_00862_, _21099_, _41806_);
  and (_00893_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _41806_);
  not (_21130_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_21141_, _17410_, _21130_);
  and (_21152_, _17094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21162_, _21152_, _21141_);
  nor (_21173_, _21162_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21184_, _17247_, _21130_);
  and (_21195_, _17584_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_21206_, _21195_, _21184_);
  and (_21217_, _21206_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21228_, _21217_, _21173_);
  nor (_21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_21250_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and (_21261_, _21239_, _17758_);
  nor (_21271_, _21261_, _21250_);
  not (_21282_, _21271_);
  and (_21293_, _16425_, _21130_);
  and (_21304_, _16096_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21315_, _21304_, _21293_);
  nor (_21326_, _21315_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21337_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21348_, _16260_, _21130_);
  and (_21359_, _16601_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21370_, _21359_, _21348_);
  nor (_21380_, _21370_, _21337_);
  nor (_21391_, _21380_, _21326_);
  nor (_21402_, _21391_, _21282_);
  and (_21413_, _21391_, _21282_);
  nor (_21424_, _21413_, _21402_);
  nor (_21435_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and (_21446_, _21239_, _16919_);
  nor (_21457_, _21446_, _21435_);
  not (_21468_, _21457_);
  nor (_21489_, _17410_, _21130_);
  nor (_21501_, _21489_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21513_, _17094_, _21130_);
  and (_21525_, _17247_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21537_, _21525_, _21513_);
  nor (_21549_, _21537_, _21337_);
  nor (_21550_, _21549_, _21501_);
  nor (_21561_, _21550_, _21468_);
  and (_21572_, _21550_, _21468_);
  nor (_21583_, _21572_, _21561_);
  not (_21594_, _21583_);
  nor (_21604_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_21615_, _21239_, _17943_);
  nor (_21626_, _21615_, _21604_);
  not (_21637_, _21626_);
  nor (_21648_, _16425_, _21130_);
  nor (_21659_, _21648_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21670_, _16096_, _21130_);
  and (_21681_, _16260_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21692_, _21681_, _21670_);
  nor (_21703_, _21692_, _21337_);
  nor (_21713_, _21703_, _21659_);
  nor (_21724_, _21713_, _21637_);
  and (_21735_, _21713_, _21637_);
  nor (_21746_, _21735_, _21724_);
  not (_21757_, _21746_);
  and (_21768_, _21162_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21779_, _21768_);
  nor (_21790_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_21801_, _21239_, _18107_);
  nor (_21812_, _21801_, _21790_);
  and (_21822_, _21812_, _21779_);
  and (_21833_, _21315_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21844_, _21833_);
  and (_21855_, _21239_, _18477_);
  nor (_21866_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_21877_, _21866_, _21855_);
  and (_21888_, _21877_, _21844_);
  nor (_21899_, _21877_, _21844_);
  nor (_21910_, _21899_, _21888_);
  not (_21921_, _21910_);
  and (_21931_, _21489_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21942_, _21931_);
  and (_21953_, _21239_, _18978_);
  nor (_21964_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_21975_, _21964_, _21953_);
  and (_21986_, _21975_, _21942_);
  and (_21997_, _21648_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_22008_, _21997_);
  nor (_22019_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_22030_, _21239_, _18815_);
  nor (_22040_, _22030_, _22019_);
  nor (_22061_, _22040_, _22008_);
  not (_22062_, _22061_);
  nor (_22073_, _21975_, _21942_);
  nor (_22084_, _22073_, _21986_);
  and (_22095_, _22084_, _22062_);
  nor (_22106_, _22095_, _21986_);
  nor (_22117_, _22106_, _21921_);
  nor (_22128_, _22117_, _21888_);
  nor (_22139_, _21812_, _21779_);
  nor (_22150_, _22139_, _21822_);
  not (_22160_, _22150_);
  nor (_22171_, _22160_, _22128_);
  nor (_22182_, _22171_, _21822_);
  nor (_22193_, _22182_, _21757_);
  nor (_22204_, _22193_, _21724_);
  nor (_22215_, _22204_, _21594_);
  nor (_22226_, _22215_, _21561_);
  not (_22237_, _22226_);
  and (_22248_, _22237_, _21424_);
  or (_22259_, _22248_, _21402_);
  and (_22269_, _17584_, _16601_);
  or (_22280_, _22269_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_22291_, _21370_);
  and (_22302_, _21206_, _22291_);
  nor (_22324_, _21692_, _21537_);
  and (_22325_, _22324_, _22302_);
  or (_22336_, _22325_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_22347_, _22336_, _22280_);
  and (_22358_, _22347_, _22259_);
  and (_22369_, _22358_, _21228_);
  nor (_22379_, _22237_, _21424_);
  or (_22390_, _22379_, _22248_);
  and (_22401_, _22390_, _22369_);
  nor (_22412_, _22369_, _21271_);
  nor (_22423_, _22412_, _22401_);
  not (_22435_, _22423_);
  and (_22446_, _22423_, _21228_);
  not (_22457_, _21391_);
  and (_22468_, _22204_, _21594_);
  or (_22478_, _22468_, _22215_);
  and (_22489_, _22478_, _22369_);
  nor (_22500_, _22369_, _21457_);
  nor (_22511_, _22500_, _22489_);
  and (_22522_, _22511_, _22457_);
  nor (_22533_, _22511_, _22457_);
  nor (_22544_, _22533_, _22522_);
  not (_22555_, _22544_);
  not (_22566_, _21550_);
  nor (_22577_, _22369_, _21637_);
  and (_22588_, _22182_, _21757_);
  nor (_22598_, _22588_, _22193_);
  and (_22609_, _22598_, _22369_);
  or (_22620_, _22609_, _22577_);
  and (_22631_, _22620_, _22566_);
  nor (_22642_, _22620_, _22566_);
  nor (_22653_, _22642_, _22631_);
  not (_22664_, _22653_);
  not (_22675_, _21713_);
  and (_22686_, _22160_, _22128_);
  or (_22697_, _22686_, _22171_);
  and (_22707_, _22697_, _22369_);
  nor (_22718_, _22369_, _21812_);
  nor (_22729_, _22718_, _22707_);
  and (_22740_, _22729_, _22675_);
  and (_22751_, _22106_, _21921_);
  nor (_22762_, _22751_, _22117_);
  not (_22773_, _22762_);
  and (_22784_, _22773_, _22369_);
  nor (_22795_, _22369_, _21877_);
  nor (_22806_, _22795_, _22784_);
  and (_22816_, _22806_, _21779_);
  nor (_22827_, _22806_, _21779_);
  nor (_22838_, _22827_, _22816_);
  not (_22849_, _22838_);
  nor (_22860_, _22084_, _22062_);
  nor (_22871_, _22860_, _22095_);
  not (_22882_, _22871_);
  and (_22893_, _22882_, _22369_);
  nor (_22904_, _22369_, _21975_);
  nor (_22915_, _22904_, _22893_);
  and (_22925_, _22915_, _21844_);
  not (_22936_, _22040_);
  and (_22947_, _22369_, _21997_);
  or (_22958_, _22947_, _22936_);
  nand (_22969_, _22369_, _21997_);
  or (_22980_, _22969_, _22040_);
  and (_23001_, _22980_, _22958_);
  nor (_23002_, _23001_, _21931_);
  and (_23013_, _23001_, _21931_);
  nor (_23033_, _23013_, _23002_);
  and (_23034_, _21239_, _19360_);
  nor (_23045_, _21239_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_23066_, _23045_, _23034_);
  nor (_23067_, _23066_, _22008_);
  not (_23078_, _23067_);
  and (_23099_, _23078_, _23033_);
  nor (_23100_, _23099_, _23002_);
  nor (_23111_, _22915_, _21844_);
  nor (_23132_, _23111_, _22925_);
  not (_23133_, _23132_);
  nor (_23143_, _23133_, _23100_);
  nor (_23164_, _23143_, _22925_);
  nor (_23165_, _23164_, _22849_);
  nor (_23176_, _23165_, _22816_);
  nor (_23197_, _22729_, _22675_);
  nor (_23198_, _23197_, _22740_);
  not (_23209_, _23198_);
  nor (_23220_, _23209_, _23176_);
  nor (_23231_, _23220_, _22740_);
  nor (_23242_, _23231_, _22664_);
  nor (_23253_, _23242_, _22631_);
  nor (_23264_, _23253_, _22555_);
  or (_23275_, _23264_, _22522_);
  or (_23286_, _23275_, _22446_);
  and (_23297_, _23286_, _22347_);
  nor (_23308_, _23297_, _22435_);
  and (_23319_, _22446_, _22347_);
  and (_23330_, _23319_, _23275_);
  or (_23341_, _23330_, _23308_);
  and (_00914_, _23341_, _41806_);
  or (_23362_, _22423_, _21228_);
  and (_23373_, _23362_, _23297_);
  and (_03014_, _23373_, _41806_);
  and (_03025_, _22369_, _41806_);
  and (_03046_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _41806_);
  and (_03068_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _41806_);
  and (_03089_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _41806_);
  or (_23434_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23445_, _21066_, rst);
  and (_03100_, _23445_, _23434_);
  and (_23466_, _23373_, _21997_);
  or (_23477_, _23466_, _23066_);
  nand (_23488_, _23466_, _23066_);
  and (_23499_, _23488_, _23477_);
  and (_03111_, _23499_, _41806_);
  nor (_23520_, _23373_, _23001_);
  nor (_23531_, _23078_, _23033_);
  nor (_23542_, _23531_, _23099_);
  and (_23553_, _23542_, _23373_);
  or (_23564_, _23553_, _23520_);
  and (_03122_, _23564_, _41806_);
  and (_23585_, _23133_, _23100_);
  or (_23596_, _23585_, _23143_);
  nand (_23607_, _23596_, _23373_);
  or (_23618_, _23373_, _22915_);
  and (_23629_, _23618_, _23607_);
  and (_03133_, _23629_, _41806_);
  and (_23650_, _23164_, _22849_);
  or (_23661_, _23650_, _23165_);
  nand (_23672_, _23661_, _23373_);
  or (_23683_, _23373_, _22806_);
  and (_23694_, _23683_, _23672_);
  and (_03144_, _23694_, _41806_);
  and (_23715_, _23209_, _23176_);
  or (_23726_, _23715_, _23220_);
  nand (_23737_, _23726_, _23373_);
  or (_23748_, _23373_, _22729_);
  and (_23759_, _23748_, _23737_);
  and (_03155_, _23759_, _41806_);
  and (_23780_, _23231_, _22664_);
  or (_23791_, _23780_, _23242_);
  nand (_23802_, _23791_, _23373_);
  or (_23813_, _23373_, _22620_);
  and (_23824_, _23813_, _23802_);
  and (_03166_, _23824_, _41806_);
  and (_23845_, _23253_, _22555_);
  or (_23856_, _23845_, _23264_);
  nand (_23867_, _23856_, _23373_);
  or (_23878_, _23373_, _22511_);
  and (_23889_, _23878_, _23867_);
  and (_03177_, _23889_, _41806_);
  not (_23910_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23921_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15636_);
  and (_23932_, _23921_, _23910_);
  and (_23943_, _23932_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_23954_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23965_, _23954_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_23976_, _23954_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_23987_, _23976_, _23965_);
  and (_23998_, _23987_, _23943_);
  nor (_24009_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24020_, _24009_, _23921_);
  and (_24031_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24042_, _24031_, _23998_);
  not (_24053_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_24064_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15636_);
  and (_24075_, _24064_, _24053_);
  and (_24086_, _24075_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24097_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_24108_, _24075_, _23910_);
  and (_24119_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  nor (_24130_, _24009_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_24141_, _24130_, _23921_);
  and (_24152_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_24163_, _24152_, _24119_);
  nor (_24185_, _24163_, _24097_);
  and (_24197_, _24185_, _24042_);
  and (_24209_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_24221_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24233_, _24221_, _23954_);
  and (_24245_, _24233_, _23943_);
  nor (_24257_, _24245_, _24209_);
  and (_24258_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_24269_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_24280_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_24291_, _24280_, _24269_);
  nor (_24302_, _24291_, _24258_);
  and (_24313_, _24302_, _24257_);
  and (_24324_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_24335_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_24346_, _24335_, _24324_);
  and (_24357_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_24368_, _24357_);
  not (_24379_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24390_, _23943_, _24379_);
  and (_24401_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_24412_, _24401_, _24390_);
  and (_24423_, _24412_, _24368_);
  and (_24434_, _24423_, _24346_);
  and (_24445_, _24434_, _24313_);
  and (_24456_, _24445_, _24197_);
  and (_24467_, _23965_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_24478_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_24489_, _24478_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_24500_, _24489_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_24511_, _24500_);
  not (_24522_, _23943_);
  nor (_24533_, _24489_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_24544_, _24533_, _24522_);
  and (_24555_, _24544_, _24511_);
  not (_24566_, _24555_);
  and (_24577_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24587_, _24577_, _23921_);
  and (_24598_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_24609_, _24598_, _24587_);
  and (_24621_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_24632_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_24643_, _24632_, _24621_);
  and (_24654_, _24643_, _24609_);
  and (_24665_, _24654_, _24566_);
  nor (_24676_, _24478_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_24687_, _24676_);
  nor (_24697_, _24489_, _24522_);
  and (_24708_, _24697_, _24687_);
  not (_24719_, _24708_);
  and (_24730_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_24741_, _24730_, _24587_);
  and (_24752_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_24763_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_24774_, _24763_, _24752_);
  and (_24785_, _24774_, _24741_);
  and (_24796_, _24785_, _24719_);
  nor (_24807_, _24796_, _24665_);
  not (_24818_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_24829_, _24500_, _24818_);
  and (_24840_, _24500_, _24818_);
  nor (_24851_, _24840_, _24829_);
  nor (_24862_, _24851_, _24522_);
  not (_24873_, _24862_);
  and (_24884_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_24895_, _24884_, _24587_);
  and (_24906_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_24917_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_24928_, _24917_, _24906_);
  and (_24938_, _24928_, _24895_);
  and (_24949_, _24938_, _24873_);
  not (_24960_, _24949_);
  not (_24971_, _24467_);
  nor (_24982_, _23965_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_24993_, _24982_, _24522_);
  and (_25004_, _24993_, _24971_);
  not (_25015_, _25004_);
  and (_25026_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and (_25037_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_25048_, _25037_, _25026_);
  and (_25058_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_25069_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_25080_, _25069_, _25058_);
  and (_25091_, _25080_, _25048_);
  and (_25112_, _25091_, _25015_);
  not (_25113_, _25112_);
  nor (_25124_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_25135_, _25124_, _24522_);
  nor (_25156_, _25135_, _24478_);
  and (_25157_, _24086_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_25168_, _25157_, _25156_);
  and (_25188_, _24108_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and (_25189_, _24141_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_25200_, _25189_, _25188_);
  and (_25211_, _24020_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_25222_, _25211_, _24587_);
  and (_25243_, _25222_, _25200_);
  and (_25244_, _25243_, _25168_);
  nor (_25255_, _25244_, _25113_);
  and (_25266_, _25255_, _24960_);
  and (_25277_, _25266_, _24807_);
  nand (_25287_, _25277_, _24456_);
  and (_25298_, _23341_, _21055_);
  not (_25309_, _25298_);
  and (_25320_, _20451_, _15702_);
  not (_25331_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_25342_, _15647_, _25331_);
  and (_25353_, _25342_, _15691_);
  not (_25374_, _25353_);
  nor (_25375_, _17758_, _17584_);
  and (_25386_, _17758_, _17584_);
  nor (_25397_, _25386_, _25375_);
  not (_25408_, _16601_);
  nor (_25419_, _16919_, _25408_);
  nor (_25430_, _16919_, _16601_);
  and (_25441_, _16919_, _16601_);
  nor (_25452_, _25441_, _25430_);
  not (_25462_, _17247_);
  nor (_25473_, _17943_, _25462_);
  nor (_25484_, _17943_, _17247_);
  and (_25495_, _17943_, _17247_);
  nor (_25506_, _25495_, _25484_);
  not (_25517_, _16260_);
  and (_25528_, _18107_, _25517_);
  nor (_25548_, _25528_, _25506_);
  nor (_25549_, _25548_, _25473_);
  nor (_25560_, _25549_, _25452_);
  nor (_25571_, _25560_, _25419_);
  and (_25582_, _25549_, _25452_);
  nor (_25593_, _25582_, _25560_);
  not (_25604_, _25593_);
  and (_25615_, _25528_, _25506_);
  nor (_25626_, _25615_, _25548_);
  not (_25636_, _25626_);
  nor (_25647_, _18107_, _16260_);
  and (_25658_, _18107_, _16260_);
  nor (_25669_, _25658_, _25647_);
  not (_25680_, _25669_);
  and (_25691_, _18477_, _17094_);
  nor (_25702_, _18477_, _17094_);
  nor (_25713_, _25702_, _25691_);
  nor (_25723_, _18978_, _16096_);
  and (_25744_, _18978_, _16096_);
  nor (_25745_, _25744_, _25723_);
  nor (_25756_, _18815_, _17410_);
  and (_25767_, _18815_, _17410_);
  nor (_25778_, _25767_, _25756_);
  not (_25789_, _16425_);
  and (_25800_, _19360_, _25789_);
  nor (_25810_, _25800_, _25778_);
  not (_25821_, _17410_);
  nor (_25832_, _18815_, _25821_);
  nor (_25843_, _25832_, _25810_);
  nor (_25854_, _25843_, _25745_);
  not (_25865_, _16096_);
  nor (_25876_, _18978_, _25865_);
  nor (_25887_, _25876_, _25854_);
  nor (_25897_, _25887_, _25713_);
  and (_25908_, _25887_, _25713_);
  nor (_25919_, _25908_, _25897_);
  not (_25930_, _25919_);
  and (_25941_, _25843_, _25745_);
  nor (_25952_, _25941_, _25854_);
  not (_25963_, _25952_);
  and (_25974_, _25800_, _25778_);
  nor (_25984_, _25974_, _25810_);
  not (_25995_, _25984_);
  nor (_26006_, _19360_, _16425_);
  and (_26017_, _19360_, _16425_);
  nor (_26028_, _26017_, _26006_);
  not (_26039_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_26050_, _15909_, _26039_);
  not (_26061_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26071_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26092_, _26071_, _17475_);
  nor (_26093_, _26092_, _26061_);
  nor (_26104_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26115_, _26104_, _16150_);
  not (_26126_, _26115_);
  not (_26137_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_26147_, _26137_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26158_, _26147_, _16490_);
  not (_26169_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26180_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _26169_);
  and (_26201_, _26180_, _17138_);
  nor (_26202_, _26201_, _26158_);
  and (_26213_, _26202_, _26126_);
  and (_26224_, _26213_, _26093_);
  and (_26234_, _26071_, _16985_);
  nor (_26245_, _26234_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26256_, _26180_, _17301_);
  not (_26267_, _26256_);
  and (_26278_, _26147_, _15953_);
  and (_26289_, _26104_, _16315_);
  nor (_26300_, _26289_, _26278_);
  and (_26311_, _26300_, _26267_);
  and (_26321_, _26311_, _26245_);
  nor (_26332_, _26321_, _26224_);
  nor (_26343_, _26332_, _15909_);
  nor (_26354_, _26343_, _26050_);
  and (_26365_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_26376_, _26365_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_26387_, _26376_);
  and (_26398_, _26387_, _26354_);
  and (_26408_, _26387_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_26419_, _26408_, _26398_);
  nor (_26430_, _26419_, _26028_);
  and (_26441_, _26430_, _25995_);
  and (_26452_, _26441_, _25963_);
  and (_26463_, _26452_, _25930_);
  not (_26474_, _17094_);
  or (_26485_, _18477_, _26474_);
  and (_26496_, _18477_, _26474_);
  or (_26506_, _25887_, _26496_);
  and (_26517_, _26506_, _26485_);
  or (_26528_, _26517_, _26463_);
  and (_26539_, _26528_, _25680_);
  and (_26550_, _26539_, _25636_);
  and (_26561_, _26550_, _25604_);
  nor (_26572_, _26561_, _25571_);
  nor (_26583_, _26572_, _25397_);
  and (_26593_, _26572_, _25397_);
  nor (_26604_, _26593_, _26583_);
  nor (_26615_, _26604_, _25374_);
  not (_26626_, _26615_);
  not (_26647_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_26648_, _21012_, _26647_);
  and (_26659_, _26648_, _15691_);
  not (_26670_, _25452_);
  and (_26680_, _25647_, _25506_);
  nor (_26691_, _26680_, _25484_);
  nor (_26702_, _26691_, _26670_);
  not (_26713_, _25745_);
  and (_26724_, _26006_, _25778_);
  nor (_26735_, _26724_, _25756_);
  nor (_26746_, _26735_, _26713_);
  nor (_26757_, _26746_, _25723_);
  nor (_26768_, _26757_, _25713_);
  and (_26778_, _26757_, _25713_);
  nor (_26789_, _26778_, _26768_);
  not (_26800_, _26028_);
  nor (_26811_, _26419_, _26800_);
  and (_26822_, _26811_, _25778_);
  and (_26833_, _26735_, _26713_);
  nor (_26844_, _26833_, _26746_);
  and (_26855_, _26844_, _26822_);
  not (_26866_, _26855_);
  nor (_26877_, _26866_, _26789_);
  nor (_26888_, _26757_, _25691_);
  or (_26898_, _26888_, _25702_);
  or (_26909_, _26898_, _26877_);
  and (_26920_, _26909_, _25669_);
  nor (_26941_, _25647_, _25506_);
  nor (_26942_, _26941_, _26680_);
  and (_26953_, _26942_, _26920_);
  and (_26964_, _26691_, _26670_);
  nor (_26975_, _26964_, _26702_);
  and (_26986_, _26975_, _26953_);
  or (_26997_, _26986_, _26702_);
  nor (_27007_, _26997_, _25430_);
  and (_27018_, _27007_, _25397_);
  nor (_27029_, _27007_, _25397_);
  or (_27050_, _27029_, _27018_);
  and (_27051_, _27050_, _26659_);
  and (_27062_, _15680_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27073_, _27062_, _25342_);
  nor (_27084_, _19360_, _18815_);
  and (_27095_, _27084_, _18989_);
  and (_27106_, _27095_, _18488_);
  and (_27117_, _27106_, _18117_);
  and (_27127_, _27117_, _18520_);
  and (_27138_, _27127_, _16930_);
  and (_27149_, _27138_, _26419_);
  not (_27160_, _26419_);
  and (_27171_, _16919_, _17943_);
  and (_27182_, _19360_, _18815_);
  and (_27193_, _27182_, _18978_);
  and (_27204_, _27193_, _18477_);
  and (_27215_, _27204_, _18107_);
  and (_27226_, _27215_, _27171_);
  and (_27237_, _27226_, _27160_);
  nor (_27247_, _27237_, _27149_);
  and (_27268_, _27247_, _17758_);
  nor (_27269_, _27247_, _17758_);
  nor (_27280_, _27269_, _27268_);
  and (_27291_, _27280_, _27073_);
  not (_27302_, _17584_);
  nor (_27313_, _26419_, _27302_);
  not (_27324_, _27313_);
  and (_27335_, _26419_, _17758_);
  and (_27346_, _27062_, _15658_);
  not (_27356_, _27346_);
  nor (_27367_, _27356_, _27335_);
  and (_27378_, _27367_, _27324_);
  nor (_27389_, _27378_, _27291_);
  and (_27400_, _26648_, _21044_);
  not (_27411_, _27400_);
  and (_27422_, _18978_, _18815_);
  nor (_27433_, _27422_, _18477_);
  and (_27444_, _27433_, _27400_);
  and (_27455_, _27444_, _18117_);
  nor (_27466_, _27455_, _18520_);
  and (_27476_, _27466_, _16919_);
  nor (_27487_, _27171_, _17758_);
  nor (_27498_, _27487_, _27444_);
  and (_27509_, _27498_, _26419_);
  nor (_27530_, _27509_, _27476_);
  nor (_27531_, _27530_, _17758_);
  and (_27542_, _27530_, _17758_);
  nor (_27552_, _27542_, _27531_);
  nor (_27563_, _27552_, _27411_);
  not (_27574_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27585_, _15680_, _27574_);
  and (_27596_, _27585_, _21023_);
  and (_27607_, _27596_, _25397_);
  and (_27618_, _21044_, _15658_);
  and (_27629_, _27618_, _25375_);
  and (_27640_, _27585_, _26648_);
  not (_27651_, _27640_);
  nor (_27662_, _27651_, _25386_);
  and (_27672_, _25342_, _21044_);
  and (_27683_, _27672_, _17758_);
  or (_27694_, _27683_, _27662_);
  or (_27705_, _27694_, _27629_);
  nor (_27716_, _27705_, _27607_);
  and (_27727_, _27062_, _26648_);
  not (_27738_, _27727_);
  nor (_27749_, _27738_, _26419_);
  and (_27760_, _27585_, _15647_);
  not (_27771_, _27760_);
  nor (_27782_, _27771_, _16919_);
  not (_27793_, _27782_);
  and (_27813_, _21023_, _15691_);
  not (_27814_, _27813_);
  nor (_27825_, _27814_, _17758_);
  and (_27836_, _27062_, _21023_);
  not (_27847_, _27836_);
  nor (_27858_, _27847_, _19360_);
  nor (_27869_, _27858_, _27825_);
  and (_27880_, _27869_, _27793_);
  not (_27891_, _27880_);
  nor (_27902_, _27891_, _27749_);
  and (_27913_, _27902_, _27716_);
  not (_27923_, _27913_);
  nor (_27934_, _27923_, _27563_);
  and (_27945_, _27934_, _27389_);
  not (_27956_, _27945_);
  nor (_27967_, _27956_, _27051_);
  and (_27978_, _27967_, _26626_);
  not (_27989_, _27978_);
  nor (_28000_, _27989_, _25320_);
  and (_28011_, _28000_, _25309_);
  not (_28022_, _28011_);
  or (_28033_, _28022_, _25287_);
  not (_28044_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_28054_, \oc8051_top_1.oc8051_decoder1.wr , _15636_);
  not (_28065_, _28054_);
  nor (_28076_, _28065_, _23932_);
  and (_28087_, _28076_, _28044_);
  not (_28098_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_28109_, _25287_, _28098_);
  and (_28120_, _28109_, _28087_);
  and (_28131_, _28120_, _28033_);
  nor (_28142_, _28076_, _28098_);
  not (_28153_, _26659_);
  nor (_28164_, _27007_, _25386_);
  nor (_28175_, _28164_, _25375_);
  nor (_28185_, _28175_, _28153_);
  not (_28196_, _28185_);
  and (_28207_, _17758_, _27302_);
  nor (_28218_, _28207_, _26583_);
  nor (_28229_, _28218_, _25374_);
  and (_28250_, _26419_, _16919_);
  and (_28251_, _28250_, _27466_);
  nor (_28262_, _28251_, _27335_);
  nor (_28273_, _26419_, _17758_);
  not (_28284_, _28273_);
  nor (_28295_, _28284_, _27476_);
  nor (_28306_, _28295_, _27411_);
  and (_28317_, _28306_, _28262_);
  or (_28327_, _28317_, _27444_);
  nor (_28338_, _27814_, _26419_);
  not (_28349_, _28338_);
  and (_28360_, _26376_, _26354_);
  and (_28371_, _27585_, _25342_);
  and (_28382_, _27618_, _26354_);
  nor (_28393_, _28382_, _28371_);
  nor (_28404_, _28393_, _28360_);
  nor (_28415_, _27738_, _19360_);
  and (_28435_, _27585_, _15658_);
  not (_28436_, _28435_);
  nor (_28447_, _28436_, _17758_);
  nor (_28458_, _28447_, _28415_);
  not (_28469_, _28458_);
  nor (_28480_, _28469_, _28404_);
  and (_28491_, _28480_, _28349_);
  nor (_28502_, _26408_, _26354_);
  not (_28513_, _27596_);
  nor (_28524_, _28513_, _26398_);
  nor (_28535_, _28524_, _27640_);
  nor (_28545_, _28535_, _28502_);
  nor (_28556_, _27672_, _27160_);
  and (_28567_, _27847_, _26408_);
  nor (_28578_, _28567_, _26398_);
  not (_28589_, _28578_);
  nor (_28600_, _28589_, _28556_);
  nor (_28611_, _28600_, _28545_);
  and (_28622_, _28611_, _28491_);
  not (_28633_, _28622_);
  nor (_28644_, _28633_, _28327_);
  not (_28654_, _28644_);
  nor (_28665_, _28654_, _28229_);
  and (_28676_, _28665_, _28196_);
  not (_28687_, _24197_);
  nor (_28698_, _24434_, _24313_);
  and (_28709_, _28698_, _28687_);
  and (_28720_, _28709_, _25277_);
  nand (_28731_, _28720_, _28676_);
  and (_28742_, _28076_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_28753_, _28720_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_28764_, _28753_, _28742_);
  and (_28774_, _28764_, _28731_);
  or (_28785_, _28774_, _28142_);
  or (_28796_, _28785_, _28131_);
  and (_06695_, _28796_, _41806_);
  and (_28817_, _23499_, _21055_);
  not (_28828_, _28817_);
  and (_28839_, _20779_, _15702_);
  and (_28850_, _26419_, _26800_);
  nor (_28861_, _28850_, _26811_);
  not (_28872_, _28861_);
  nor (_28883_, _26659_, _25353_);
  nor (_28893_, _28883_, _28872_);
  not (_28904_, _28893_);
  and (_28915_, _27596_, _26028_);
  not (_28926_, _28915_);
  and (_28937_, _27618_, _26006_);
  not (_28948_, _28937_);
  nor (_28969_, _27651_, _26017_);
  and (_28970_, _27672_, _19360_);
  nor (_28981_, _28970_, _28969_);
  and (_28992_, _28981_, _28948_);
  and (_29002_, _28992_, _28926_);
  nor (_29013_, _28436_, _26419_);
  not (_29024_, _29013_);
  nor (_29035_, _27356_, _16425_);
  and (_29046_, _27073_, _19360_);
  nor (_29057_, _29046_, _29035_);
  and (_29068_, _27062_, _26647_);
  not (_29079_, _29068_);
  nor (_29090_, _29079_, _18815_);
  not (_29101_, _29090_);
  and (_29112_, _28371_, _18215_);
  nor (_29122_, _27813_, _27400_);
  nor (_29133_, _29122_, _19360_);
  nor (_29144_, _29133_, _29112_);
  and (_29155_, _29144_, _29101_);
  and (_29166_, _29155_, _29057_);
  and (_29177_, _29166_, _29024_);
  and (_29188_, _29177_, _29002_);
  and (_29198_, _29188_, _28904_);
  not (_29209_, _29198_);
  nor (_29220_, _29209_, _28839_);
  and (_29231_, _29220_, _28828_);
  not (_29242_, _29231_);
  or (_29253_, _29242_, _25287_);
  not (_29264_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_29275_, _25287_, _29264_);
  and (_29285_, _29275_, _28087_);
  and (_29296_, _29285_, _29253_);
  nor (_29307_, _28076_, _29264_);
  not (_29318_, _28676_);
  or (_29329_, _29318_, _25287_);
  and (_29340_, _29275_, _28742_);
  and (_29351_, _29340_, _29329_);
  or (_29362_, _29351_, _29307_);
  or (_29372_, _29362_, _29296_);
  and (_08932_, _29372_, _41806_);
  and (_29393_, _20811_, _15702_);
  not (_29404_, _29393_);
  and (_29415_, _23564_, _21055_);
  nor (_29426_, _26006_, _25778_);
  or (_29437_, _29426_, _26724_);
  and (_29448_, _29437_, _26811_);
  nor (_29458_, _29437_, _26811_);
  or (_29469_, _29458_, _29448_);
  and (_29480_, _29469_, _26659_);
  nor (_29491_, _26430_, _25995_);
  nor (_29512_, _29491_, _26441_);
  nor (_29513_, _29512_, _25374_);
  not (_29524_, _29513_);
  nor (_29535_, _27433_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_29546_, _29535_, _27400_);
  and (_29556_, _29546_, _27814_);
  or (_29567_, _29556_, _18815_);
  and (_29578_, _27596_, _25778_);
  nor (_29589_, _27651_, _25767_);
  or (_29600_, _29589_, _29578_);
  not (_29611_, _29600_);
  and (_29622_, _27618_, _25756_);
  and (_29633_, _27672_, _18815_);
  nor (_29643_, _29633_, _29622_);
  and (_29654_, _29643_, _29611_);
  nor (_29665_, _29535_, _19022_);
  nand (_29676_, _29665_, _27400_);
  nor (_29687_, _29079_, _18978_);
  nor (_29698_, _27771_, _19360_);
  nor (_29709_, _29698_, _29687_);
  and (_29720_, _29709_, _29676_);
  and (_29730_, _29720_, _29654_);
  and (_29741_, _29730_, _29567_);
  and (_29752_, _29741_, _29524_);
  nor (_29773_, _27356_, _17410_);
  nor (_29774_, _27182_, _27084_);
  not (_29785_, _29774_);
  nor (_29796_, _29785_, _26419_);
  and (_29806_, _29785_, _26419_);
  nor (_29817_, _29806_, _29796_);
  and (_29828_, _29817_, _27073_);
  nor (_29839_, _29828_, _29773_);
  nand (_29850_, _29839_, _29752_);
  nor (_29861_, _29850_, _29480_);
  not (_29872_, _29861_);
  nor (_29883_, _29872_, _29415_);
  and (_29893_, _29883_, _29404_);
  not (_29904_, _29893_);
  or (_29915_, _29904_, _25287_);
  not (_29926_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_29937_, _25287_, _29926_);
  and (_29948_, _29937_, _28087_);
  and (_29959_, _29948_, _29915_);
  nor (_29970_, _28076_, _29926_);
  not (_29980_, _24434_);
  and (_29991_, _29980_, _24313_);
  and (_30002_, _29991_, _24197_);
  and (_30013_, _30002_, _25277_);
  or (_30024_, _30013_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_30035_, _30024_, _28742_);
  nand (_30046_, _30013_, _28676_);
  and (_30057_, _30046_, _30035_);
  or (_30077_, _30057_, _29970_);
  or (_30078_, _30077_, _29959_);
  and (_08943_, _30078_, _41806_);
  and (_30099_, _20842_, _15702_);
  not (_30110_, _30099_);
  and (_30121_, _23629_, _21055_);
  nor (_30132_, _27356_, _16096_);
  and (_30143_, _27084_, _26419_);
  and (_30153_, _27182_, _27160_);
  nor (_30164_, _30153_, _30143_);
  and (_30175_, _30164_, _18978_);
  nor (_30186_, _30164_, _18978_);
  nor (_30197_, _30186_, _30175_);
  and (_30208_, _30197_, _27073_);
  nor (_30219_, _30208_, _30132_);
  nor (_30230_, _26441_, _25963_);
  nor (_30240_, _30230_, _26452_);
  nor (_30251_, _30240_, _25374_);
  not (_30262_, _30251_);
  nor (_30273_, _29079_, _18477_);
  and (_30284_, _27618_, _25723_);
  and (_30295_, _27672_, _18978_);
  nor (_30306_, _30295_, _30284_);
  nor (_30317_, _27651_, _25744_);
  and (_30327_, _27596_, _25745_);
  nor (_30338_, _30327_, _30317_);
  nor (_30349_, _27771_, _18815_);
  nor (_30360_, _27814_, _18978_);
  nor (_30371_, _30360_, _30349_);
  and (_30382_, _30371_, _30338_);
  nand (_30402_, _30382_, _30306_);
  nor (_30403_, _30402_, _30273_);
  and (_30414_, _30403_, _30262_);
  nor (_30425_, _26844_, _26822_);
  nor (_30436_, _30425_, _28153_);
  and (_30447_, _30436_, _26866_);
  and (_30458_, _27422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_30470_, _29665_, _18978_);
  nor (_30491_, _30470_, _30458_);
  nor (_30501_, _30491_, _27411_);
  nor (_30512_, _30501_, _30447_);
  and (_30523_, _30512_, _30414_);
  and (_30534_, _30523_, _30219_);
  not (_30545_, _30534_);
  nor (_30556_, _30545_, _30121_);
  and (_30567_, _30556_, _30110_);
  not (_30578_, _30567_);
  or (_30589_, _30578_, _25287_);
  not (_30599_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_30610_, _25287_, _30599_);
  and (_30621_, _30610_, _28087_);
  and (_30632_, _30621_, _30589_);
  nor (_30643_, _28076_, _30599_);
  nand (_30654_, _25277_, _24197_);
  or (_30665_, _28698_, _30654_);
  and (_30676_, _30665_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_30686_, _24313_);
  and (_30697_, _24197_, _24434_);
  and (_30708_, _30697_, _30686_);
  and (_30719_, _30708_, _29318_);
  and (_30730_, _24197_, _24313_);
  and (_30741_, _30730_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_30752_, _30741_, _30719_);
  and (_30763_, _30752_, _25277_);
  or (_30773_, _30763_, _30676_);
  and (_30784_, _30773_, _28742_);
  or (_30795_, _30784_, _30643_);
  or (_30806_, _30795_, _30632_);
  and (_08954_, _30806_, _41806_);
  and (_30827_, _20885_, _15702_);
  not (_30838_, _30827_);
  and (_30849_, _23694_, _21055_);
  and (_30859_, _26866_, _26789_);
  or (_30870_, _30859_, _28153_);
  nor (_30891_, _30870_, _26877_);
  not (_30892_, _30891_);
  nor (_30903_, _26452_, _25930_);
  nor (_30914_, _30903_, _26463_);
  nor (_30925_, _30914_, _25374_);
  not (_30936_, _30925_);
  nor (_30946_, _27356_, _17094_);
  nor (_30957_, _27193_, _26419_);
  nor (_30968_, _27095_, _27160_);
  nor (_30979_, _30968_, _30957_);
  and (_30990_, _30979_, _18488_);
  not (_31001_, _30990_);
  not (_31012_, _27073_);
  nor (_31022_, _30979_, _18488_);
  nor (_31033_, _31022_, _31012_);
  and (_31044_, _31033_, _31001_);
  nor (_31055_, _31044_, _30946_);
  not (_31066_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_31077_, _27422_, _31066_);
  nor (_31088_, _31077_, _18488_);
  nor (_31099_, _27814_, _18477_);
  nor (_31119_, _27433_, _27411_);
  nor (_31120_, _31119_, _31099_);
  nor (_31131_, _31120_, _31088_);
  not (_31142_, _31131_);
  nor (_31153_, _27651_, _25691_);
  and (_31164_, _27596_, _25713_);
  nor (_31175_, _31164_, _31153_);
  and (_31186_, _27618_, _25702_);
  and (_31197_, _27672_, _18477_);
  nor (_31207_, _31197_, _31186_);
  nor (_31218_, _29079_, _18107_);
  nor (_31229_, _27771_, _18978_);
  nor (_31240_, _31229_, _31218_);
  and (_31251_, _31240_, _31207_);
  and (_31262_, _31251_, _31175_);
  and (_31273_, _31262_, _31142_);
  and (_31284_, _31273_, _31055_);
  and (_31294_, _31284_, _30936_);
  and (_31305_, _31294_, _30892_);
  not (_31316_, _31305_);
  nor (_31327_, _31316_, _30849_);
  and (_31338_, _31327_, _30838_);
  not (_31349_, _31338_);
  or (_31360_, _31349_, _25287_);
  not (_31371_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_31381_, _25287_, _31371_);
  and (_31392_, _31381_, _28087_);
  and (_31403_, _31392_, _31360_);
  nor (_31414_, _28076_, _31371_);
  and (_31425_, _30654_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_31436_, _28698_, _24197_);
  not (_31447_, _31436_);
  nor (_31458_, _31447_, _28676_);
  nor (_31468_, _30730_, _30697_);
  nor (_31479_, _31468_, _31371_);
  or (_31490_, _31479_, _31458_);
  and (_31501_, _31490_, _25277_);
  or (_31512_, _31501_, _31425_);
  and (_31523_, _31512_, _28742_);
  or (_31534_, _31523_, _31414_);
  or (_31545_, _31534_, _31403_);
  and (_08965_, _31545_, _41806_);
  and (_31565_, _23759_, _21055_);
  not (_31576_, _31565_);
  and (_31587_, _20917_, _15702_);
  or (_31598_, _26909_, _25669_);
  nor (_31609_, _28153_, _26920_);
  and (_31620_, _31609_, _31598_);
  nor (_31630_, _26528_, _25669_);
  and (_31641_, _26528_, _25669_);
  nor (_31652_, _31641_, _31630_);
  and (_31663_, _31652_, _25353_);
  and (_31674_, _26419_, _18117_);
  nor (_31695_, _26419_, _16260_);
  or (_31696_, _31695_, _31674_);
  and (_31707_, _31696_, _27346_);
  and (_31717_, _27106_, _26419_);
  and (_31728_, _27204_, _27160_);
  nor (_31739_, _31728_, _31717_);
  nor (_31750_, _31739_, _18107_);
  and (_31761_, _31739_, _18107_);
  or (_31772_, _31761_, _31012_);
  nor (_31783_, _31772_, _31750_);
  nor (_31794_, _31783_, _31707_);
  or (_31804_, _27444_, _18117_);
  nor (_31815_, _27455_, _27411_);
  and (_31826_, _31815_, _31804_);
  and (_31837_, _27596_, _25669_);
  nor (_31848_, _27651_, _25658_);
  not (_31859_, _31848_);
  and (_31870_, _27618_, _25647_);
  and (_31881_, _27672_, _18107_);
  nor (_31891_, _31881_, _31870_);
  nand (_31902_, _31891_, _31859_);
  nor (_31913_, _31902_, _31837_);
  nor (_31924_, _29079_, _17943_);
  nor (_31935_, _27814_, _18107_);
  nor (_31946_, _27771_, _18477_);
  or (_31957_, _31946_, _31935_);
  nor (_31968_, _31957_, _31924_);
  nand (_31979_, _31968_, _31913_);
  nor (_31989_, _31979_, _31826_);
  nand (_32000_, _31989_, _31794_);
  or (_32011_, _32000_, _31663_);
  or (_32022_, _32011_, _31620_);
  nor (_32033_, _32022_, _31587_);
  and (_32044_, _32033_, _31576_);
  not (_32055_, _32044_);
  or (_32065_, _32055_, _25287_);
  not (_32076_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_32087_, _25287_, _32076_);
  and (_32098_, _32087_, _28087_);
  and (_32109_, _32098_, _32065_);
  nor (_32120_, _28076_, _32076_);
  and (_32131_, _24445_, _28687_);
  nor (_32142_, _24445_, _28687_);
  nor (_32152_, _32142_, _32131_);
  not (_32163_, _32152_);
  nand (_32174_, _32163_, _25277_);
  and (_32185_, _32174_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_32196_, _32131_, _29318_);
  and (_32207_, _32142_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_32218_, _32207_, _32196_);
  and (_32229_, _32218_, _25277_);
  or (_32240_, _32229_, _32185_);
  and (_32251_, _32240_, _28742_);
  or (_32262_, _32251_, _32120_);
  or (_32273_, _32262_, _32109_);
  and (_08976_, _32273_, _41806_);
  and (_32294_, _23824_, _21055_);
  not (_32305_, _32294_);
  and (_32326_, _20959_, _15702_);
  nor (_32327_, _26942_, _26920_);
  not (_32338_, _32327_);
  nor (_32349_, _28153_, _26953_);
  and (_32360_, _32349_, _32338_);
  not (_32371_, _32360_);
  nor (_32382_, _26539_, _25636_);
  nor (_32393_, _32382_, _26550_);
  nor (_32404_, _32393_, _25374_);
  nor (_32415_, _26419_, _17247_);
  and (_32425_, _26419_, _18520_);
  nor (_32436_, _32425_, _32415_);
  nor (_32447_, _32436_, _27356_);
  nor (_32458_, _27117_, _27160_);
  nor (_32469_, _27215_, _26419_);
  nor (_32480_, _32469_, _32458_);
  and (_32491_, _32480_, _18520_);
  nor (_32502_, _32480_, _18520_);
  or (_32513_, _32502_, _31012_);
  nor (_32524_, _32513_, _32491_);
  nor (_32535_, _32524_, _32447_);
  not (_32546_, _27509_);
  and (_32557_, _32546_, _27466_);
  nor (_32568_, _27509_, _27455_);
  nor (_32579_, _32568_, _17943_);
  nor (_32590_, _32579_, _32557_);
  nor (_32601_, _32590_, _27411_);
  nor (_32612_, _27651_, _25495_);
  and (_32633_, _27596_, _25506_);
  nor (_32634_, _32633_, _32612_);
  and (_32645_, _27618_, _25484_);
  and (_32656_, _27672_, _17943_);
  nor (_32667_, _32656_, _32645_);
  nor (_32678_, _29079_, _16919_);
  not (_32689_, _32678_);
  nor (_32700_, _27814_, _17943_);
  nor (_32711_, _27771_, _18107_);
  nor (_32722_, _32711_, _32700_);
  and (_32733_, _32722_, _32689_);
  and (_32744_, _32733_, _32667_);
  and (_32755_, _32744_, _32634_);
  not (_32766_, _32755_);
  nor (_32777_, _32766_, _32601_);
  and (_32788_, _32777_, _32535_);
  not (_32798_, _32788_);
  nor (_32809_, _32798_, _32404_);
  and (_32820_, _32809_, _32371_);
  not (_32831_, _32820_);
  nor (_32842_, _32831_, _32326_);
  and (_32853_, _32842_, _32305_);
  not (_32864_, _32853_);
  or (_32875_, _32864_, _25287_);
  not (_32886_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_32897_, _25287_, _32886_);
  and (_32908_, _32897_, _28087_);
  and (_32919_, _32908_, _32875_);
  nor (_32930_, _28076_, _32886_);
  and (_32941_, _29991_, _28687_);
  and (_32952_, _32941_, _25277_);
  nand (_32963_, _32952_, _28676_);
  or (_32984_, _32952_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_32985_, _32984_, _28742_);
  and (_32996_, _32985_, _32963_);
  or (_33007_, _32996_, _32930_);
  or (_33018_, _33007_, _32919_);
  and (_08987_, _33018_, _41806_);
  and (_33039_, _23889_, _21055_);
  not (_33050_, _33039_);
  and (_33061_, _20991_, _15702_);
  nor (_33072_, _26975_, _26953_);
  not (_33083_, _33072_);
  nor (_33094_, _28153_, _26986_);
  and (_33105_, _33094_, _33083_);
  not (_33116_, _33105_);
  nor (_33127_, _26550_, _25604_);
  nor (_33138_, _33127_, _26561_);
  nor (_33148_, _33138_, _25374_);
  nor (_33159_, _26419_, _25408_);
  or (_33170_, _33159_, _27356_);
  nor (_33181_, _33170_, _28250_);
  nor (_33192_, _26419_, _18520_);
  nand (_33203_, _33192_, _27215_);
  nand (_33214_, _27127_, _26419_);
  and (_33225_, _33214_, _33203_);
  nor (_33236_, _33225_, _16919_);
  not (_33247_, _33236_);
  and (_33258_, _33225_, _16919_);
  nor (_33269_, _33258_, _31012_);
  and (_33280_, _33269_, _33247_);
  nor (_33291_, _33280_, _33181_);
  nor (_33302_, _32557_, _16919_);
  and (_33313_, _32557_, _16919_);
  nor (_33324_, _33313_, _33302_);
  nor (_33335_, _33324_, _27411_);
  and (_33356_, _27596_, _25452_);
  nor (_33357_, _27651_, _25441_);
  not (_33368_, _33357_);
  and (_33379_, _27618_, _25430_);
  and (_33390_, _27672_, _16919_);
  nor (_33401_, _33390_, _33379_);
  nand (_33412_, _33401_, _33368_);
  nor (_33423_, _33412_, _33356_);
  nor (_33434_, _29079_, _17758_);
  not (_33445_, _33434_);
  nor (_33456_, _27814_, _16919_);
  nor (_33467_, _27771_, _17943_);
  nor (_33478_, _33467_, _33456_);
  and (_33489_, _33478_, _33445_);
  and (_33499_, _33489_, _33423_);
  not (_33510_, _33499_);
  nor (_33521_, _33510_, _33335_);
  and (_33532_, _33521_, _33291_);
  not (_33543_, _33532_);
  nor (_33554_, _33543_, _33148_);
  and (_33565_, _33554_, _33116_);
  not (_33576_, _33565_);
  nor (_33587_, _33576_, _33061_);
  and (_33598_, _33587_, _33050_);
  not (_33609_, _33598_);
  or (_33620_, _33609_, _25287_);
  not (_33631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_33642_, _25287_, _33631_);
  and (_33653_, _33642_, _28087_);
  and (_33664_, _33653_, _33620_);
  nor (_33675_, _28076_, _33631_);
  nor (_33686_, _24197_, _24313_);
  and (_33697_, _33686_, _24434_);
  and (_33708_, _33697_, _25277_);
  nand (_33719_, _33708_, _28676_);
  or (_33730_, _33708_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_33741_, _33730_, _28742_);
  and (_33752_, _33741_, _33719_);
  or (_33763_, _33752_, _33675_);
  or (_33774_, _33763_, _33664_);
  and (_08998_, _33774_, _41806_);
  and (_33795_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_33806_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_33817_, _33806_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_33828_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_33839_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_33849_, _33839_, _33828_);
  and (_33860_, _33806_, _15636_);
  and (_33881_, _33860_, _33849_);
  not (_33882_, _33881_);
  and (_33893_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_33904_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_33915_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_33926_, _33915_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_33937_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_33948_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_33959_, _33948_, _33937_);
  and (_33970_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not (_33981_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_33992_, _33981_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34003_, _33992_, _33937_);
  and (_34014_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_34025_, _34014_, _33970_);
  and (_34036_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34047_, _34036_, _33937_);
  and (_34058_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not (_34069_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34080_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _34069_);
  and (_34091_, _34080_, _33937_);
  and (_34102_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_34113_, _34102_, _34058_);
  and (_34124_, _33948_, _33937_);
  and (_34135_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_34156_, _33948_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_34157_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_34168_, _34157_, _34135_);
  and (_34179_, _34168_, _34113_);
  and (_34190_, _34179_, _34025_);
  nor (_34200_, _34190_, _33926_);
  nor (_34211_, _34200_, _33904_);
  nor (_34222_, _34211_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34233_, _34222_, _33893_);
  nor (_34244_, _34233_, _33882_);
  and (_34255_, _33849_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_34266_, _34255_, _33882_);
  nor (_34277_, _34266_, _34244_);
  and (_34288_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34299_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_34310_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34321_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_34332_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_34343_, _34332_, _34321_);
  and (_34354_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34365_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_34376_, _34365_, _34354_);
  and (_34387_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_34398_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_34409_, _34398_, _34387_);
  and (_34420_, _34409_, _34376_);
  and (_34431_, _34420_, _34343_);
  nor (_34442_, _34431_, _33915_);
  and (_34453_, _34442_, _34310_);
  nor (_34464_, _34453_, _34299_);
  nor (_34475_, _34464_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34486_, _34475_, _34288_);
  nor (_34497_, _34486_, _33882_);
  and (_34508_, _33849_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_34519_, _34508_, _33882_);
  nor (_34530_, _34519_, _34497_);
  not (_34540_, _34530_);
  and (_34551_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34562_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34573_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_34584_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_34595_, _34584_, _34573_);
  and (_34606_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_34617_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_34628_, _34617_, _34606_);
  and (_34639_, _34628_, _34595_);
  and (_34650_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_34661_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_34672_, _34661_, _34650_);
  and (_34683_, _34672_, _34639_);
  nor (_34694_, _34683_, _33926_);
  nor (_34705_, _34694_, _34562_);
  nor (_34716_, _34705_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34727_, _34716_, _34551_);
  nor (_34738_, _34727_, _33882_);
  and (_34749_, _33849_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_34760_, _34749_, _33882_);
  nor (_34781_, _34760_, _34738_);
  nor (_34782_, _34781_, _34540_);
  and (_34793_, _34782_, _34277_);
  and (_34804_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not (_34815_, _34804_);
  and (_34826_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_34837_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_34848_, _34837_, _34826_);
  and (_34859_, _34848_, _34815_);
  and (_34870_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_34881_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_34891_, _34881_, _34870_);
  and (_34902_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_34913_, _33915_, _34902_);
  and (_34924_, _34913_, _34891_);
  and (_34935_, _34924_, _34859_);
  and (_34946_, _34935_, _34310_);
  nor (_34957_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _34310_);
  nor (_34968_, _34957_, _34946_);
  nor (_34979_, _34968_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_34990_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35001_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _34990_);
  nor (_35012_, _35001_, _34979_);
  and (_35023_, _35012_, _33881_);
  and (_35034_, _33849_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_35045_, _35034_, _33882_);
  nor (_35056_, _35045_, _35023_);
  and (_35067_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35078_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35089_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_35100_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_35111_, _35100_, _35089_);
  and (_35122_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_35133_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_35144_, _35133_, _35122_);
  and (_35155_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_35166_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_35177_, _35166_, _35155_);
  and (_35188_, _35177_, _35144_);
  and (_35199_, _35188_, _35111_);
  nor (_35209_, _35199_, _33926_);
  nor (_35220_, _35209_, _35078_);
  nor (_35231_, _35220_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35242_, _35231_, _35067_);
  nor (_35253_, _35242_, _33882_);
  and (_35264_, _33849_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_35275_, _35264_, _33882_);
  nor (_35286_, _35275_, _35253_);
  nor (_35297_, _35286_, _35056_);
  and (_35308_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35319_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35330_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_35341_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_35352_, _35341_, _35330_);
  and (_35363_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_35374_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_35385_, _35374_, _35363_);
  and (_35396_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_35407_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_35418_, _35407_, _35396_);
  and (_35429_, _35418_, _35385_);
  and (_35440_, _35429_, _35352_);
  nor (_35451_, _35440_, _33915_);
  and (_35462_, _35451_, _34310_);
  or (_35473_, _35462_, _35319_);
  and (_35495_, _35473_, _34990_);
  nor (_35496_, _35495_, _35308_);
  nor (_35518_, _35496_, _33882_);
  and (_35519_, _33849_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_35541_, _35519_, _33882_);
  nor (_35542_, _35541_, _35518_);
  and (_35563_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_35564_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_35575_, _35564_, _35563_);
  and (_35586_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_35597_, _35586_, _33915_);
  and (_35608_, _35597_, _35575_);
  and (_35619_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_35630_, _35619_);
  and (_35641_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_35652_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_35663_, _35652_, _35641_);
  and (_35674_, _35663_, _35630_);
  and (_35685_, _35674_, _35608_);
  and (_35696_, _35685_, _34310_);
  nor (_35707_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _34310_);
  or (_35718_, _35707_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35729_, _35718_, _35696_);
  and (_35740_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_35751_, _35740_, _35729_);
  and (_35762_, _35751_, _33881_);
  and (_35773_, _33849_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_35784_, _35773_, _33882_);
  nor (_35795_, _35784_, _35762_);
  not (_35806_, _35795_);
  and (_35817_, _35806_, _35542_);
  and (_35828_, _35817_, _35297_);
  and (_35839_, _35828_, _34793_);
  and (_35850_, _35297_, _35542_);
  and (_35860_, _34781_, _34277_);
  and (_35871_, _35860_, _34540_);
  and (_35882_, _35871_, _35850_);
  or (_35893_, _35882_, _35839_);
  not (_35904_, _35893_);
  and (_35915_, _35860_, _34530_);
  and (_35926_, _35915_, _35850_);
  not (_35937_, _34277_);
  and (_35948_, _34781_, _35937_);
  and (_35959_, _35948_, _34540_);
  and (_35970_, _35959_, _35828_);
  nor (_35981_, _35970_, _35926_);
  and (_35992_, _35948_, _34530_);
  and (_36003_, _35992_, _35806_);
  and (_36014_, _36003_, _35850_);
  and (_36025_, _34782_, _35937_);
  and (_36036_, _36025_, _35850_);
  nor (_36047_, _36036_, _36014_);
  and (_36058_, _36047_, _35981_);
  and (_36069_, _35795_, _35850_);
  nor (_36080_, _34781_, _34530_);
  and (_36091_, _36080_, _35937_);
  or (_36102_, _36091_, _34793_);
  and (_36113_, _36102_, _36069_);
  and (_36124_, _35992_, _35795_);
  and (_36135_, _36124_, _35850_);
  nor (_36146_, _36135_, _36113_);
  and (_36157_, _36146_, _36058_);
  and (_36167_, _36157_, _35904_);
  and (_36178_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_36189_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_36200_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_36211_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_36222_, _36211_, _36200_);
  and (_36233_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_36244_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_36255_, _36244_, _36233_);
  and (_36266_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_36277_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_36288_, _36277_, _36266_);
  and (_36299_, _36288_, _36255_);
  and (_36310_, _36299_, _36222_);
  nor (_36321_, _36310_, _33915_);
  and (_36332_, _36321_, _34310_);
  nor (_36343_, _36332_, _36189_);
  nor (_36354_, _36343_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_36365_, _36354_, _36178_);
  nor (_36376_, _36365_, _33882_);
  and (_36387_, _33849_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_36398_, _36387_, _33882_);
  nor (_36409_, _36398_, _36376_);
  not (_36420_, _36409_);
  not (_36431_, _35056_);
  and (_36442_, _35542_, _35286_);
  and (_36453_, _36442_, _36431_);
  and (_36464_, _36453_, _36420_);
  and (_36474_, _35959_, _35795_);
  and (_36485_, _36474_, _36464_);
  and (_36496_, _36464_, _36003_);
  and (_36507_, _36080_, _34277_);
  and (_36518_, _36507_, _35806_);
  and (_36529_, _36518_, _36464_);
  nor (_36540_, _36529_, _36496_);
  not (_36551_, _36540_);
  nor (_36562_, _36551_, _36485_);
  and (_36573_, _36409_, _35056_);
  and (_36584_, _36573_, _36442_);
  and (_36595_, _36025_, _35806_);
  and (_36606_, _36595_, _36584_);
  not (_36617_, _36606_);
  and (_36628_, _36453_, _36409_);
  and (_36639_, _36628_, _35871_);
  and (_36650_, _36507_, _35795_);
  and (_36661_, _36650_, _35850_);
  nor (_36672_, _36661_, _36639_);
  and (_36683_, _36672_, _36617_);
  and (_36694_, _36683_, _36562_);
  and (_36705_, _36694_, _36167_);
  nor (_36716_, _36705_, _33817_);
  not (_36727_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_36738_, _15636_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_36749_, _36738_, _36727_);
  and (_36760_, _36749_, _36507_);
  and (_36771_, _36760_, _36584_);
  and (_36781_, _36639_, _36738_);
  and (_36792_, _36781_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_36803_, _36792_, _36771_);
  nor (_36814_, _36803_, _36716_);
  nor (_36825_, _36814_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36836_, _36825_, _33795_);
  and (_36847_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_36858_, _33817_);
  not (_36869_, _35286_);
  and (_36880_, _35542_, _36869_);
  nor (_36891_, _36409_, _36431_);
  and (_36902_, _36891_, _36880_);
  and (_36913_, _35948_, _35806_);
  and (_36924_, _36913_, _36902_);
  and (_36935_, _36091_, _35795_);
  and (_36946_, _36935_, _36902_);
  and (_36957_, _35959_, _36069_);
  or (_36968_, _36957_, _36946_);
  or (_36979_, _36968_, _36924_);
  and (_36990_, _34793_, _35806_);
  or (_37001_, _36990_, _35871_);
  and (_37012_, _36902_, _37001_);
  nor (_37023_, _35806_, _35542_);
  and (_37034_, _37023_, _35959_);
  and (_37045_, _35915_, _35795_);
  and (_37056_, _37045_, _36902_);
  or (_37067_, _37056_, _37034_);
  or (_37078_, _37067_, _36639_);
  or (_37087_, _37078_, _37012_);
  and (_37095_, _36902_, _36650_);
  and (_37102_, _36025_, _35795_);
  and (_37110_, _37102_, _36902_);
  or (_37118_, _37110_, _37095_);
  and (_37125_, _36628_, _36474_);
  and (_37133_, _36628_, _36595_);
  nor (_37141_, _37133_, _37125_);
  not (_37148_, _37141_);
  or (_37149_, _37148_, _37118_);
  or (_37150_, _37149_, _37087_);
  or (_37153_, _37150_, _36979_);
  and (_37164_, _34793_, _35795_);
  and (_37175_, _37164_, _36453_);
  and (_37186_, _35915_, _35806_);
  and (_37197_, _37186_, _36902_);
  and (_37208_, _35959_, _35806_);
  and (_37219_, _36584_, _37208_);
  or (_37230_, _37219_, _37197_);
  nor (_37241_, _37230_, _37175_);
  and (_37252_, _36628_, _36518_);
  and (_37263_, _36902_, _36595_);
  nor (_37274_, _37263_, _37252_);
  and (_37285_, _37274_, _37241_);
  and (_37296_, _36584_, _36474_);
  and (_37307_, _37164_, _36902_);
  nor (_37318_, _37307_, _37296_);
  and (_37329_, _36628_, _37208_);
  and (_37340_, _37102_, _36628_);
  nor (_37351_, _37340_, _37329_);
  and (_37362_, _37351_, _37318_);
  and (_37373_, _37362_, _37285_);
  and (_37384_, _36628_, _36003_);
  and (_37394_, _36902_, _36124_);
  or (_37405_, _37394_, _37384_);
  and (_37416_, _36584_, _36025_);
  and (_37421_, _36650_, _36453_);
  or (_37432_, _37421_, _37416_);
  or (_37443_, _37432_, _37405_);
  and (_37454_, _36628_, _36124_);
  and (_37464_, _36453_, _36990_);
  or (_37475_, _37464_, _37454_);
  and (_37485_, _36584_, _35871_);
  and (_37496_, _37485_, _35795_);
  and (_37507_, _35806_, _35871_);
  or (_37518_, _37186_, _37507_);
  and (_37528_, _37518_, _36584_);
  nor (_37539_, _37528_, _37496_);
  not (_37550_, _37539_);
  or (_37560_, _37550_, _37475_);
  nor (_37571_, _37560_, _37443_);
  nand (_37582_, _37571_, _37373_);
  or (_37592_, _37582_, _37153_);
  and (_37603_, _37592_, _36858_);
  and (_37614_, _36738_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_37624_, _37614_, _36639_);
  not (_37635_, _37624_);
  nor (_37646_, _34781_, _35937_);
  and (_37657_, _36584_, _37646_);
  and (_37668_, _37657_, _36749_);
  not (_37679_, _36749_);
  and (_37690_, _35795_, _35871_);
  and (_37701_, _37690_, _36584_);
  and (_37712_, _37186_, _36584_);
  nor (_37723_, _37712_, _37701_);
  nor (_37734_, _37723_, _37679_);
  nor (_37745_, _37734_, _37668_);
  and (_37756_, _37745_, _37635_);
  not (_37767_, _37756_);
  nor (_37778_, _37767_, _37603_);
  nor (_37789_, _37778_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37800_, _37789_, _36847_);
  nor (_37811_, _37800_, _36836_);
  and (_37822_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_37833_, _36573_, _36880_);
  and (_37844_, _37833_, _36124_);
  and (_37855_, _37833_, _36474_);
  nor (_37866_, _37855_, _37844_);
  and (_37877_, _37866_, _36562_);
  nor (_37888_, _37877_, _33817_);
  nor (_37899_, _37888_, _37668_);
  nor (_37910_, _37866_, _36858_);
  not (_37921_, _37910_);
  and (_37932_, _37921_, _37899_);
  nor (_37943_, _37932_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37954_, _37943_, _37822_);
  and (_37965_, _37954_, _41806_);
  and (_09544_, _37965_, _37811_);
  and (_37986_, _24796_, _24665_);
  and (_37997_, _37986_, _25244_);
  and (_38008_, _37997_, _24960_);
  and (_38019_, _38008_, _25112_);
  and (_38030_, _38019_, _30002_);
  and (_38041_, _38030_, _28076_);
  and (_38052_, _38041_, _28044_);
  nor (_38063_, _21055_, _15702_);
  and (_38074_, _26648_, _21034_);
  nor (_38085_, _27813_, _38074_);
  and (_38096_, _38085_, _27771_);
  and (_38107_, _38096_, _38063_);
  and (_38118_, _38107_, _29079_);
  nor (_38129_, _38118_, _17758_);
  not (_38140_, _38129_);
  and (_38151_, _38140_, _27716_);
  and (_38162_, _38151_, _27389_);
  not (_38173_, _38162_);
  and (_38183_, _38173_, _38052_);
  and (_38194_, _38019_, _24197_);
  and (_38205_, _38194_, _29991_);
  and (_38216_, _38205_, _28087_);
  not (_38226_, _38216_);
  and (_38237_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_38248_, _38118_, _16919_);
  not (_38258_, _38248_);
  and (_38269_, _38258_, _33423_);
  and (_38280_, _38269_, _33291_);
  nor (_38290_, _38280_, _38226_);
  nor (_38301_, _38290_, _38237_);
  and (_38312_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38322_, _38118_, _17943_);
  not (_38333_, _38322_);
  and (_38344_, _38333_, _32667_);
  and (_38355_, _38344_, _32634_);
  and (_38366_, _38355_, _32535_);
  nor (_38377_, _38366_, _38226_);
  nor (_38388_, _38377_, _38312_);
  and (_38390_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38391_, _38118_, _18107_);
  not (_38392_, _38391_);
  and (_38393_, _38392_, _31913_);
  and (_38394_, _38393_, _31794_);
  nor (_38395_, _38394_, _38226_);
  nor (_38396_, _38395_, _38390_);
  and (_38397_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38398_, _38118_, _18477_);
  not (_38399_, _38398_);
  and (_38400_, _38399_, _31207_);
  and (_38401_, _38400_, _31175_);
  and (_38402_, _38401_, _31055_);
  nor (_38403_, _38402_, _38226_);
  nor (_38404_, _38403_, _38397_);
  and (_38405_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38406_, _38118_, _18978_);
  not (_38407_, _38406_);
  and (_38408_, _38407_, _30306_);
  and (_38409_, _38408_, _30338_);
  and (_38410_, _38409_, _30219_);
  nor (_38411_, _38410_, _38226_);
  nor (_38412_, _38411_, _38405_);
  and (_38413_, _38226_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38414_, _38118_, _18815_);
  not (_38415_, _38414_);
  and (_38416_, _38415_, _29654_);
  and (_38417_, _38416_, _29839_);
  not (_38418_, _38417_);
  and (_38419_, _38418_, _38216_);
  nor (_38420_, _38419_, _38413_);
  nor (_38421_, _38216_, _24379_);
  nor (_38422_, _38118_, _19360_);
  not (_38423_, _38422_);
  and (_38424_, _38423_, _29057_);
  and (_38425_, _38424_, _29002_);
  not (_38426_, _38425_);
  and (_38427_, _38426_, _38216_);
  nor (_38428_, _38427_, _38421_);
  and (_38429_, _38428_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38430_, _38429_, _38420_);
  and (_38431_, _38430_, _38412_);
  and (_38432_, _38431_, _38404_);
  and (_38433_, _38432_, _38396_);
  and (_38434_, _38433_, _38388_);
  and (_38435_, _38434_, _38301_);
  nor (_38436_, _38216_, _24818_);
  and (_38437_, _38436_, _38435_);
  nor (_38438_, _38436_, _38435_);
  nor (_38439_, _38438_, _38437_);
  and (_38440_, _38439_, _24522_);
  nor (_38441_, _38440_, _24862_);
  nor (_38442_, _38441_, _38216_);
  nor (_38443_, _38442_, _38183_);
  nor (_09564_, _38443_, rst);
  not (_38444_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38445_, _38428_, _38444_);
  nor (_38446_, _38428_, _38444_);
  nor (_38447_, _38446_, _38445_);
  and (_38448_, _38447_, _24522_);
  nor (_38449_, _38448_, _24390_);
  nor (_38450_, _38449_, _38216_);
  nor (_38451_, _38450_, _38427_);
  nand (_10690_, _38451_, _41806_);
  nor (_38452_, _38429_, _38420_);
  nor (_38453_, _38452_, _38430_);
  nor (_38454_, _38453_, _23943_);
  nor (_38455_, _38454_, _24245_);
  nor (_38456_, _38455_, _38216_);
  nor (_38457_, _38456_, _38419_);
  nand (_10701_, _38457_, _41806_);
  nor (_38458_, _38430_, _38412_);
  nor (_38459_, _38458_, _38431_);
  nor (_38460_, _38459_, _23943_);
  nor (_38461_, _38460_, _23998_);
  nor (_38462_, _38461_, _38216_);
  nor (_38463_, _38462_, _38411_);
  nand (_10712_, _38463_, _41806_);
  nor (_38464_, _38431_, _38404_);
  nor (_38465_, _38464_, _38432_);
  nor (_38466_, _38465_, _23943_);
  nor (_38467_, _38466_, _25004_);
  nor (_38468_, _38467_, _38216_);
  nor (_38469_, _38468_, _38403_);
  nor (_10723_, _38469_, rst);
  nor (_38470_, _38432_, _38396_);
  nor (_38471_, _38470_, _38433_);
  nor (_38472_, _38471_, _23943_);
  nor (_38473_, _38472_, _25156_);
  nor (_38474_, _38473_, _38216_);
  nor (_38475_, _38474_, _38395_);
  nor (_10734_, _38475_, rst);
  nor (_38476_, _38433_, _38388_);
  nor (_38477_, _38476_, _38434_);
  nor (_38478_, _38477_, _23943_);
  nor (_38479_, _38478_, _24708_);
  nor (_38480_, _38479_, _38216_);
  nor (_38481_, _38480_, _38377_);
  nor (_10745_, _38481_, rst);
  nor (_38482_, _38434_, _38301_);
  nor (_38483_, _38482_, _38435_);
  nor (_38484_, _38483_, _23943_);
  nor (_38485_, _38484_, _24555_);
  nor (_38486_, _38485_, _38216_);
  nor (_38487_, _38486_, _38290_);
  nor (_10756_, _38487_, rst);
  and (_38488_, _28087_, _25112_);
  and (_38489_, _38488_, _31436_);
  nand (_38490_, _38489_, _38008_);
  nor (_38491_, _38490_, _28011_);
  and (_38492_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15636_);
  and (_38493_, _38492_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38494_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38495_, _38494_, _38493_);
  or (_38496_, _38495_, _38491_);
  nor (_38497_, _27814_, _17584_);
  nor (_38498_, _28436_, _18477_);
  and (_38499_, _26419_, _17247_);
  not (_38500_, _38499_);
  nor (_38501_, _17758_, _16425_);
  and (_38502_, _38501_, _27138_);
  and (_38503_, _38502_, _25821_);
  and (_38504_, _38503_, _25865_);
  and (_38505_, _38504_, _26474_);
  nor (_38506_, _38505_, _27160_);
  and (_38507_, _26419_, _16260_);
  nor (_38508_, _38507_, _38506_);
  and (_38509_, _38508_, _38500_);
  and (_38510_, _27226_, _17758_);
  and (_38511_, _17094_, _16096_);
  and (_38512_, _17410_, _16425_);
  and (_38513_, _38512_, _38511_);
  and (_38514_, _38513_, _38510_);
  and (_38515_, _17247_, _16260_);
  and (_38516_, _38515_, _38514_);
  nor (_38517_, _38516_, _26419_);
  not (_38518_, _38517_);
  and (_38519_, _38518_, _38509_);
  nor (_38520_, _26419_, _16601_);
  and (_38521_, _26419_, _16601_);
  nor (_38522_, _38521_, _38520_);
  and (_38523_, _38522_, _38519_);
  nor (_38524_, _38523_, _27302_);
  and (_38525_, _38523_, _27302_);
  nor (_38526_, _38525_, _38524_);
  and (_38527_, _38526_, _27073_);
  and (_38528_, _26419_, _27302_);
  nor (_38529_, _38528_, _28273_);
  nor (_38530_, _38529_, _27356_);
  or (_38531_, _38530_, _38527_);
  or (_38532_, _38531_, _38498_);
  and (_38533_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_38534_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38535_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38536_, _38535_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38537_, _38536_, _38534_);
  nor (_38538_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38539_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38540_, _38539_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38541_, _38540_, _38538_);
  nor (_38542_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38543_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38544_, _38543_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38545_, _38544_, _38542_);
  not (_38546_, _38545_);
  nor (_38547_, _38546_, _28175_);
  nor (_38548_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38549_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38550_, _38549_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38551_, _38550_, _38548_);
  and (_38552_, _38551_, _38547_);
  nor (_38553_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38554_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38555_, _38554_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38556_, _38555_, _38553_);
  and (_38557_, _38556_, _38552_);
  and (_38558_, _38557_, _38541_);
  nor (_38559_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38560_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38561_, _38560_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38562_, _38561_, _38559_);
  and (_38563_, _38562_, _38558_);
  and (_38564_, _38563_, _38537_);
  nor (_38565_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38566_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38567_, _38566_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38568_, _38567_, _38565_);
  and (_38569_, _38568_, _38564_);
  nor (_38570_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38571_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38572_, _38571_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38573_, _38572_, _38570_);
  nor (_38574_, _38573_, _38569_);
  and (_38575_, _38573_, _38569_);
  or (_38576_, _38575_, _38574_);
  nor (_38577_, _38576_, _28153_);
  and (_38578_, _20747_, _15702_);
  or (_38579_, _38578_, _38577_);
  or (_38580_, _38579_, _38533_);
  or (_38581_, _38580_, _38532_);
  nor (_38582_, _38581_, _38497_);
  nand (_38583_, _38582_, _38493_);
  and (_38584_, _38583_, _41806_);
  and (_12702_, _38584_, _38496_);
  and (_38585_, _38488_, _30708_);
  and (_38586_, _38585_, _38008_);
  nor (_38587_, _38586_, _38493_);
  not (_38588_, _38587_);
  nand (_38589_, _38588_, _28011_);
  not (_38590_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_38591_, _38587_, _38590_);
  and (_38592_, _38591_, _41806_);
  and (_12723_, _38592_, _38589_);
  nor (_38593_, _38490_, _29231_);
  and (_38594_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38595_, _38594_, _38493_);
  or (_38596_, _38595_, _38593_);
  nor (_38597_, _27814_, _16425_);
  nor (_38598_, _28436_, _18107_);
  nor (_38599_, _27356_, _19360_);
  nor (_38600_, _28273_, _27335_);
  not (_38601_, _38600_);
  nor (_38602_, _38601_, _27247_);
  nor (_38603_, _38602_, _25789_);
  and (_38604_, _38602_, _25789_);
  nor (_38605_, _38604_, _38603_);
  and (_38606_, _38605_, _27073_);
  or (_38607_, _38606_, _38599_);
  or (_38608_, _38607_, _38598_);
  and (_38609_, _23373_, _21055_);
  and (_38610_, _38546_, _28175_);
  nor (_38611_, _38610_, _38547_);
  and (_38612_, _38611_, _26659_);
  and (_38613_, _20525_, _15702_);
  or (_38614_, _38613_, _38612_);
  or (_38615_, _38614_, _38609_);
  or (_38616_, _38615_, _38608_);
  nor (_38617_, _38616_, _38597_);
  nand (_38618_, _38617_, _38493_);
  and (_38619_, _38618_, _41806_);
  and (_13612_, _38619_, _38596_);
  nor (_38620_, _38490_, _29893_);
  and (_38621_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38622_, _38621_, _38493_);
  or (_38623_, _38622_, _38620_);
  nor (_38624_, _27814_, _17410_);
  nor (_38625_, _28436_, _17943_);
  and (_38626_, _38502_, _26419_);
  and (_38627_, _38510_, _16425_);
  and (_38628_, _38627_, _27160_);
  nor (_38629_, _38628_, _38626_);
  and (_38630_, _38629_, _17410_);
  nor (_38631_, _38629_, _17410_);
  or (_38632_, _38631_, _31012_);
  nor (_38633_, _38632_, _38630_);
  nor (_38634_, _27356_, _18815_);
  or (_38635_, _38634_, _38633_);
  or (_38636_, _38635_, _38625_);
  and (_38637_, _22369_, _21055_);
  nor (_38638_, _38551_, _38547_);
  nor (_38639_, _38638_, _38552_);
  and (_38640_, _38639_, _26659_);
  and (_38641_, _20557_, _15702_);
  or (_38642_, _38641_, _38640_);
  or (_38643_, _38642_, _38637_);
  or (_38644_, _38643_, _38636_);
  nor (_38645_, _38644_, _38624_);
  nand (_38646_, _38645_, _38493_);
  and (_38647_, _38646_, _41806_);
  and (_13621_, _38647_, _38623_);
  nor (_38648_, _38490_, _30567_);
  and (_38649_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38650_, _38649_, _38493_);
  or (_38651_, _38650_, _38648_);
  nor (_38652_, _27814_, _16096_);
  nor (_38653_, _28436_, _16919_);
  and (_38654_, _38627_, _17410_);
  and (_38655_, _38654_, _27160_);
  and (_38656_, _38503_, _26419_);
  nor (_38657_, _38656_, _38655_);
  and (_38658_, _38657_, _16096_);
  nor (_38659_, _38657_, _16096_);
  nor (_38660_, _38659_, _38658_);
  and (_38661_, _38660_, _27073_);
  nor (_38662_, _27356_, _18978_);
  or (_38663_, _38662_, _38661_);
  or (_38664_, _38663_, _38653_);
  and (_38665_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38666_, _38556_, _38552_);
  nor (_38667_, _38666_, _38557_);
  and (_38668_, _38667_, _26659_);
  and (_38669_, _20589_, _15702_);
  or (_38670_, _38669_, _38668_);
  or (_38671_, _38670_, _38665_);
  or (_38672_, _38671_, _38664_);
  nor (_38673_, _38672_, _38652_);
  nand (_38674_, _38673_, _38493_);
  and (_38675_, _38674_, _41806_);
  and (_13631_, _38675_, _38651_);
  nor (_38676_, _38490_, _31338_);
  and (_38677_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38678_, _38677_, _38493_);
  or (_38679_, _38678_, _38676_);
  nor (_38680_, _27814_, _17094_);
  nor (_38681_, _38504_, _26474_);
  not (_38682_, _38681_);
  and (_38683_, _38682_, _38506_);
  and (_38684_, _38654_, _16096_);
  nor (_38685_, _38684_, _17094_);
  nor (_38686_, _38685_, _38514_);
  nor (_38687_, _38686_, _26419_);
  nor (_38688_, _38687_, _38683_);
  nor (_38689_, _38688_, _31012_);
  nor (_38690_, _27356_, _18477_);
  or (_38691_, _38690_, _38689_);
  or (_38692_, _38691_, _28447_);
  and (_38693_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_38694_, _38557_, _38541_);
  not (_38695_, _38694_);
  nor (_38696_, _38558_, _28153_);
  and (_38697_, _38696_, _38695_);
  and (_38698_, _20620_, _15702_);
  or (_38699_, _38698_, _38697_);
  or (_38700_, _38699_, _38693_);
  or (_38701_, _38700_, _38692_);
  nor (_38702_, _38701_, _38680_);
  nand (_38703_, _38702_, _38493_);
  and (_38704_, _38703_, _41806_);
  and (_13640_, _38704_, _38679_);
  nor (_38705_, _38490_, _32044_);
  and (_38706_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38707_, _38706_, _38493_);
  or (_38708_, _38707_, _38705_);
  nor (_38709_, _27814_, _16260_);
  nor (_38710_, _28436_, _19360_);
  nor (_38711_, _38514_, _26419_);
  nor (_38712_, _38711_, _38506_);
  nor (_38713_, _38712_, _25517_);
  and (_38714_, _38712_, _25517_);
  nor (_38715_, _38714_, _38713_);
  and (_38716_, _38715_, _27073_);
  nor (_38717_, _26419_, _18117_);
  or (_38718_, _38717_, _27356_);
  nor (_38719_, _38718_, _38507_);
  or (_38720_, _38719_, _38716_);
  or (_38721_, _38720_, _38710_);
  and (_38722_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38723_, _38562_, _38558_);
  not (_38724_, _38723_);
  nor (_38725_, _38563_, _28153_);
  and (_38726_, _38725_, _38724_);
  and (_38727_, _20652_, _15702_);
  or (_38728_, _38727_, _38726_);
  or (_38729_, _38728_, _38722_);
  or (_38730_, _38729_, _38721_);
  nor (_38731_, _38730_, _38709_);
  nand (_38732_, _38731_, _38493_);
  and (_38733_, _38732_, _41806_);
  and (_13650_, _38733_, _38708_);
  nor (_38734_, _38490_, _32853_);
  and (_38735_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38736_, _38735_, _38493_);
  or (_38737_, _38736_, _38734_);
  nor (_38738_, _27814_, _17247_);
  nor (_38739_, _28436_, _18815_);
  and (_38740_, _38514_, _16260_);
  nor (_38741_, _38740_, _26419_);
  not (_38742_, _38741_);
  and (_38743_, _38742_, _38508_);
  and (_38744_, _38743_, _17247_);
  nor (_38745_, _38743_, _17247_);
  or (_38746_, _38745_, _38744_);
  and (_38747_, _38746_, _27073_);
  nor (_38748_, _33192_, _27356_);
  and (_38749_, _38748_, _38500_);
  or (_38750_, _38749_, _38747_);
  or (_38751_, _38750_, _38739_);
  and (_38752_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_38753_, _38563_, _38537_);
  nor (_38754_, _38753_, _38564_);
  and (_38755_, _38754_, _26659_);
  and (_38756_, _20684_, _15702_);
  or (_38757_, _38756_, _38755_);
  or (_38758_, _38757_, _38752_);
  or (_38759_, _38758_, _38751_);
  nor (_38760_, _38759_, _38738_);
  nand (_38761_, _38760_, _38493_);
  and (_38762_, _38761_, _41806_);
  and (_13660_, _38762_, _38737_);
  nor (_38763_, _38490_, _33598_);
  and (_38764_, _38490_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38765_, _38764_, _38493_);
  or (_38766_, _38765_, _38763_);
  nor (_38767_, _27814_, _16601_);
  nor (_38768_, _28436_, _18978_);
  and (_38769_, _38519_, _16601_);
  nor (_38770_, _38519_, _16601_);
  nor (_38771_, _38770_, _38769_);
  nor (_38772_, _38771_, _31012_);
  nor (_38773_, _26419_, _16930_);
  or (_38774_, _38773_, _27356_);
  nor (_38775_, _38774_, _38521_);
  or (_38776_, _38775_, _38772_);
  or (_38777_, _38776_, _38768_);
  and (_38778_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_38779_, _38568_, _38564_);
  not (_38780_, _38779_);
  nor (_38781_, _38569_, _28153_);
  and (_38782_, _38781_, _38780_);
  and (_38783_, _20715_, _15702_);
  or (_38784_, _38783_, _38782_);
  or (_38785_, _38784_, _38778_);
  or (_38786_, _38785_, _38777_);
  nor (_38787_, _38786_, _38767_);
  nand (_38788_, _38787_, _38493_);
  and (_38789_, _38788_, _41806_);
  and (_13670_, _38789_, _38766_);
  nand (_38790_, _38588_, _29231_);
  not (_38791_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_38792_, _38587_, _38791_);
  and (_38793_, _38792_, _41806_);
  and (_13679_, _38793_, _38790_);
  nand (_38794_, _38588_, _29893_);
  not (_38795_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand (_38796_, _38587_, _38795_);
  and (_38797_, _38796_, _41806_);
  and (_13688_, _38797_, _38794_);
  nand (_38798_, _38588_, _30567_);
  not (_38799_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_38800_, _38587_, _38799_);
  and (_38801_, _38800_, _41806_);
  and (_13698_, _38801_, _38798_);
  nand (_38802_, _38588_, _31338_);
  or (_38803_, _38588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38804_, _38803_, _41806_);
  and (_13708_, _38804_, _38802_);
  nand (_38805_, _38588_, _32044_);
  or (_38806_, _38588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38807_, _38806_, _41806_);
  and (_13718_, _38807_, _38805_);
  nand (_38808_, _38588_, _32853_);
  or (_38809_, _38588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38810_, _38809_, _41806_);
  and (_13727_, _38810_, _38808_);
  nand (_38812_, _38588_, _33598_);
  or (_38815_, _38588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38816_, _38815_, _41806_);
  and (_13736_, _38816_, _38812_);
  and (_38817_, _28087_, _24456_);
  nor (_38818_, _24665_, _24949_);
  and (_38819_, _25255_, _24796_);
  and (_38820_, _38819_, _38818_);
  and (_38821_, _38820_, _38817_);
  nor (_38822_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_38823_, _38822_);
  and (_38824_, _38823_, _28676_);
  and (_38833_, _38820_, _28742_);
  not (_38839_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_38845_, _38822_, _38839_);
  nor (_38849_, _38845_, _38833_);
  not (_38850_, _38849_);
  nor (_38851_, _38850_, _38824_);
  not (_38852_, _38833_);
  not (_38853_, _28709_);
  nor (_38854_, _38853_, _28676_);
  nor (_38855_, _28709_, _38839_);
  nor (_38856_, _38855_, _38854_);
  nor (_38857_, _38856_, _38852_);
  nor (_38858_, _38857_, _38851_);
  or (_38859_, _38858_, _38821_);
  not (_38860_, _38821_);
  or (_38861_, _38860_, _38162_);
  and (_38862_, _38861_, _38859_);
  nor (_16545_, _38862_, rst);
  nor (_38863_, _38860_, _38417_);
  not (_38864_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_38865_, _38833_, _30002_);
  nand (_38866_, _38865_, _38864_);
  and (_38867_, _38866_, _38860_);
  or (_38868_, _38865_, _29318_);
  and (_38869_, _38868_, _38867_);
  or (_38870_, _38869_, _38863_);
  and (_21479_, _38870_, _41806_);
  nand (_38871_, _38821_, _38410_);
  or (_38873_, _20811_, _20779_);
  or (_38875_, _38873_, _20842_);
  or (_38876_, _38875_, _20885_);
  or (_38877_, _38876_, _20959_);
  or (_38878_, _38877_, _20991_);
  or (_38879_, _38878_, _20451_);
  and (_38880_, _38879_, _15702_);
  or (_38881_, _28218_, _26572_);
  not (_38882_, _28207_);
  nand (_38883_, _38882_, _26572_);
  and (_38884_, _38883_, _25353_);
  and (_38885_, _38884_, _38881_);
  not (_38886_, _25375_);
  nand (_38887_, _27007_, _38886_);
  nor (_38888_, _28153_, _28164_);
  and (_38889_, _38888_, _38887_);
  and (_38890_, _38515_, _22269_);
  and (_38891_, _38513_, _21055_);
  nand (_38892_, _38891_, _38890_);
  nand (_38893_, _38892_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_38894_, _38893_, _38889_);
  or (_38895_, _38894_, _38885_);
  or (_38896_, _38895_, _31587_);
  or (_38897_, _38896_, _38880_);
  nor (_38898_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_38899_, _38898_, _38833_);
  and (_38900_, _38899_, _38897_);
  not (_38901_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_38902_, _30708_, _38901_);
  or (_38903_, _38902_, _30719_);
  and (_38904_, _38903_, _38833_);
  or (_38905_, _38904_, _38821_);
  or (_38906_, _38905_, _38900_);
  and (_38907_, _38906_, _38871_);
  and (_21490_, _38907_, _41806_);
  nor (_38908_, _38860_, _38402_);
  and (_38909_, _38833_, _31436_);
  and (_38910_, _38909_, _28676_);
  nor (_38912_, _38909_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_38915_, _38912_, _38821_);
  not (_38921_, _38915_);
  nor (_38926_, _38921_, _38910_);
  nor (_38933_, _38926_, _38908_);
  nor (_21502_, _38933_, rst);
  not (_38949_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  not (_38950_, _24665_);
  nand (_38951_, _38819_, _38950_);
  not (_38952_, _28742_);
  nor (_38953_, _38952_, _24949_);
  not (_38954_, _38953_);
  nor (_38955_, _38954_, _38951_);
  and (_38956_, _38955_, _32163_);
  nor (_38957_, _38956_, _38949_);
  and (_38958_, _32142_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_38959_, _38958_, _32196_);
  nor (_38960_, _38959_, _38852_);
  nor (_38961_, _38960_, _38957_);
  nor (_38962_, _38961_, _38821_);
  nor (_38963_, _38860_, _38394_);
  nor (_38964_, _38963_, _38962_);
  nor (_21514_, _38964_, rst);
  nand (_38965_, _38833_, _32941_);
  nor (_38966_, _38965_, _28676_);
  and (_38967_, _38965_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_38968_, _38967_, _38821_);
  or (_38969_, _38968_, _38966_);
  nand (_38970_, _38821_, _38366_);
  and (_38971_, _38970_, _38969_);
  and (_21526_, _38971_, _41806_);
  and (_38972_, _33697_, _29318_);
  nor (_38973_, _33697_, _31066_);
  nor (_38974_, _38973_, _38972_);
  nor (_38975_, _38974_, _38852_);
  and (_38976_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_38977_, _38976_);
  nor (_38978_, _38977_, _27813_);
  nor (_38979_, _38978_, _31066_);
  and (_38980_, _26659_, _26909_);
  and (_38981_, _26528_, _25353_);
  nor (_38982_, _38981_, _38980_);
  nor (_38983_, _38982_, _38977_);
  nor (_38984_, _38983_, _38979_);
  nor (_38988_, _38984_, _38833_);
  nor (_38999_, _38988_, _38975_);
  nor (_39002_, _38999_, _38821_);
  nor (_39003_, _38860_, _38280_);
  nor (_39004_, _39003_, _39002_);
  nor (_21538_, _39004_, rst);
  not (_39020_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39021_, _38492_, _39020_);
  not (_39022_, _39021_);
  or (_39023_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_39024_, _39023_, _39020_);
  and (_39025_, _24197_, _25112_);
  and (_39026_, _39025_, _24445_);
  not (_39027_, _24796_);
  and (_39028_, _25244_, _39027_);
  and (_39029_, _39028_, _28087_);
  and (_39030_, _39029_, _39026_);
  nand (_39031_, _39030_, _38818_);
  and (_39032_, _39031_, _39024_);
  nor (_39033_, _39032_, _28011_);
  and (_39034_, _25244_, _25112_);
  and (_39035_, _39034_, _24807_);
  and (_39036_, _39035_, _38953_);
  and (_39037_, _39036_, _28709_);
  and (_39038_, _39037_, _28676_);
  nor (_39039_, _39037_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_39040_, _39039_);
  and (_39041_, _39032_, _39022_);
  and (_39042_, _39041_, _39040_);
  not (_39043_, _39042_);
  nor (_39044_, _39043_, _39038_);
  or (_39045_, _39044_, _39033_);
  and (_39046_, _39045_, _39022_);
  nor (_39047_, _39022_, _38582_);
  or (_39048_, _39047_, _39046_);
  and (_22313_, _39048_, _41806_);
  nor (_39049_, _39032_, _29231_);
  and (_39050_, _39036_, _24456_);
  and (_39051_, _39050_, _28676_);
  nor (_39052_, _39050_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not (_39053_, _39052_);
  and (_39054_, _39053_, _39041_);
  not (_39055_, _39054_);
  nor (_39056_, _39055_, _39051_);
  or (_39057_, _39056_, _39049_);
  and (_39058_, _39057_, _39022_);
  nor (_39059_, _39022_, _38617_);
  or (_39060_, _39059_, _39058_);
  and (_24174_, _39060_, _41806_);
  and (_39061_, _39021_, _38645_);
  nor (_39062_, _39032_, _29893_);
  and (_39063_, _39036_, _30002_);
  and (_39064_, _39063_, _28676_);
  nor (_39065_, _39063_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not (_39066_, _39065_);
  and (_39067_, _39066_, _39041_);
  not (_39068_, _39067_);
  nor (_39069_, _39068_, _39064_);
  nor (_39070_, _39069_, _39021_);
  not (_39071_, _39070_);
  nor (_39072_, _39071_, _39062_);
  nor (_39073_, _39072_, _39061_);
  and (_24186_, _39073_, _41806_);
  nor (_39074_, _39032_, _30567_);
  nor (_39075_, _25113_, _24949_);
  and (_39076_, _39075_, _25244_);
  and (_39077_, _28742_, _24807_);
  and (_39078_, _39077_, _39076_);
  not (_39079_, _39078_);
  and (_39080_, _39041_, _39079_);
  and (_39081_, _39080_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_39082_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_39083_, _30708_, _39082_);
  nor (_39084_, _39083_, _30719_);
  and (_39085_, _39041_, _39078_);
  not (_39086_, _39085_);
  nor (_39087_, _39086_, _39084_);
  nor (_39088_, _39087_, _39081_);
  and (_39089_, _39088_, _39022_);
  not (_39090_, _39089_);
  nor (_39091_, _39090_, _39074_);
  and (_39092_, _39021_, _38673_);
  or (_39093_, _39092_, _39091_);
  nor (_24198_, _39093_, rst);
  nor (_39094_, _39032_, _31338_);
  and (_39095_, _39080_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_39096_, _31447_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39097_, _39096_, _31458_);
  nor (_39098_, _39097_, _39086_);
  nor (_39099_, _39098_, _39095_);
  not (_39100_, _39099_);
  nor (_39101_, _39100_, _39094_);
  nor (_39102_, _39101_, _39021_);
  nor (_39103_, _39022_, _38702_);
  nor (_39104_, _39103_, _39102_);
  nor (_24210_, _39104_, rst);
  nor (_39105_, _39032_, _32044_);
  and (_39106_, _39036_, _32131_);
  and (_39107_, _39106_, _28676_);
  nor (_39108_, _39106_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_39109_, _39108_);
  and (_39110_, _39109_, _39041_);
  not (_39111_, _39110_);
  nor (_39112_, _39111_, _39107_);
  or (_39113_, _39112_, _39105_);
  and (_39114_, _39113_, _39022_);
  nor (_39115_, _39022_, _38731_);
  or (_39116_, _39115_, _39114_);
  and (_24222_, _39116_, _41806_);
  nor (_39117_, _39032_, _32853_);
  and (_39118_, _39036_, _32941_);
  and (_39119_, _39118_, _28676_);
  nor (_39120_, _39118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_39121_, _39120_);
  and (_39122_, _39121_, _39041_);
  not (_39123_, _39122_);
  nor (_39124_, _39123_, _39119_);
  or (_39125_, _39124_, _39117_);
  and (_39126_, _39125_, _39022_);
  nor (_39127_, _39022_, _38760_);
  or (_39128_, _39127_, _39126_);
  and (_24234_, _39128_, _41806_);
  nor (_39129_, _39032_, _33598_);
  and (_39130_, _39036_, _33697_);
  and (_39131_, _39130_, _28676_);
  nor (_39132_, _39130_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not (_39133_, _39132_);
  and (_39134_, _39133_, _39041_);
  not (_39135_, _39134_);
  nor (_39136_, _39135_, _39131_);
  or (_39137_, _39136_, _39129_);
  and (_39138_, _39137_, _39022_);
  nor (_39139_, _39022_, _38787_);
  or (_39140_, _39139_, _39138_);
  and (_24246_, _39140_, _41806_);
  and (_39141_, _38019_, _28709_);
  nand (_39142_, _39141_, _28676_);
  or (_39143_, _39141_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39144_, _39143_, _28742_);
  and (_39145_, _39144_, _39142_);
  and (_39146_, _38008_, _39026_);
  nand (_39147_, _39146_, _38162_);
  or (_39148_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39149_, _39148_, _28087_);
  and (_39150_, _39149_, _39147_);
  not (_39151_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_39152_, _28076_, _39151_);
  or (_39153_, _39152_, rst);
  or (_39154_, _39153_, _39150_);
  or (_35484_, _39154_, _39145_);
  nor (_39155_, _38950_, _24949_);
  and (_39156_, _38819_, _39155_);
  and (_39157_, _39156_, _28709_);
  nand (_39158_, _39157_, _28676_);
  or (_39159_, _39157_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39160_, _39159_, _28742_);
  and (_39161_, _39160_, _39158_);
  and (_39162_, _39156_, _24456_);
  not (_39163_, _39162_);
  nor (_39164_, _39163_, _38162_);
  not (_39165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_39166_, _39162_, _39165_);
  or (_39167_, _39166_, _39164_);
  and (_39168_, _39167_, _28087_);
  nor (_39169_, _28076_, _39165_);
  or (_39170_, _39169_, rst);
  or (_39171_, _39170_, _39168_);
  or (_35507_, _39171_, _39161_);
  and (_39172_, _39027_, _24665_);
  and (_39173_, _39172_, _39076_);
  and (_39174_, _39173_, _28709_);
  nand (_39175_, _39174_, _28676_);
  or (_39176_, _39174_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39177_, _39176_, _28742_);
  and (_39178_, _39177_, _39175_);
  and (_39179_, _39028_, _39155_);
  and (_39180_, _39179_, _39026_);
  not (_39181_, _39180_);
  nor (_39182_, _39181_, _38162_);
  not (_39183_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_39184_, _39180_, _39183_);
  or (_39185_, _39184_, _39182_);
  and (_39186_, _39185_, _28087_);
  nor (_39187_, _28076_, _39183_);
  or (_39188_, _39187_, rst);
  or (_39189_, _39188_, _39186_);
  or (_35530_, _39189_, _39178_);
  and (_39190_, _39172_, _25266_);
  and (_39191_, _39190_, _28709_);
  nand (_39192_, _39191_, _28676_);
  or (_39193_, _39191_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_39194_, _39193_, _28742_);
  and (_39195_, _39194_, _39192_);
  nor (_39196_, _25244_, _24796_);
  and (_39203_, _39155_, _39196_);
  and (_39214_, _39203_, _39026_);
  not (_39225_, _39214_);
  nor (_39235_, _39225_, _38162_);
  not (_39241_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_39251_, _39214_, _39241_);
  or (_39262_, _39251_, _39235_);
  and (_39273_, _39262_, _28087_);
  nor (_39284_, _28076_, _39241_);
  or (_39295_, _39284_, rst);
  or (_39306_, _39295_, _39273_);
  or (_35552_, _39306_, _39195_);
  not (_39327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39338_, _39146_, _39327_);
  nand (_39349_, _38019_, _24456_);
  nor (_39360_, _39349_, _28676_);
  or (_39371_, _39360_, _39338_);
  and (_39382_, _39371_, _28742_);
  and (_39393_, _39146_, _38426_);
  or (_39404_, _39393_, _39338_);
  and (_39410_, _39404_, _28087_);
  nor (_39411_, _28076_, _39327_);
  or (_39412_, _39411_, rst);
  or (_39413_, _39412_, _39410_);
  or (_41207_, _39413_, _39382_);
  or (_39414_, _38030_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39415_, _39414_, _28742_);
  nand (_39416_, _38205_, _28676_);
  and (_39417_, _39416_, _39415_);
  nand (_39418_, _39146_, _38417_);
  or (_39419_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39420_, _39419_, _28087_);
  and (_39421_, _39420_, _39418_);
  not (_39422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_39423_, _28076_, _39422_);
  or (_39424_, _39423_, rst);
  or (_39425_, _39424_, _39421_);
  or (_41209_, _39425_, _39417_);
  not (_39426_, _31468_);
  nand (_39427_, _38019_, _39426_);
  and (_39428_, _39427_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39429_, _30730_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39430_, _39429_, _30719_);
  and (_39431_, _39430_, _38019_);
  or (_39432_, _39431_, _39428_);
  and (_39433_, _39432_, _28742_);
  nand (_39434_, _39146_, _38410_);
  or (_39435_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39436_, _39435_, _28087_);
  and (_39437_, _39436_, _39434_);
  not (_39438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_39439_, _28076_, _39438_);
  or (_39440_, _39439_, rst);
  or (_39441_, _39440_, _39437_);
  or (_41211_, _39441_, _39433_);
  not (_39442_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_39443_, _38194_, _39442_);
  nor (_39444_, _31468_, _39442_);
  or (_39445_, _39444_, _31458_);
  and (_39446_, _39445_, _38019_);
  or (_39447_, _39446_, _39443_);
  and (_39448_, _39447_, _28742_);
  nand (_39449_, _39146_, _38402_);
  or (_39450_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39451_, _39450_, _28087_);
  and (_39452_, _39451_, _39449_);
  nor (_39453_, _28076_, _39442_);
  or (_39454_, _39453_, rst);
  or (_39455_, _39454_, _39452_);
  or (_41213_, _39455_, _39448_);
  nand (_39456_, _38019_, _32163_);
  and (_39457_, _39456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39458_, _32142_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39459_, _39458_, _32196_);
  and (_39460_, _39459_, _38019_);
  or (_39461_, _39460_, _39457_);
  and (_39462_, _39461_, _28742_);
  nand (_39463_, _39146_, _38394_);
  or (_39464_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39465_, _39464_, _28087_);
  and (_39466_, _39465_, _39463_);
  not (_39467_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_39468_, _28076_, _39467_);
  or (_39469_, _39468_, rst);
  or (_39470_, _39469_, _39466_);
  or (_41214_, _39470_, _39462_);
  and (_39471_, _38019_, _32941_);
  nand (_39472_, _39471_, _28676_);
  or (_39473_, _39471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39474_, _39473_, _28742_);
  and (_39475_, _39474_, _39472_);
  nand (_39476_, _39146_, _38366_);
  or (_39477_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39478_, _39477_, _28087_);
  and (_39479_, _39478_, _39476_);
  not (_39480_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_39481_, _28076_, _39480_);
  or (_39482_, _39481_, rst);
  or (_39483_, _39482_, _39479_);
  or (_41216_, _39483_, _39475_);
  and (_39484_, _38019_, _33697_);
  nand (_39485_, _39484_, _28676_);
  or (_39486_, _39484_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39487_, _39486_, _28742_);
  and (_39488_, _39487_, _39485_);
  nand (_39489_, _39146_, _38280_);
  or (_39490_, _39146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39491_, _39490_, _28087_);
  and (_39492_, _39491_, _39489_);
  not (_39493_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_39494_, _28076_, _39493_);
  or (_39495_, _39494_, rst);
  or (_39496_, _39495_, _39492_);
  or (_41218_, _39496_, _39488_);
  nand (_39497_, _39162_, _28676_);
  or (_39498_, _39162_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39499_, _39498_, _28742_);
  and (_39500_, _39499_, _39497_);
  nor (_39501_, _39163_, _38425_);
  not (_39502_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_39503_, _39162_, _39502_);
  or (_39504_, _39503_, _39501_);
  and (_39505_, _39504_, _28087_);
  nor (_39506_, _28076_, _39502_);
  or (_39507_, _39506_, rst);
  or (_39508_, _39507_, _39505_);
  or (_41220_, _39508_, _39500_);
  and (_39509_, _39156_, _30002_);
  nand (_39510_, _39509_, _28676_);
  or (_39511_, _39509_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39512_, _39511_, _28742_);
  and (_39513_, _39512_, _39510_);
  nor (_39514_, _39163_, _38417_);
  not (_39515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_39516_, _39162_, _39515_);
  or (_39517_, _39516_, _39514_);
  and (_39518_, _39517_, _28087_);
  nor (_39519_, _28076_, _39515_);
  or (_39520_, _39519_, rst);
  or (_39521_, _39520_, _39518_);
  or (_41221_, _39521_, _39513_);
  and (_39522_, _39156_, _30708_);
  nand (_39523_, _39522_, _28676_);
  or (_39524_, _39522_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39525_, _39524_, _28742_);
  and (_39526_, _39525_, _39523_);
  nor (_39527_, _39163_, _38410_);
  not (_39528_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_39529_, _39162_, _39528_);
  or (_39530_, _39529_, _39527_);
  and (_39531_, _39530_, _28087_);
  nor (_39532_, _28076_, _39528_);
  or (_39533_, _39532_, rst);
  or (_39534_, _39533_, _39531_);
  or (_41223_, _39534_, _39526_);
  and (_39535_, _39156_, _31436_);
  nand (_39536_, _39535_, _28676_);
  or (_39537_, _39535_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39538_, _39537_, _28742_);
  and (_39539_, _39538_, _39536_);
  nor (_39540_, _39163_, _38402_);
  not (_39541_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_39542_, _39162_, _39541_);
  or (_39543_, _39542_, _39540_);
  and (_39544_, _39543_, _28087_);
  nor (_39545_, _28076_, _39541_);
  or (_39546_, _39545_, rst);
  or (_39547_, _39546_, _39544_);
  or (_41225_, _39547_, _39539_);
  and (_39548_, _39156_, _32131_);
  nand (_39549_, _39548_, _28676_);
  or (_39550_, _39548_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39551_, _39550_, _28742_);
  and (_39552_, _39551_, _39549_);
  nor (_39553_, _39163_, _38394_);
  not (_39554_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_39555_, _39162_, _39554_);
  or (_39556_, _39555_, _39553_);
  and (_39557_, _39556_, _28087_);
  nor (_39558_, _28076_, _39554_);
  or (_39559_, _39558_, rst);
  or (_39560_, _39559_, _39557_);
  or (_41227_, _39560_, _39552_);
  and (_39561_, _39156_, _32941_);
  nand (_39562_, _39561_, _28676_);
  or (_39563_, _39561_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39564_, _39563_, _28742_);
  and (_39565_, _39564_, _39562_);
  nor (_39566_, _39163_, _38366_);
  not (_39567_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_39568_, _39162_, _39567_);
  or (_39569_, _39568_, _39566_);
  and (_39570_, _39569_, _28087_);
  nor (_39571_, _28076_, _39567_);
  or (_39572_, _39571_, rst);
  or (_39573_, _39572_, _39570_);
  or (_41228_, _39573_, _39565_);
  and (_39574_, _39156_, _33697_);
  nand (_39575_, _39574_, _28676_);
  or (_39576_, _39574_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39577_, _39576_, _28742_);
  and (_39578_, _39577_, _39575_);
  nor (_39579_, _39163_, _38280_);
  not (_39580_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_39581_, _39162_, _39580_);
  or (_39582_, _39581_, _39579_);
  and (_39583_, _39582_, _28087_);
  nor (_39584_, _28076_, _39580_);
  or (_39585_, _39584_, rst);
  or (_39586_, _39585_, _39583_);
  or (_41230_, _39586_, _39578_);
  nand (_39587_, _39180_, _28676_);
  or (_39588_, _39180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39589_, _39588_, _28742_);
  and (_39590_, _39589_, _39587_);
  nor (_39591_, _39181_, _38425_);
  not (_39592_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_39593_, _39180_, _39592_);
  or (_39594_, _39593_, _39591_);
  and (_39595_, _39594_, _28087_);
  nor (_39596_, _28076_, _39592_);
  or (_39597_, _39596_, rst);
  or (_39598_, _39597_, _39595_);
  or (_41232_, _39598_, _39590_);
  and (_39599_, _39173_, _30002_);
  nand (_39600_, _39599_, _28676_);
  or (_39601_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39602_, _39601_, _28742_);
  and (_39603_, _39602_, _39600_);
  nor (_39604_, _39181_, _38417_);
  not (_39605_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_39606_, _39180_, _39605_);
  or (_39607_, _39606_, _39604_);
  and (_39608_, _39607_, _28087_);
  nor (_39609_, _28076_, _39605_);
  or (_39610_, _39609_, rst);
  or (_39611_, _39610_, _39608_);
  or (_41234_, _39611_, _39603_);
  and (_39612_, _39173_, _30708_);
  nand (_39613_, _39612_, _28676_);
  or (_39614_, _39612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39615_, _39614_, _28742_);
  and (_39616_, _39615_, _39613_);
  nor (_39618_, _39181_, _38410_);
  not (_39619_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_39620_, _39180_, _39619_);
  or (_39621_, _39620_, _39618_);
  and (_39622_, _39621_, _28087_);
  nor (_39623_, _28076_, _39619_);
  or (_39624_, _39623_, rst);
  or (_39625_, _39624_, _39622_);
  or (_41235_, _39625_, _39616_);
  and (_39626_, _39173_, _31436_);
  nand (_39627_, _39626_, _28676_);
  or (_39628_, _39626_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39629_, _39628_, _28742_);
  and (_39630_, _39629_, _39627_);
  nor (_39631_, _39181_, _38402_);
  not (_39632_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_39633_, _39180_, _39632_);
  or (_39634_, _39633_, _39631_);
  and (_39635_, _39634_, _28087_);
  nor (_39636_, _28076_, _39632_);
  or (_39637_, _39636_, rst);
  or (_39638_, _39637_, _39635_);
  or (_41237_, _39638_, _39630_);
  and (_39639_, _39173_, _32131_);
  nand (_39640_, _39639_, _28676_);
  or (_39641_, _39639_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39642_, _39641_, _28742_);
  and (_39643_, _39642_, _39640_);
  nor (_39644_, _39181_, _38394_);
  not (_39645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_39646_, _39180_, _39645_);
  or (_39647_, _39646_, _39644_);
  and (_39652_, _39647_, _28087_);
  nor (_39653_, _28076_, _39645_);
  or (_39654_, _39653_, rst);
  or (_39655_, _39654_, _39652_);
  or (_41239_, _39655_, _39643_);
  and (_39656_, _39173_, _32941_);
  nand (_39657_, _39656_, _28676_);
  or (_39658_, _39656_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39659_, _39658_, _28742_);
  and (_39660_, _39659_, _39657_);
  nor (_39661_, _39181_, _38366_);
  not (_39662_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_39663_, _39180_, _39662_);
  or (_39664_, _39663_, _39661_);
  and (_39665_, _39664_, _28087_);
  nor (_39666_, _28076_, _39662_);
  or (_39667_, _39666_, rst);
  or (_39668_, _39667_, _39665_);
  or (_41240_, _39668_, _39660_);
  and (_39669_, _39173_, _33697_);
  nand (_39670_, _39669_, _28676_);
  or (_39671_, _39669_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39672_, _39671_, _28742_);
  and (_39673_, _39672_, _39670_);
  nor (_39674_, _39181_, _38280_);
  not (_39675_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_39676_, _39180_, _39675_);
  or (_39677_, _39676_, _39674_);
  and (_39678_, _39677_, _28087_);
  nor (_39679_, _28076_, _39675_);
  or (_39680_, _39679_, rst);
  or (_39681_, _39680_, _39678_);
  or (_41242_, _39681_, _39673_);
  and (_39682_, _39190_, _24456_);
  nand (_39683_, _39682_, _28676_);
  or (_39684_, _39682_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39685_, _39684_, _28742_);
  and (_39686_, _39685_, _39683_);
  nor (_39687_, _39225_, _38425_);
  not (_39688_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_39689_, _39214_, _39688_);
  or (_39690_, _39689_, _39687_);
  and (_39691_, _39690_, _28087_);
  nor (_39692_, _28076_, _39688_);
  or (_39693_, _39692_, rst);
  or (_39694_, _39693_, _39691_);
  or (_41244_, _39694_, _39686_);
  and (_39695_, _39190_, _30002_);
  nand (_39696_, _39695_, _28676_);
  or (_39697_, _39695_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39698_, _39697_, _28742_);
  and (_39699_, _39698_, _39696_);
  nor (_39700_, _39225_, _38417_);
  not (_39701_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_39702_, _39214_, _39701_);
  or (_39703_, _39702_, _39700_);
  and (_39704_, _39703_, _28087_);
  nor (_39705_, _28076_, _39701_);
  or (_39706_, _39705_, rst);
  or (_39707_, _39706_, _39704_);
  or (_41245_, _39707_, _39699_);
  and (_39708_, _39190_, _30708_);
  nand (_39709_, _39708_, _28676_);
  or (_39710_, _39708_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39711_, _39710_, _28742_);
  and (_39712_, _39711_, _39709_);
  nor (_39720_, _39225_, _38410_);
  not (_39721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_39722_, _39214_, _39721_);
  or (_39723_, _39722_, _39720_);
  and (_39724_, _39723_, _28087_);
  nor (_39725_, _28076_, _39721_);
  or (_39726_, _39725_, rst);
  or (_39727_, _39726_, _39724_);
  or (_41247_, _39727_, _39712_);
  and (_39728_, _39190_, _31436_);
  nand (_39729_, _39728_, _28676_);
  or (_39730_, _39728_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39731_, _39730_, _28742_);
  and (_39732_, _39731_, _39729_);
  nor (_39733_, _39225_, _38402_);
  not (_39734_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_39735_, _39214_, _39734_);
  or (_39736_, _39735_, _39733_);
  and (_39737_, _39736_, _28087_);
  nor (_39738_, _28076_, _39734_);
  or (_39739_, _39738_, rst);
  or (_39740_, _39739_, _39737_);
  or (_41249_, _39740_, _39732_);
  and (_39741_, _39190_, _32131_);
  nand (_39742_, _39741_, _28676_);
  or (_39743_, _39741_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39744_, _39743_, _28742_);
  and (_39745_, _39744_, _39742_);
  nor (_39746_, _39225_, _38394_);
  not (_39747_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_39748_, _39214_, _39747_);
  or (_39749_, _39748_, _39746_);
  and (_39750_, _39749_, _28087_);
  nor (_39751_, _28076_, _39747_);
  or (_39752_, _39751_, rst);
  or (_39753_, _39752_, _39750_);
  or (_41251_, _39753_, _39745_);
  and (_39754_, _39190_, _32941_);
  nand (_39755_, _39754_, _28676_);
  or (_39756_, _39754_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39757_, _39756_, _28742_);
  and (_39758_, _39757_, _39755_);
  nor (_39759_, _39225_, _38366_);
  not (_39760_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_39761_, _39214_, _39760_);
  or (_39762_, _39761_, _39759_);
  and (_39763_, _39762_, _28087_);
  nor (_39768_, _28076_, _39760_);
  or (_39769_, _39768_, rst);
  or (_39770_, _39769_, _39763_);
  or (_41252_, _39770_, _39758_);
  and (_39771_, _39190_, _33697_);
  nand (_39772_, _39771_, _28676_);
  or (_39773_, _39771_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39774_, _39773_, _28742_);
  and (_39775_, _39774_, _39772_);
  nor (_39776_, _39225_, _38280_);
  not (_39777_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_39778_, _39214_, _39777_);
  or (_39779_, _39778_, _39776_);
  and (_39780_, _39779_, _28087_);
  nor (_39781_, _28076_, _39777_);
  or (_39782_, _39781_, rst);
  or (_39792_, _39782_, _39780_);
  or (_41254_, _39792_, _39775_);
  and (_39793_, _38817_, _25113_);
  and (_39794_, _39793_, _39203_);
  nor (_39795_, _25244_, _25112_);
  and (_39796_, _39795_, _39172_);
  and (_39797_, _39796_, _38953_);
  and (_39798_, _39797_, _28709_);
  nand (_39799_, _39798_, _28676_);
  or (_39800_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_39801_, _39800_, _39799_);
  or (_39802_, _39801_, _39794_);
  nand (_39803_, _39794_, _38162_);
  and (_39804_, _39803_, _41806_);
  and (_41748_, _39804_, _39802_);
  and (_39805_, _39793_, _39179_);
  and (_39806_, _25244_, _25113_);
  and (_39807_, _39806_, _38953_);
  and (_39808_, _39807_, _39172_);
  and (_39809_, _39808_, _28709_);
  nand (_39810_, _39809_, _28676_);
  or (_39811_, _39809_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_39812_, _39811_, _39810_);
  or (_39813_, _39812_, _39805_);
  nand (_39814_, _39805_, _38162_);
  and (_39815_, _39814_, _41806_);
  and (_41751_, _39815_, _39813_);
  or (_39816_, _24445_, _30697_);
  and (_39817_, _39816_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39818_, _39817_, _38972_);
  and (_39819_, _39807_, _37986_);
  and (_39820_, _39819_, _39818_);
  and (_39821_, _39793_, _38008_);
  nand (_39822_, _39819_, _24434_);
  and (_39823_, _39822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39824_, _39823_, _39821_);
  or (_39825_, _39824_, _39820_);
  nand (_39826_, _39821_, _38280_);
  and (_39827_, _39826_, _41806_);
  and (_41753_, _39827_, _39825_);
  not (_39828_, _39821_);
  not (_39829_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_39830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_39831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_39832_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _39831_);
  and (_39833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39834_, _39833_, _39832_);
  nor (_39835_, _39834_, _39830_);
  or (_39836_, _39835_, _39829_);
  and (_39837_, _39831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_39838_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_39839_, _39838_, _39837_);
  nor (_39840_, _39839_, _39830_);
  and (_39841_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _39831_);
  and (_39842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39843_, _39842_, _39841_);
  nand (_39844_, _39843_, _39840_);
  or (_39845_, _39844_, _39836_);
  and (_39846_, _39845_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor (_39847_, _24197_, _25112_);
  and (_39848_, _28742_, _28698_);
  and (_39849_, _39848_, _38008_);
  and (_39850_, _39849_, _39847_);
  or (_39851_, _39850_, _39846_);
  and (_39852_, _39851_, _39828_);
  nand (_39853_, _39850_, _28676_);
  and (_39854_, _39853_, _39852_);
  nor (_39855_, _39828_, _38162_);
  or (_39856_, _39855_, _39854_);
  and (_41755_, _39856_, _41806_);
  nor (_39857_, _39843_, _39830_);
  nand (_39858_, _39857_, _39839_);
  or (_39859_, _39858_, _39836_);
  and (_39860_, _39859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_39861_, _28742_, _29991_);
  and (_39862_, _39861_, _38008_);
  and (_39863_, _39862_, _39847_);
  or (_39864_, _39863_, _39860_);
  and (_39865_, _39864_, _39828_);
  nand (_39866_, _39863_, _28676_);
  and (_39867_, _39866_, _39865_);
  nor (_39868_, _39828_, _38366_);
  or (_39869_, _39868_, _39867_);
  and (_41757_, _39869_, _41806_);
  not (_39870_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_39871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _39870_);
  nand (_39872_, _39835_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_39873_, _39857_, _39840_);
  or (_39874_, _39873_, _39872_);
  and (_39875_, _39874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_39876_, _39875_, _39871_);
  nor (_39877_, _28687_, _25112_);
  and (_39878_, _39862_, _39877_);
  or (_39879_, _39878_, _39876_);
  and (_39880_, _39879_, _39828_);
  nand (_39881_, _39878_, _28676_);
  and (_39882_, _39881_, _39880_);
  nor (_39883_, _39828_, _38417_);
  or (_39884_, _39883_, _39882_);
  and (_41759_, _39884_, _41806_);
  and (_39885_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_39886_, _39872_, _39858_);
  and (_39887_, _39886_, _39885_);
  and (_39888_, _39849_, _39877_);
  or (_39889_, _39888_, _39887_);
  and (_39890_, _39889_, _39828_);
  nand (_39891_, _39888_, _28676_);
  and (_39892_, _39891_, _39890_);
  nor (_39893_, _39828_, _38402_);
  or (_39894_, _39893_, _39892_);
  and (_41761_, _39894_, _41806_);
  and (_39895_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_39896_, _39895_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_39897_, _39896_);
  and (_39898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_39899_, _39898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_39900_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_39901_, _39900_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_39902_, _39901_, _39899_);
  and (_39903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_39904_, _39903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  not (_39905_, _39904_);
  and (_39906_, _39905_, _39902_);
  and (_39907_, _39906_, _39897_);
  not (_39908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_39909_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_39910_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _39831_);
  or (_39911_, _39910_, _39909_);
  nor (_39912_, _39911_, _39908_);
  nor (_39913_, _39912_, _39830_);
  nor (_39914_, _39913_, _39907_);
  and (_39915_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_39916_, _39915_, _39831_);
  and (_39917_, _39916_, _39914_);
  and (_39918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _39830_);
  not (_39919_, _39918_);
  not (_39920_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_39921_, _39898_, _39920_);
  not (_39922_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_39923_, _39900_, _39922_);
  nor (_39924_, _39923_, _39921_);
  not (_39925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_39926_, _39903_, _39925_);
  not (_39927_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_39928_, _39895_, _39927_);
  nor (_39929_, _39928_, _39926_);
  and (_39930_, _39929_, _39924_);
  nor (_39931_, _39930_, _39919_);
  nand (_39932_, _39931_, _39916_);
  and (_39933_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41806_);
  nand (_39934_, _39933_, _39932_);
  nor (_41793_, _39934_, _39917_);
  nor (_39935_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_39936_, _39935_);
  nor (_39937_, _39931_, _39914_);
  nor (_39938_, _39937_, _39936_);
  nand (_39939_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41806_);
  nor (_41795_, _39939_, _39938_);
  and (_39940_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_39941_, _39902_);
  or (_39942_, _39941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_39943_, _39942_, _39940_);
  or (_39944_, _39906_, _39837_);
  and (_39945_, _39944_, _39943_);
  and (_39946_, _39945_, _39914_);
  or (_39947_, _39946_, _39915_);
  and (_39948_, _39937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_39949_, _39914_);
  and (_39950_, _39931_, _39949_);
  and (_39951_, _39928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_39952_, _39951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_39953_, _39924_);
  and (_39954_, _39926_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39955_, _39954_, _39953_);
  and (_39956_, _39955_, _39952_);
  and (_39957_, _39953_, _39837_);
  or (_39958_, _39957_, _39956_);
  and (_39959_, _39958_, _39950_);
  or (_39960_, _39959_, _39948_);
  or (_39961_, _39960_, _39947_);
  not (_39962_, _39915_);
  or (_39963_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_39964_, _39963_, _41806_);
  and (_41796_, _39964_, _39961_);
  and (_39965_, _39896_, _39831_);
  or (_39966_, _39941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_39967_, _39966_, _39965_);
  or (_39968_, _39906_, _39838_);
  and (_39969_, _39968_, _39967_);
  and (_39970_, _39969_, _39914_);
  or (_39971_, _39970_, _39915_);
  and (_39972_, _39937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_39973_, _39928_, _39831_);
  or (_39974_, _39973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_39975_, _39926_, _39831_);
  nor (_39976_, _39975_, _39953_);
  and (_39977_, _39976_, _39974_);
  and (_39978_, _39953_, _39838_);
  or (_39979_, _39978_, _39977_);
  and (_39980_, _39979_, _39950_);
  or (_39981_, _39980_, _39972_);
  or (_39982_, _39981_, _39971_);
  or (_39983_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_39984_, _39983_, _41806_);
  and (_41798_, _39984_, _39982_);
  nand (_39985_, _39937_, _39830_);
  nor (_39986_, _39831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_39987_, _39986_, _39915_);
  and (_39988_, _39987_, _41806_);
  and (_41800_, _39988_, _39985_);
  and (_39989_, _39937_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_39990_, _39831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_39991_, _39990_, _39986_);
  nor (_39992_, _39991_, _39949_);
  or (_39993_, _39992_, _39915_);
  or (_39994_, _39993_, _39989_);
  or (_39995_, _39991_, _39962_);
  and (_39996_, _39995_, _41806_);
  and (_41802_, _39996_, _39994_);
  and (_39997_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41806_);
  and (_41804_, _39997_, _39915_);
  nor (_39998_, _39937_, _39915_);
  and (_39999_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_40000_, _39999_, _39998_);
  and (_42729_, _40000_, _41806_);
  and (_40001_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_40002_, _40001_, _39998_);
  and (_42731_, _40002_, _41806_);
  and (_40003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _41806_);
  and (_42733_, _40003_, _39915_);
  not (_40004_, _39921_);
  nor (_40005_, _39928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_40006_, _40005_, _39926_);
  or (_40007_, _40006_, _39923_);
  and (_40008_, _40007_, _40004_);
  and (_40009_, _40008_, _39950_);
  not (_40010_, _39899_);
  or (_40011_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40012_, _40011_, _39905_);
  or (_40013_, _40012_, _39901_);
  and (_40014_, _40013_, _40010_);
  and (_40015_, _40014_, _39914_);
  or (_40016_, _40015_, _39915_);
  or (_40017_, _40016_, _40009_);
  or (_40018_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40019_, _40018_, _41806_);
  and (_42734_, _40019_, _40017_);
  nand (_40020_, _39924_, _39918_);
  nor (_40021_, _40020_, _39929_);
  or (_40022_, _40021_, _39914_);
  nand (_40023_, _39914_, _39941_);
  and (_40024_, _40023_, _40022_);
  or (_40025_, _40024_, _39915_);
  or (_40026_, _39962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_40027_, _40026_, _41806_);
  and (_42736_, _40027_, _40025_);
  and (_40028_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _41806_);
  and (_42738_, _40028_, _39915_);
  and (_40029_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _41806_);
  and (_42740_, _40029_, _39915_);
  nand (_40030_, _39937_, _39935_);
  nor (_40031_, _39915_, _39914_);
  or (_40032_, _40031_, _39831_);
  and (_40033_, _40032_, _41806_);
  and (_42742_, _40033_, _40030_);
  not (_40034_, _39998_);
  and (_40035_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_40036_, _39965_);
  and (_40037_, _40036_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_40038_, _39904_, _39831_);
  or (_40039_, _40038_, _39901_);
  or (_40040_, _40039_, _40037_);
  not (_40041_, _39901_);
  or (_40042_, _40041_, _39833_);
  and (_40043_, _40042_, _40040_);
  or (_40044_, _40043_, _39899_);
  or (_40045_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _39831_);
  or (_40046_, _40045_, _40010_);
  and (_40047_, _40046_, _39914_);
  and (_40048_, _40047_, _40044_);
  not (_40049_, _39973_);
  and (_40050_, _40049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_40051_, _39975_, _39923_);
  or (_40052_, _40051_, _40050_);
  not (_40053_, _39923_);
  or (_40054_, _40053_, _39833_);
  and (_40055_, _40054_, _40004_);
  and (_40056_, _40055_, _40052_);
  and (_40057_, _40045_, _39921_);
  or (_40058_, _40057_, _40056_);
  and (_40059_, _40058_, _39950_);
  or (_40060_, _40059_, _40048_);
  and (_40061_, _40060_, _39962_);
  or (_40062_, _40061_, _40035_);
  and (_42744_, _40062_, _41806_);
  and (_40063_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40064_, _40036_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40065_, _40064_, _40039_);
  or (_40066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _39831_);
  or (_40067_, _40066_, _40041_);
  and (_40068_, _40067_, _40010_);
  and (_40069_, _40068_, _40065_);
  and (_40070_, _39899_, _39842_);
  or (_40071_, _40070_, _40069_);
  and (_40072_, _40071_, _39914_);
  and (_40073_, _40049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40074_, _40073_, _40051_);
  or (_40075_, _40066_, _40053_);
  and (_40076_, _40075_, _40004_);
  and (_40077_, _40076_, _40074_);
  and (_40078_, _39921_, _39842_);
  or (_40079_, _40078_, _40077_);
  and (_40080_, _40079_, _39950_);
  or (_40081_, _40080_, _40072_);
  and (_40082_, _40081_, _39962_);
  or (_40083_, _40082_, _40063_);
  and (_42746_, _40083_, _41806_);
  and (_40084_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_40085_, _39940_);
  and (_40086_, _40085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_40087_, _39904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40088_, _40087_, _39901_);
  or (_40089_, _40088_, _40086_);
  or (_40090_, _40041_, _39832_);
  and (_40091_, _40090_, _40089_);
  or (_40092_, _40091_, _39899_);
  or (_40093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40094_, _40093_, _40010_);
  and (_40095_, _40094_, _39914_);
  and (_40096_, _40095_, _40092_);
  not (_40097_, _39951_);
  and (_40098_, _40097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_40099_, _39954_, _39923_);
  or (_40100_, _40099_, _40098_);
  or (_40101_, _40053_, _39832_);
  and (_40102_, _40101_, _40004_);
  and (_40103_, _40102_, _40100_);
  and (_40104_, _40093_, _39921_);
  or (_40105_, _40104_, _40103_);
  and (_40106_, _40105_, _39950_);
  or (_40107_, _40106_, _40096_);
  and (_40108_, _40107_, _39962_);
  or (_40109_, _40108_, _40084_);
  and (_42748_, _40109_, _41806_);
  and (_40110_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40111_, _40085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40112_, _40111_, _40088_);
  or (_40113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40114_, _40113_, _40041_);
  and (_40115_, _40114_, _40010_);
  and (_40116_, _40115_, _40112_);
  and (_40117_, _39899_, _39841_);
  or (_40118_, _40117_, _40116_);
  and (_40119_, _40118_, _39914_);
  and (_40120_, _40097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40121_, _40120_, _40099_);
  or (_40122_, _40113_, _40053_);
  and (_40123_, _40122_, _40004_);
  and (_40124_, _40123_, _40121_);
  and (_40125_, _39921_, _39841_);
  or (_40126_, _40125_, _40124_);
  and (_40127_, _40126_, _39950_);
  or (_40128_, _40127_, _40119_);
  and (_40129_, _40128_, _39962_);
  or (_40130_, _40129_, _40110_);
  and (_42750_, _40130_, _41806_);
  and (_40131_, _39935_, _39914_);
  nand (_40132_, _39935_, _39931_);
  and (_40133_, _40132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_40134_, _40133_, _40131_);
  and (_42752_, _40134_, _41806_);
  and (_40135_, _39932_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_40136_, _40135_, _39917_);
  and (_42754_, _40136_, _41806_);
  and (_40137_, _39819_, _24456_);
  or (_40138_, _40137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_40139_, _40138_, _39828_);
  nand (_40140_, _40137_, _28676_);
  and (_40141_, _40140_, _40139_);
  nor (_40142_, _39828_, _38425_);
  or (_40143_, _40142_, _40141_);
  and (_42756_, _40143_, _41806_);
  and (_40144_, _39819_, _30708_);
  nand (_40145_, _40144_, _28676_);
  or (_40146_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_40147_, _40146_, _39828_);
  and (_40148_, _40147_, _40145_);
  nor (_40149_, _39828_, _38410_);
  or (_40150_, _40149_, _40148_);
  and (_42758_, _40150_, _41806_);
  and (_40151_, _39819_, _32131_);
  nand (_40152_, _40151_, _28676_);
  or (_40153_, _40151_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_40154_, _40153_, _39828_);
  and (_40155_, _40154_, _40152_);
  nor (_40156_, _39828_, _38394_);
  or (_40157_, _40156_, _40155_);
  and (_42760_, _40157_, _41806_);
  and (_40158_, _39808_, _24456_);
  nand (_40159_, _40158_, _28676_);
  not (_40160_, _39805_);
  or (_40161_, _40158_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40162_, _40161_, _40160_);
  and (_40163_, _40162_, _40159_);
  nor (_40164_, _40160_, _38425_);
  or (_40165_, _40164_, _40163_);
  and (_42762_, _40165_, _41806_);
  and (_40166_, _39808_, _30002_);
  nand (_40167_, _40166_, _28676_);
  or (_40168_, _40166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40169_, _40168_, _40160_);
  and (_40170_, _40169_, _40167_);
  nor (_40171_, _40160_, _38417_);
  or (_40172_, _40171_, _40170_);
  and (_42764_, _40172_, _41806_);
  and (_40173_, _30730_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40174_, _40173_, _30719_);
  and (_40175_, _40174_, _39808_);
  nand (_40176_, _39808_, _39426_);
  and (_40177_, _40176_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40178_, _40177_, _39805_);
  or (_40179_, _40178_, _40175_);
  nand (_40180_, _39805_, _38410_);
  and (_40181_, _40180_, _41806_);
  and (_42766_, _40181_, _40179_);
  and (_40182_, _39808_, _31436_);
  nand (_40183_, _40182_, _28676_);
  or (_40184_, _40182_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40185_, _40184_, _40183_);
  or (_40186_, _40185_, _39805_);
  nand (_40187_, _39805_, _38402_);
  and (_40188_, _40187_, _41806_);
  and (_42768_, _40188_, _40186_);
  and (_40189_, _39808_, _32131_);
  nand (_40190_, _40189_, _28676_);
  or (_40191_, _40189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_40192_, _40191_, _40160_);
  and (_40193_, _40192_, _40190_);
  nor (_40194_, _40160_, _38394_);
  or (_40195_, _40194_, _40193_);
  and (_42770_, _40195_, _41806_);
  and (_40196_, _39808_, _32941_);
  nand (_40197_, _40196_, _28676_);
  or (_40198_, _40196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_40199_, _40198_, _40160_);
  and (_40200_, _40199_, _40197_);
  nor (_40201_, _40160_, _38366_);
  or (_40202_, _40201_, _40200_);
  and (_42772_, _40202_, _41806_);
  and (_40203_, _39808_, _33697_);
  nand (_40204_, _40203_, _28676_);
  or (_40205_, _40203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_40206_, _40205_, _40160_);
  and (_40207_, _40206_, _40204_);
  nor (_40208_, _40160_, _38280_);
  or (_40209_, _40208_, _40207_);
  and (_42774_, _40209_, _41806_);
  and (_40210_, _39797_, _24456_);
  nand (_40211_, _40210_, _28676_);
  or (_40212_, _40210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40213_, _40212_, _40211_);
  or (_40214_, _40213_, _39794_);
  nand (_40215_, _39794_, _38425_);
  and (_40216_, _40215_, _41806_);
  and (_42776_, _40216_, _40214_);
  and (_40217_, _39797_, _30002_);
  nand (_40218_, _40217_, _28676_);
  not (_40219_, _39794_);
  or (_40220_, _40217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40221_, _40220_, _40219_);
  and (_40222_, _40221_, _40218_);
  nor (_40223_, _40219_, _38417_);
  or (_40224_, _40223_, _40222_);
  and (_42778_, _40224_, _41806_);
  and (_40225_, _30730_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40226_, _40225_, _30719_);
  and (_40227_, _40226_, _39797_);
  nand (_40228_, _39797_, _39426_);
  and (_40229_, _40228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40230_, _40229_, _39794_);
  or (_40231_, _40230_, _40227_);
  nand (_40232_, _39794_, _38410_);
  and (_40233_, _40232_, _41806_);
  and (_42780_, _40233_, _40231_);
  and (_40234_, _39797_, _31436_);
  nand (_40235_, _40234_, _28676_);
  or (_40236_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40237_, _40236_, _40219_);
  and (_40238_, _40237_, _40235_);
  nor (_40239_, _40219_, _38402_);
  or (_40240_, _40239_, _40238_);
  and (_42782_, _40240_, _41806_);
  and (_40241_, _39797_, _32131_);
  nand (_40242_, _40241_, _28676_);
  or (_40243_, _40241_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40244_, _40243_, _40219_);
  and (_40245_, _40244_, _40242_);
  nor (_40246_, _40219_, _38394_);
  or (_40247_, _40246_, _40245_);
  and (_42784_, _40247_, _41806_);
  and (_40248_, _39797_, _32941_);
  nand (_40249_, _40248_, _28676_);
  or (_40250_, _40248_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40251_, _40250_, _40219_);
  and (_40252_, _40251_, _40249_);
  nor (_40253_, _40219_, _38366_);
  or (_40254_, _40253_, _40252_);
  and (_42786_, _40254_, _41806_);
  and (_40255_, _39797_, _33697_);
  nand (_40256_, _40255_, _28676_);
  or (_40257_, _40255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_40258_, _40257_, _40219_);
  and (_40259_, _40258_, _40256_);
  nor (_40260_, _40219_, _38280_);
  or (_40261_, _40260_, _40259_);
  and (_42788_, _40261_, _41806_);
  nor (_40262_, _24949_, _23932_);
  nor (_40263_, _40262_, _28065_);
  not (_40264_, _40263_);
  and (_40265_, _37954_, _37811_);
  not (_40266_, _38443_);
  and (_40267_, _40266_, _40265_);
  not (_40268_, _40267_);
  not (_40269_, _36836_);
  and (_40270_, _37800_, _40269_);
  and (_40271_, _40270_, _37954_);
  not (_40272_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_40273_, _36409_, _29980_);
  nor (_40274_, _36409_, _29980_);
  nor (_40275_, _40274_, _40273_);
  and (_40276_, _40275_, _24313_);
  not (_40277_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_40278_, _38821_, _40277_);
  nor (_40279_, _40278_, _38908_);
  and (_40280_, _40279_, _25113_);
  nor (_40281_, _40279_, _25113_);
  nor (_40282_, _40281_, _40280_);
  and (_40283_, _40282_, _24197_);
  and (_40284_, _40283_, _40276_);
  and (_40285_, _40284_, _40263_);
  and (_40286_, _40285_, _40272_);
  and (_40287_, _40286_, _38173_);
  and (_40288_, _40279_, _36420_);
  and (_40289_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_40290_, _40279_, _36420_);
  and (_40291_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_40292_, _40291_, _40289_);
  nor (_40293_, _40279_, _36409_);
  and (_40294_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_40295_, _40279_, _36409_);
  and (_40296_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_40297_, _40296_, _40294_);
  and (_40298_, _40297_, _40292_);
  nor (_40299_, _40298_, _40286_);
  nor (_40300_, _40299_, _40287_);
  not (_40301_, _40300_);
  and (_40302_, _40301_, _40271_);
  not (_40303_, _37954_);
  nor (_40304_, _37800_, _40269_);
  not (_40305_, _33860_);
  and (_40306_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_40307_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_40308_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_40309_, _40308_, _40307_);
  and (_40310_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_40311_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_40312_, _40311_, _40310_);
  and (_40313_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_40314_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_40315_, _40314_, _40313_);
  and (_40316_, _40315_, _40312_);
  and (_40317_, _40316_, _40309_);
  nor (_40318_, _33915_, _40305_);
  not (_40319_, _40318_);
  nor (_40320_, _40319_, _40317_);
  nor (_40321_, _40320_, _40306_);
  not (_40322_, _40321_);
  and (_40323_, _40322_, _40304_);
  nor (_40324_, _40323_, _40303_);
  not (_40325_, _40324_);
  nor (_40326_, _40325_, _40302_);
  and (_40327_, _40326_, _40268_);
  nor (_40328_, _37384_, _37148_);
  nor (_40329_, _37296_, _37252_);
  nor (_40330_, _37454_, _37219_);
  and (_40331_, _40330_, _40329_);
  and (_40332_, _37539_, _37351_);
  and (_40333_, _40332_, _40331_);
  and (_40334_, _40333_, _40328_);
  nor (_40335_, _40334_, _33817_);
  and (_40336_, _37507_, _36584_);
  nor (_40337_, _37712_, _40336_);
  nor (_40338_, _40337_, _37679_);
  nor (_40339_, _40338_, _40335_);
  not (_40340_, _40339_);
  and (_40341_, _40340_, _40327_);
  and (_40342_, _40304_, _37954_);
  and (_40343_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_40344_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_40345_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_40346_, _40345_, _40344_);
  and (_40347_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_40348_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_40349_, _40348_, _40347_);
  and (_40350_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_40351_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_40352_, _40351_, _40350_);
  and (_40353_, _40352_, _40349_);
  and (_40354_, _40353_, _40346_);
  nor (_40355_, _40354_, _40319_);
  nor (_40356_, _40355_, _40343_);
  not (_40357_, _40356_);
  and (_40358_, _40357_, _40342_);
  not (_40359_, _40271_);
  not (_40360_, _38402_);
  and (_40361_, _40286_, _40360_);
  and (_40362_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_40363_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_40364_, _40363_, _40362_);
  and (_40365_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_40366_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_40367_, _40366_, _40365_);
  and (_40368_, _40367_, _40364_);
  nor (_40369_, _40368_, _40286_);
  nor (_40370_, _40369_, _40361_);
  nor (_40371_, _40370_, _40359_);
  nor (_40372_, _40371_, _40358_);
  not (_40373_, _38469_);
  and (_40374_, _40373_, _40265_);
  not (_40375_, _40279_);
  and (_40376_, _37800_, _36836_);
  and (_40377_, _40376_, _37954_);
  and (_40378_, _40377_, _40375_);
  nor (_40379_, _40378_, _40374_);
  and (_40380_, _40379_, _40372_);
  not (_40381_, _40380_);
  and (_40382_, _40381_, _40341_);
  and (_40383_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_40384_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_40385_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_40386_, _40385_, _40384_);
  and (_40387_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_40388_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_40389_, _40388_, _40387_);
  and (_40390_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_40391_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_40392_, _40391_, _40390_);
  and (_40393_, _40392_, _40389_);
  and (_40394_, _40393_, _40386_);
  nor (_40395_, _40394_, _40319_);
  nor (_40396_, _40395_, _40383_);
  not (_40397_, _40396_);
  and (_40398_, _40397_, _40342_);
  and (_40399_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_40400_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_40401_, _40400_, _40399_);
  and (_40402_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_40403_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_40404_, _40403_, _40402_);
  and (_40405_, _40404_, _40401_);
  nor (_40406_, _40405_, _40286_);
  and (_40407_, _40286_, _38426_);
  nor (_40408_, _40407_, _40406_);
  nor (_40409_, _40408_, _40359_);
  nor (_40410_, _40409_, _40398_);
  not (_40411_, _38451_);
  and (_40412_, _40411_, _40265_);
  and (_40413_, _40377_, _36420_);
  nor (_40414_, _40413_, _40412_);
  and (_40415_, _40414_, _40410_);
  nor (_40416_, _40415_, _40340_);
  nor (_40417_, _40416_, _40382_);
  and (_40418_, _24949_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40419_, _40418_, _25113_);
  nor (_40420_, _24434_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40421_, _40420_, _40419_);
  not (_40422_, _40421_);
  and (_40423_, _40422_, _40417_);
  nor (_40424_, _40423_, _40264_);
  and (_40425_, _40303_, _36836_);
  and (_40426_, _40425_, _37800_);
  not (_40427_, _38481_);
  and (_40428_, _40427_, _40265_);
  nor (_40429_, _40428_, _40426_);
  and (_40430_, _40303_, _37811_);
  not (_40431_, _40430_);
  not (_40432_, _38366_);
  and (_40433_, _40286_, _40432_);
  and (_40434_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_40435_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_40436_, _40435_, _40434_);
  and (_40437_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_40438_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_40439_, _40438_, _40437_);
  and (_40440_, _40439_, _40436_);
  nor (_40441_, _40440_, _40286_);
  nor (_40442_, _40441_, _40433_);
  not (_40443_, _40442_);
  and (_40444_, _40443_, _40271_);
  and (_40445_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_40446_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_40447_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_40448_, _40447_, _40446_);
  and (_40449_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_40450_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_40451_, _40450_, _40449_);
  and (_40452_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_40453_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_40454_, _40453_, _40452_);
  and (_40455_, _40454_, _40451_);
  and (_40456_, _40455_, _40448_);
  nor (_40457_, _40456_, _40319_);
  nor (_40458_, _40457_, _40445_);
  not (_40459_, _40458_);
  and (_40460_, _40459_, _40342_);
  nor (_40461_, _40460_, _40444_);
  and (_40462_, _40461_, _40431_);
  and (_40463_, _40462_, _40429_);
  not (_40464_, _40463_);
  and (_40465_, _40464_, _40341_);
  and (_40466_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_40467_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_40468_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_40469_, _40468_, _40467_);
  and (_40470_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_40471_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_40472_, _40471_, _40470_);
  and (_40473_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_40474_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_40475_, _40474_, _40473_);
  and (_40476_, _40475_, _40472_);
  and (_40477_, _40476_, _40469_);
  nor (_40478_, _40477_, _40319_);
  nor (_40479_, _40478_, _40466_);
  not (_40480_, _40479_);
  and (_40481_, _40480_, _40342_);
  not (_40482_, _38410_);
  and (_40483_, _40286_, _40482_);
  and (_40484_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_40485_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_40486_, _40485_, _40484_);
  and (_40487_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_40488_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_40489_, _40488_, _40487_);
  and (_40490_, _40489_, _40486_);
  nor (_40491_, _40490_, _40286_);
  nor (_40492_, _40491_, _40483_);
  not (_40493_, _40492_);
  and (_40494_, _40493_, _40271_);
  nor (_40495_, _40494_, _40481_);
  not (_40496_, _38463_);
  and (_40497_, _40496_, _40265_);
  and (_40498_, _40377_, _36869_);
  nor (_40499_, _40498_, _40497_);
  and (_40500_, _40499_, _40495_);
  nor (_40501_, _40500_, _40340_);
  nor (_40502_, _40501_, _40465_);
  and (_40503_, _40418_, _39027_);
  nor (_40504_, _24197_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40505_, _40504_, _40503_);
  not (_40506_, _40505_);
  and (_40507_, _40506_, _40502_);
  nor (_40508_, _40422_, _40417_);
  nor (_40509_, _40508_, _40507_);
  and (_40510_, _40509_, _40424_);
  not (_40511_, _38475_);
  and (_40512_, _40511_, _40265_);
  or (_40513_, _40512_, _40425_);
  and (_40514_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_40515_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_40516_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_40517_, _40516_, _40515_);
  and (_40518_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_40519_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_40520_, _40519_, _40518_);
  and (_40521_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_40522_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_40523_, _40522_, _40521_);
  and (_40524_, _40523_, _40520_);
  and (_40525_, _40524_, _40517_);
  nor (_40526_, _40525_, _40319_);
  nor (_40527_, _40526_, _40514_);
  not (_40528_, _40527_);
  and (_40529_, _40528_, _40342_);
  and (_40530_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_40531_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_40532_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_40533_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_40534_, _40533_, _40532_);
  or (_40535_, _40534_, _40531_);
  nor (_40536_, _40535_, _40530_);
  nor (_40537_, _40536_, _40286_);
  not (_40538_, _38394_);
  and (_40539_, _40286_, _40538_);
  or (_40540_, _40539_, _40537_);
  and (_40541_, _40540_, _40271_);
  or (_40542_, _40541_, _40529_);
  nor (_40543_, _38821_, _38949_);
  or (_40544_, _40543_, _38963_);
  and (_40545_, _40544_, _40377_);
  or (_40546_, _40545_, _40542_);
  or (_40547_, _40546_, _40513_);
  and (_40548_, _40547_, _40341_);
  and (_40549_, _40270_, _40303_);
  not (_40550_, _38457_);
  and (_40551_, _40550_, _40265_);
  nor (_40552_, _40551_, _40549_);
  and (_40553_, _40377_, _36431_);
  and (_40554_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  not (_40555_, _40554_);
  and (_40556_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_40557_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_40558_, _40557_, _40556_);
  and (_40559_, _40558_, _40555_);
  and (_40560_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_40561_, _40560_, _40286_);
  and (_40562_, _40561_, _40559_);
  and (_40563_, _40286_, _38417_);
  or (_40564_, _40563_, _40562_);
  nor (_40570_, _40564_, _40359_);
  and (_40576_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_40582_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_40588_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_40594_, _40588_, _40582_);
  and (_40597_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_40598_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_40599_, _40598_, _40597_);
  and (_40600_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_40601_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_40602_, _40601_, _40600_);
  and (_40603_, _40602_, _40599_);
  and (_40604_, _40603_, _40594_);
  nor (_40605_, _40604_, _40319_);
  nor (_40606_, _40605_, _40576_);
  not (_40607_, _40606_);
  and (_40608_, _40607_, _40342_);
  or (_40609_, _40608_, _40570_);
  nor (_40610_, _40609_, _40553_);
  and (_40611_, _40610_, _40552_);
  nor (_40612_, _40611_, _40340_);
  nor (_40613_, _40612_, _40548_);
  not (_40614_, _25244_);
  and (_40615_, _40418_, _40614_);
  nor (_40616_, _24313_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40617_, _40616_, _40615_);
  nand (_40618_, _40617_, _40613_);
  or (_40619_, _40617_, _40613_);
  and (_40620_, _40619_, _40618_);
  not (_40621_, _40620_);
  nor (_40622_, _40506_, _40502_);
  not (_40623_, _40622_);
  nor (_40624_, _40381_, _40341_);
  and (_40625_, _40290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_40626_, _40288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_40627_, _40626_, _40625_);
  and (_40628_, _40293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_40629_, _40295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_40630_, _40629_, _40628_);
  and (_40631_, _40630_, _40627_);
  nor (_40632_, _40631_, _40286_);
  not (_40633_, _38280_);
  and (_40636_, _40286_, _40633_);
  nor (_40639_, _40636_, _40632_);
  nor (_40643_, _40639_, _40359_);
  and (_40645_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_40646_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_40647_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_40652_, _40647_, _40646_);
  and (_40657_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_40658_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_40659_, _40658_, _40657_);
  and (_40660_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_40666_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_40670_, _40666_, _40660_);
  and (_40671_, _40670_, _40659_);
  and (_40672_, _40671_, _40652_);
  nor (_40677_, _40672_, _40319_);
  nor (_40682_, _40677_, _40645_);
  not (_40683_, _40682_);
  and (_40684_, _40683_, _40304_);
  or (_40685_, _40684_, _40425_);
  nor (_40691_, _40685_, _40643_);
  not (_40695_, _38487_);
  and (_40696_, _40695_, _40265_);
  nor (_40697_, _40696_, _40430_);
  and (_40703_, _40697_, _40691_);
  and (_40707_, _40703_, _40341_);
  nor (_40708_, _40707_, _40624_);
  nor (_40709_, _40418_, _25113_);
  and (_40714_, _40418_, _24665_);
  nor (_40719_, _40714_, _40709_);
  not (_40720_, _40719_);
  and (_40721_, _40720_, _40708_);
  nor (_40726_, _40720_, _40708_);
  nor (_40731_, _40726_, _40721_);
  and (_40732_, _40731_, _40623_);
  and (_40733_, _40732_, _40621_);
  and (_40734_, _40733_, _40510_);
  not (_40740_, _40502_);
  and (_40744_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_40745_, _40417_);
  and (_40746_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_40752_, _40746_, _40744_);
  and (_40756_, _40752_, _40613_);
  not (_40757_, _40613_);
  not (_40758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_40763_, _40417_, _40758_);
  and (_40768_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_40769_, _40768_, _40763_);
  and (_40770_, _40769_, _40757_);
  or (_40775_, _40770_, _40756_);
  or (_40780_, _40775_, _40740_);
  not (_40781_, _40708_);
  and (_40782_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_40785_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_40791_, _40785_, _40782_);
  and (_40793_, _40791_, _40613_);
  not (_40794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_40797_, _40417_, _40794_);
  and (_40803_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_40805_, _40803_, _40797_);
  and (_40806_, _40805_, _40757_);
  or (_40808_, _40806_, _40793_);
  or (_40814_, _40808_, _40502_);
  and (_40817_, _40814_, _40781_);
  and (_40818_, _40817_, _40780_);
  or (_40820_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_40826_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_40828_, _40826_, _40820_);
  and (_40829_, _40828_, _40613_);
  or (_40830_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_40831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_40832_, _40417_, _40831_);
  and (_40833_, _40832_, _40830_);
  and (_40834_, _40833_, _40757_);
  or (_40835_, _40834_, _40829_);
  or (_40836_, _40835_, _40740_);
  or (_40837_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_40838_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_40839_, _40838_, _40837_);
  and (_40840_, _40839_, _40613_);
  or (_40841_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_40842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_40843_, _40417_, _40842_);
  and (_40844_, _40843_, _40841_);
  and (_40845_, _40844_, _40757_);
  or (_40846_, _40845_, _40840_);
  or (_40847_, _40846_, _40502_);
  and (_40848_, _40847_, _40708_);
  and (_40849_, _40848_, _40836_);
  or (_40850_, _40849_, _40818_);
  or (_40851_, _40850_, _40734_);
  not (_40852_, _40734_);
  or (_40853_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_40854_, _40853_, _41806_);
  and (_42863_, _40854_, _40851_);
  nor (_40855_, _40421_, _40264_);
  nor (_40856_, _40617_, _40264_);
  and (_40857_, _40856_, _40855_);
  and (_40858_, _40719_, _40263_);
  nor (_40859_, _40505_, _40264_);
  and (_40860_, _40859_, _40858_);
  and (_40861_, _40860_, _40857_);
  and (_40862_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_40863_, _40862_, _26071_);
  nor (_40864_, _40863_, _28676_);
  nand (_40865_, _26071_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40866_, _17475_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40867_, _40866_, _40865_);
  nor (_40868_, _38162_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_40869_, _40868_, _40867_);
  or (_40870_, _40869_, _40864_);
  and (_40871_, _40870_, _40263_);
  and (_40872_, _40871_, _40861_);
  not (_40873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_40874_, _40861_, _40873_);
  or (_42875_, _40874_, _40872_);
  nor (_40875_, _40859_, _40858_);
  nor (_40876_, _40856_, _40855_);
  and (_40877_, _40876_, _40263_);
  and (_40878_, _40877_, _40875_);
  and (_40879_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _26061_);
  and (_40880_, _40879_, _26104_);
  not (_40881_, _40880_);
  nor (_40882_, _40881_, _28676_);
  not (_40883_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40884_, _38425_, _40883_);
  or (_40885_, _16315_, _40883_);
  and (_40886_, _40885_, _40881_);
  and (_40887_, _40886_, _40884_);
  or (_40888_, _40887_, _40882_);
  and (_40889_, _40888_, _40878_);
  not (_40890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_40891_, _40878_, _40890_);
  or (_43133_, _40891_, _40889_);
  nand (_40892_, _40879_, _26180_);
  nor (_40893_, _40892_, _28676_);
  nor (_40894_, _38417_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40895_, _40879_, _26137_);
  and (_40896_, _40879_, _26071_);
  or (_40897_, _40896_, _40862_);
  or (_40898_, _40897_, _40895_);
  and (_40899_, _40898_, _17301_);
  or (_40900_, _40899_, _40894_);
  or (_40901_, _40900_, _40893_);
  and (_40902_, _40901_, _40878_);
  not (_40903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_40904_, _40878_, _40903_);
  or (_43139_, _40904_, _40902_);
  not (_40905_, _40878_);
  and (_40906_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_40907_, _40879_, _26147_);
  nor (_40908_, _40907_, _28676_);
  nor (_40909_, _38410_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40910_, _40879_, _26169_);
  or (_40911_, _40910_, _40897_);
  and (_40912_, _40911_, _15953_);
  or (_40913_, _40912_, _40909_);
  or (_40914_, _40913_, _40908_);
  and (_40915_, _40914_, _40878_);
  or (_43145_, _40915_, _40906_);
  and (_40916_, _40896_, _29318_);
  nor (_40917_, _38402_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_40918_, _40895_, _40862_);
  or (_40919_, _40918_, _40910_);
  and (_40920_, _40919_, _16985_);
  or (_40921_, _40920_, _40917_);
  or (_40922_, _40921_, _40916_);
  and (_40923_, _40922_, _40878_);
  and (_40924_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_43151_, _40924_, _40923_);
  nand (_40925_, _40862_, _26104_);
  nor (_40926_, _40925_, _28676_);
  nor (_40927_, _38394_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40928_, _26104_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40929_, _16150_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40930_, _40929_, _40928_);
  or (_40931_, _40930_, _40927_);
  or (_40932_, _40931_, _40926_);
  and (_40933_, _40932_, _40878_);
  and (_40934_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_43157_, _40934_, _40933_);
  nand (_40935_, _40862_, _26180_);
  nor (_40936_, _40935_, _28676_);
  nor (_40937_, _38366_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40938_, _26180_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40939_, _17138_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40940_, _40939_, _40938_);
  or (_40941_, _40940_, _40937_);
  or (_40942_, _40941_, _40936_);
  and (_40943_, _40942_, _40878_);
  and (_40944_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_43163_, _40944_, _40943_);
  nand (_40945_, _40862_, _26147_);
  nor (_40946_, _40945_, _28676_);
  nor (_40947_, _38280_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_40948_, _26147_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_40949_, _16490_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40950_, _40949_, _40948_);
  or (_40951_, _40950_, _40947_);
  or (_40952_, _40951_, _40946_);
  and (_40953_, _40952_, _40878_);
  and (_40954_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_43169_, _40954_, _40953_);
  and (_40955_, _40878_, _40870_);
  and (_40956_, _40905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_43172_, _40956_, _40955_);
  and (_40957_, _40888_, _40263_);
  and (_40958_, _40855_, _40617_);
  and (_40959_, _40958_, _40875_);
  and (_40960_, _40959_, _40957_);
  not (_40961_, _40959_);
  and (_40962_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_43180_, _40962_, _40960_);
  and (_40963_, _40901_, _40263_);
  and (_40964_, _40959_, _40963_);
  and (_40965_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_43184_, _40965_, _40964_);
  and (_40966_, _40914_, _40263_);
  and (_40967_, _40959_, _40966_);
  and (_40968_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_43188_, _40968_, _40967_);
  and (_40969_, _40922_, _40263_);
  and (_40970_, _40959_, _40969_);
  and (_40971_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_43192_, _40971_, _40970_);
  and (_40972_, _40932_, _40263_);
  and (_40973_, _40959_, _40972_);
  not (_40974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_40975_, _40959_, _40974_);
  or (_43196_, _40975_, _40973_);
  and (_40976_, _40942_, _40263_);
  and (_40977_, _40959_, _40976_);
  not (_40978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_40979_, _40959_, _40978_);
  or (_43200_, _40979_, _40977_);
  and (_40980_, _40952_, _40263_);
  and (_40981_, _40959_, _40980_);
  and (_40982_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_43204_, _40982_, _40981_);
  and (_40983_, _40959_, _40871_);
  and (_40984_, _40961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_43207_, _40984_, _40983_);
  and (_40985_, _40856_, _40421_);
  and (_40986_, _40985_, _40875_);
  and (_40987_, _40986_, _40957_);
  not (_40988_, _40986_);
  and (_40989_, _40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_43215_, _40989_, _40987_);
  and (_40990_, _40986_, _40963_);
  and (_40991_, _40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_43219_, _40991_, _40990_);
  and (_40992_, _40986_, _40966_);
  not (_40993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_40994_, _40986_, _40993_);
  or (_43223_, _40994_, _40992_);
  and (_40995_, _40986_, _40969_);
  and (_40996_, _40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_43227_, _40996_, _40995_);
  and (_40997_, _40986_, _40972_);
  not (_40998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_40999_, _40986_, _40998_);
  or (_43231_, _40999_, _40997_);
  and (_41000_, _40986_, _40976_);
  not (_41001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_41002_, _40986_, _41001_);
  or (_43235_, _41002_, _41000_);
  and (_41003_, _40986_, _40980_);
  and (_41004_, _40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_43239_, _41004_, _41003_);
  and (_41005_, _40986_, _40871_);
  not (_41006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_41007_, _40986_, _41006_);
  or (_43242_, _41007_, _41005_);
  and (_41008_, _40875_, _40857_);
  and (_41009_, _41008_, _40957_);
  not (_41010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_41011_, _41008_, _41010_);
  or (_43248_, _41011_, _41009_);
  and (_41012_, _41008_, _40963_);
  not (_41013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_41014_, _41008_, _41013_);
  or (_43252_, _41014_, _41012_);
  and (_41015_, _41008_, _40966_);
  not (_41016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_41017_, _41008_, _41016_);
  or (_43256_, _41017_, _41015_);
  and (_41018_, _41008_, _40969_);
  not (_41019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_41020_, _41008_, _41019_);
  or (_43260_, _41020_, _41018_);
  and (_41021_, _41008_, _40972_);
  not (_41022_, _41008_);
  and (_41023_, _41022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_43264_, _41023_, _41021_);
  and (_41024_, _41008_, _40976_);
  and (_41025_, _41022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_43268_, _41025_, _41024_);
  and (_41026_, _41008_, _40980_);
  and (_41027_, _41022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_43272_, _41027_, _41026_);
  and (_41028_, _41008_, _40871_);
  nor (_41029_, _41008_, _40758_);
  or (_43275_, _41029_, _41028_);
  and (_41030_, _40859_, _40720_);
  and (_41031_, _41030_, _40876_);
  and (_41032_, _41031_, _40957_);
  not (_41033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_41034_, _41031_, _41033_);
  or (_43283_, _41034_, _41032_);
  and (_41035_, _41031_, _40963_);
  not (_41036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_41037_, _41031_, _41036_);
  or (_43287_, _41037_, _41035_);
  and (_41038_, _41031_, _40966_);
  not (_41039_, _41031_);
  and (_41040_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_43291_, _41040_, _41038_);
  and (_41041_, _41031_, _40969_);
  not (_41042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_41043_, _41031_, _41042_);
  or (_43295_, _41043_, _41041_);
  and (_41044_, _41031_, _40972_);
  and (_41045_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_43299_, _41045_, _41044_);
  and (_41046_, _41031_, _40976_);
  and (_41047_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_43303_, _41047_, _41046_);
  and (_41048_, _41031_, _40980_);
  and (_41049_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_43307_, _41049_, _41048_);
  and (_41050_, _41031_, _40871_);
  and (_41051_, _41039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_43310_, _41051_, _41050_);
  and (_41052_, _41030_, _40958_);
  and (_41053_, _41052_, _40957_);
  not (_41054_, _41052_);
  and (_41055_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_43315_, _41055_, _41053_);
  and (_41056_, _41052_, _40963_);
  and (_41057_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_43319_, _41057_, _41056_);
  and (_41058_, _41052_, _40966_);
  and (_41059_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_43322_, _41059_, _41058_);
  and (_41060_, _41052_, _40969_);
  and (_41061_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_43326_, _41061_, _41060_);
  and (_41062_, _41052_, _40972_);
  not (_41063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_41064_, _41052_, _41063_);
  or (_43330_, _41064_, _41062_);
  and (_41065_, _41052_, _40976_);
  not (_41066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_41067_, _41052_, _41066_);
  or (_43334_, _41067_, _41065_);
  and (_41068_, _41052_, _40980_);
  not (_41069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_41070_, _41052_, _41069_);
  or (_43338_, _41070_, _41068_);
  and (_41071_, _41052_, _40871_);
  and (_41072_, _41054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_43341_, _41072_, _41071_);
  and (_41073_, _41030_, _40985_);
  and (_41074_, _41073_, _40957_);
  not (_41075_, _41073_);
  and (_41076_, _41075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_43346_, _41076_, _41074_);
  and (_41077_, _41073_, _40963_);
  and (_41078_, _41075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_43350_, _41078_, _41077_);
  and (_41079_, _41073_, _40966_);
  not (_41080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_41081_, _41073_, _41080_);
  or (_43354_, _41081_, _41079_);
  and (_41082_, _41073_, _40969_);
  and (_41083_, _41075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_43358_, _41083_, _41082_);
  and (_41084_, _41073_, _40972_);
  not (_41085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_41086_, _41073_, _41085_);
  or (_43362_, _41086_, _41084_);
  and (_41087_, _41073_, _40976_);
  not (_41088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_41089_, _41073_, _41088_);
  or (_43366_, _41089_, _41087_);
  and (_41090_, _41073_, _40980_);
  not (_41091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_41092_, _41073_, _41091_);
  or (_43370_, _41092_, _41090_);
  and (_41093_, _41073_, _40871_);
  not (_41094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_41095_, _41073_, _41094_);
  or (_43373_, _41095_, _41093_);
  and (_41096_, _41030_, _40857_);
  and (_41097_, _41096_, _40957_);
  not (_41098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_41099_, _41096_, _41098_);
  or (_43378_, _41099_, _41097_);
  and (_41100_, _41096_, _40963_);
  not (_41101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_41102_, _41096_, _41101_);
  or (_43382_, _41102_, _41100_);
  and (_41103_, _41096_, _40966_);
  not (_41104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_41105_, _41096_, _41104_);
  or (_43386_, _41105_, _41103_);
  and (_41106_, _41096_, _40969_);
  not (_41107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_41108_, _41096_, _41107_);
  or (_43390_, _41108_, _41106_);
  and (_41109_, _41096_, _40972_);
  not (_41110_, _41096_);
  and (_41111_, _41110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_43394_, _41111_, _41109_);
  and (_41112_, _41096_, _40976_);
  and (_41113_, _41110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_43398_, _41113_, _41112_);
  and (_41114_, _41096_, _40980_);
  and (_41115_, _41110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_43402_, _41115_, _41114_);
  and (_41116_, _41096_, _40871_);
  nor (_41117_, _41096_, _40794_);
  or (_43405_, _41117_, _41116_);
  and (_41118_, _40858_, _40505_);
  and (_41119_, _41118_, _40876_);
  and (_41120_, _41119_, _40957_);
  not (_41121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_41122_, _41119_, _41121_);
  or (_43413_, _41122_, _41120_);
  and (_41123_, _41119_, _40963_);
  not (_41124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_41125_, _41119_, _41124_);
  or (_43417_, _41125_, _41123_);
  and (_41126_, _41119_, _40966_);
  not (_41127_, _41119_);
  and (_41128_, _41127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_43421_, _41128_, _41126_);
  and (_41129_, _41119_, _40969_);
  not (_41130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_41131_, _41119_, _41130_);
  or (_43425_, _41131_, _41129_);
  and (_41132_, _41119_, _40972_);
  and (_41133_, _41127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_43429_, _41133_, _41132_);
  and (_41134_, _41119_, _40976_);
  and (_41135_, _41127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_43433_, _41135_, _41134_);
  and (_41136_, _41119_, _40980_);
  not (_41137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_41138_, _41119_, _41137_);
  or (_43437_, _41138_, _41136_);
  and (_41139_, _41119_, _40871_);
  and (_41140_, _41127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_43440_, _41140_, _41139_);
  and (_41141_, _41118_, _40958_);
  and (_41142_, _41141_, _40957_);
  not (_41143_, _41141_);
  and (_41144_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_43445_, _41144_, _41142_);
  and (_41145_, _41141_, _40963_);
  and (_41146_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_43449_, _41146_, _41145_);
  and (_41147_, _41141_, _40966_);
  and (_41148_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_43453_, _41148_, _41147_);
  and (_41149_, _41141_, _40969_);
  and (_41150_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_43457_, _41150_, _41149_);
  and (_41151_, _41141_, _40972_);
  not (_41152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_41153_, _41141_, _41152_);
  or (_43461_, _41153_, _41151_);
  and (_41154_, _41141_, _40976_);
  not (_41155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_41156_, _41141_, _41155_);
  or (_43465_, _41156_, _41154_);
  and (_41157_, _41141_, _40980_);
  and (_41158_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_43469_, _41158_, _41157_);
  and (_41159_, _41141_, _40871_);
  and (_41160_, _41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_43472_, _41160_, _41159_);
  and (_41161_, _41118_, _40985_);
  and (_41162_, _41161_, _40957_);
  not (_41163_, _41161_);
  and (_41164_, _41163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_43477_, _41164_, _41162_);
  and (_41165_, _41161_, _40963_);
  and (_41166_, _41163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_43484_, _41166_, _41165_);
  and (_41167_, _41161_, _40966_);
  not (_41168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_41169_, _41161_, _41168_);
  or (_43504_, _41169_, _41167_);
  and (_41170_, _41161_, _40969_);
  not (_41171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_41172_, _41161_, _41171_);
  or (_43524_, _41172_, _41170_);
  and (_41173_, _41161_, _40972_);
  not (_41174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_41175_, _41161_, _41174_);
  or (_43542_, _41175_, _41173_);
  and (_41176_, _41161_, _40976_);
  not (_41177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_41178_, _41161_, _41177_);
  or (_43560_, _41178_, _41176_);
  and (_41179_, _41161_, _40980_);
  not (_41180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_41181_, _41161_, _41180_);
  or (_43578_, _41181_, _41179_);
  and (_41182_, _41161_, _40871_);
  nor (_41183_, _41161_, _40831_);
  or (_43593_, _41183_, _41182_);
  and (_41184_, _41118_, _40857_);
  and (_41185_, _41184_, _40957_);
  not (_41186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_41187_, _41184_, _41186_);
  or (_43617_, _41187_, _41185_);
  and (_41188_, _41184_, _40963_);
  not (_41189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_41190_, _41184_, _41189_);
  or (_43637_, _41190_, _41188_);
  and (_41191_, _41184_, _40966_);
  not (_41192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_41193_, _41184_, _41192_);
  or (_43657_, _41193_, _41191_);
  and (_41194_, _41184_, _40969_);
  not (_41195_, _41184_);
  and (_41196_, _41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_43669_, _41196_, _41194_);
  and (_41197_, _41184_, _40972_);
  and (_41198_, _41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_43694_, _41198_, _41197_);
  and (_41199_, _41184_, _40976_);
  and (_41200_, _41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_43712_, _41200_, _41199_);
  and (_41201_, _41184_, _40980_);
  and (_41202_, _41195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_43723_, _41202_, _41201_);
  and (_41203_, _41184_, _40871_);
  not (_41204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_41205_, _41184_, _41204_);
  or (_43726_, _41205_, _41203_);
  and (_41206_, _40876_, _40860_);
  and (_41208_, _41206_, _40957_);
  not (_41210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_41212_, _41206_, _41210_);
  or (_43732_, _41212_, _41208_);
  and (_41215_, _41206_, _40963_);
  not (_41217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_41219_, _41206_, _41217_);
  or (_43736_, _41219_, _41215_);
  and (_41222_, _41206_, _40966_);
  not (_41224_, _41206_);
  and (_41226_, _41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_43740_, _41226_, _41222_);
  and (_41229_, _41206_, _40969_);
  not (_41231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_41233_, _41206_, _41231_);
  or (_43744_, _41233_, _41229_);
  and (_41236_, _41206_, _40972_);
  and (_41238_, _41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_43748_, _41238_, _41236_);
  and (_41241_, _41206_, _40976_);
  and (_41243_, _41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_43752_, _41243_, _41241_);
  and (_41246_, _41206_, _40980_);
  not (_41248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_41250_, _41206_, _41248_);
  or (_43756_, _41250_, _41246_);
  and (_41253_, _41206_, _40871_);
  and (_41255_, _41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_43759_, _41255_, _41253_);
  and (_41256_, _40958_, _40860_);
  and (_41257_, _41256_, _40957_);
  not (_41258_, _41256_);
  and (_41259_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_43764_, _41259_, _41257_);
  and (_41260_, _41256_, _40963_);
  and (_41261_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_43768_, _41261_, _41260_);
  and (_41262_, _41256_, _40966_);
  and (_41263_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_43772_, _41263_, _41262_);
  and (_41264_, _41256_, _40969_);
  and (_41265_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_43776_, _41265_, _41264_);
  and (_41266_, _41256_, _40972_);
  not (_41267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_41268_, _41256_, _41267_);
  or (_43780_, _41268_, _41266_);
  and (_41269_, _41256_, _40976_);
  not (_41270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_41271_, _41256_, _41270_);
  or (_43784_, _41271_, _41269_);
  and (_41272_, _41256_, _40980_);
  and (_41273_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_43788_, _41273_, _41272_);
  and (_41274_, _41256_, _40871_);
  and (_41275_, _41258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_43791_, _41275_, _41274_);
  and (_41276_, _40985_, _40860_);
  and (_41277_, _41276_, _40957_);
  not (_41278_, _41276_);
  and (_41279_, _41278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_43796_, _41279_, _41277_);
  and (_41280_, _41276_, _40963_);
  and (_41281_, _41278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_43800_, _41281_, _41280_);
  and (_41282_, _41276_, _40966_);
  not (_41283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_41284_, _41276_, _41283_);
  or (_43804_, _41284_, _41282_);
  and (_41285_, _41276_, _40969_);
  not (_41286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_41287_, _41276_, _41286_);
  or (_43808_, _41287_, _41285_);
  and (_41288_, _41276_, _40972_);
  not (_41289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_41290_, _41276_, _41289_);
  or (_43812_, _41290_, _41288_);
  and (_41291_, _41276_, _40976_);
  not (_41292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_41293_, _41276_, _41292_);
  or (_43816_, _41293_, _41291_);
  and (_41294_, _41276_, _40980_);
  not (_41295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_41296_, _41276_, _41295_);
  or (_43820_, _41296_, _41294_);
  and (_41297_, _41276_, _40871_);
  nor (_41298_, _41276_, _40842_);
  or (_43823_, _41298_, _41297_);
  and (_41299_, _40957_, _40861_);
  not (_41300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_41301_, _40861_, _41300_);
  or (_43826_, _41301_, _41299_);
  and (_41302_, _40963_, _40861_);
  not (_41303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_41304_, _40861_, _41303_);
  or (_43829_, _41304_, _41302_);
  and (_41305_, _40966_, _40861_);
  not (_41306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_41307_, _40861_, _41306_);
  or (_43833_, _41307_, _41305_);
  and (_41308_, _40969_, _40861_);
  not (_41309_, _40861_);
  and (_41310_, _41309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_43837_, _41310_, _41308_);
  and (_41311_, _40972_, _40861_);
  and (_41312_, _41309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_43841_, _41312_, _41311_);
  and (_41313_, _40976_, _40861_);
  and (_41314_, _41309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_43844_, _41314_, _41313_);
  and (_41315_, _40980_, _40861_);
  and (_41316_, _41309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_43847_, _41316_, _41315_);
  or (_41317_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_41318_, _40417_, _40890_);
  and (_41319_, _41318_, _40613_);
  and (_41320_, _41319_, _41317_);
  nor (_41321_, _40417_, _41010_);
  and (_41322_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_41323_, _41322_, _41321_);
  and (_41324_, _41323_, _40757_);
  or (_41325_, _41324_, _41320_);
  or (_41326_, _41325_, _40740_);
  or (_41327_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_41328_, _40417_, _41033_);
  and (_41329_, _41328_, _40613_);
  and (_41330_, _41329_, _41327_);
  nor (_41331_, _40417_, _41098_);
  and (_41332_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_41333_, _41332_, _41331_);
  and (_41334_, _41333_, _40757_);
  or (_41335_, _41334_, _41330_);
  or (_41336_, _41335_, _40502_);
  and (_41337_, _41336_, _40781_);
  and (_41338_, _41337_, _41326_);
  nand (_41339_, _40417_, _41121_);
  or (_41340_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_41341_, _41340_, _41339_);
  and (_41342_, _41341_, _40613_);
  and (_41343_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_41344_, _40417_, _41186_);
  or (_41345_, _41344_, _41343_);
  and (_41346_, _41345_, _40757_);
  or (_41347_, _41346_, _41342_);
  or (_41348_, _41347_, _40740_);
  nand (_41349_, _40417_, _41210_);
  or (_41350_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_41351_, _41350_, _41349_);
  and (_41352_, _41351_, _40613_);
  and (_41353_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_41354_, _40417_, _41300_);
  or (_41355_, _41354_, _41353_);
  and (_41356_, _41355_, _40757_);
  or (_41357_, _41356_, _41352_);
  or (_41358_, _41357_, _40502_);
  and (_41359_, _41358_, _40708_);
  and (_41360_, _41359_, _41348_);
  or (_41361_, _41360_, _41338_);
  or (_41362_, _41361_, _40734_);
  or (_41363_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_41364_, _41363_, _41806_);
  and (_01406_, _41364_, _41362_);
  or (_41365_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_41366_, _40417_, _40903_);
  and (_41367_, _41366_, _40613_);
  and (_41368_, _41367_, _41365_);
  nor (_41369_, _40417_, _41013_);
  and (_41370_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_41371_, _41370_, _41369_);
  and (_41372_, _41371_, _40757_);
  or (_41373_, _41372_, _41368_);
  or (_41374_, _41373_, _40740_);
  or (_41375_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_41376_, _40417_, _41036_);
  and (_41377_, _41376_, _40613_);
  and (_41378_, _41377_, _41375_);
  nor (_41379_, _40417_, _41101_);
  and (_41380_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_41381_, _41380_, _41379_);
  and (_41382_, _41381_, _40757_);
  or (_41383_, _41382_, _41378_);
  or (_41384_, _41383_, _40502_);
  and (_41385_, _41384_, _40781_);
  and (_41386_, _41385_, _41374_);
  nand (_41387_, _40417_, _41124_);
  or (_41388_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_41389_, _41388_, _41387_);
  and (_41390_, _41389_, _40613_);
  and (_41391_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_41392_, _40417_, _41189_);
  or (_41393_, _41392_, _41391_);
  and (_41394_, _41393_, _40757_);
  or (_41395_, _41394_, _41390_);
  or (_41396_, _41395_, _40740_);
  nand (_41397_, _40417_, _41217_);
  or (_41398_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_41399_, _41398_, _41397_);
  and (_41400_, _41399_, _40613_);
  and (_41401_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_41402_, _40417_, _41303_);
  or (_41403_, _41402_, _41401_);
  and (_41404_, _41403_, _40757_);
  or (_41405_, _41404_, _41400_);
  or (_41406_, _41405_, _40502_);
  and (_41407_, _41406_, _40708_);
  and (_41408_, _41407_, _41396_);
  or (_41409_, _41408_, _41386_);
  or (_41410_, _41409_, _40734_);
  or (_41411_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_41412_, _41411_, _41806_);
  and (_01408_, _41412_, _41410_);
  and (_41413_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_41414_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_41415_, _41414_, _41413_);
  and (_41416_, _41415_, _40613_);
  nor (_41417_, _40417_, _41016_);
  and (_41418_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_41419_, _41418_, _41417_);
  and (_41420_, _41419_, _40757_);
  or (_41421_, _41420_, _41416_);
  or (_41422_, _41421_, _40740_);
  and (_41423_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_41424_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_41425_, _41424_, _41423_);
  and (_41426_, _41425_, _40613_);
  nor (_41427_, _40417_, _41104_);
  and (_41428_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_41429_, _41428_, _41427_);
  and (_41430_, _41429_, _40757_);
  or (_41431_, _41430_, _41426_);
  or (_41432_, _41431_, _40502_);
  and (_41433_, _41432_, _40781_);
  and (_41434_, _41433_, _41422_);
  or (_41435_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_41436_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_41437_, _41436_, _41435_);
  and (_41438_, _41437_, _40613_);
  or (_41439_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_41440_, _40417_, _41168_);
  and (_41441_, _41440_, _41439_);
  and (_41442_, _41441_, _40757_);
  or (_41443_, _41442_, _41438_);
  or (_41444_, _41443_, _40740_);
  or (_41445_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_41446_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_41447_, _41446_, _41445_);
  and (_41448_, _41447_, _40613_);
  or (_41449_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_41450_, _40417_, _41283_);
  and (_41451_, _41450_, _41449_);
  and (_41452_, _41451_, _40757_);
  or (_41453_, _41452_, _41448_);
  or (_41454_, _41453_, _40502_);
  and (_41455_, _41454_, _40708_);
  and (_41456_, _41455_, _41444_);
  or (_41457_, _41456_, _41434_);
  or (_41458_, _41457_, _40734_);
  or (_41459_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_41460_, _41459_, _41806_);
  and (_01410_, _41460_, _41458_);
  and (_41461_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_41462_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_41463_, _41462_, _41461_);
  and (_41464_, _41463_, _40613_);
  nor (_41465_, _40417_, _41019_);
  and (_41466_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_41467_, _41466_, _41465_);
  and (_41468_, _41467_, _40757_);
  or (_41469_, _41468_, _41464_);
  or (_41470_, _41469_, _40740_);
  or (_41471_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nand (_41472_, _40417_, _41042_);
  and (_41473_, _41472_, _40613_);
  and (_41474_, _41473_, _41471_);
  nor (_41475_, _40417_, _41107_);
  and (_41476_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_41477_, _41476_, _41475_);
  and (_41478_, _41477_, _40757_);
  or (_41479_, _41478_, _41474_);
  or (_41480_, _41479_, _40502_);
  and (_41481_, _41480_, _40781_);
  and (_41482_, _41481_, _41470_);
  nand (_41483_, _40417_, _41130_);
  or (_41484_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_41485_, _41484_, _41483_);
  and (_41486_, _41485_, _40613_);
  or (_41487_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_41488_, _40417_, _41171_);
  and (_41489_, _41488_, _41487_);
  and (_41490_, _41489_, _40757_);
  or (_41491_, _41490_, _41486_);
  or (_41492_, _41491_, _40740_);
  nand (_41493_, _40417_, _41231_);
  or (_41494_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_41495_, _41494_, _41493_);
  and (_41496_, _41495_, _40613_);
  or (_41497_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_41498_, _40417_, _41286_);
  and (_41499_, _41498_, _41497_);
  and (_41500_, _41499_, _40757_);
  or (_41501_, _41500_, _41496_);
  or (_41502_, _41501_, _40502_);
  and (_41503_, _41502_, _40708_);
  and (_41504_, _41503_, _41492_);
  or (_41505_, _41504_, _41482_);
  or (_41506_, _41505_, _40734_);
  or (_41507_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_41508_, _41507_, _41806_);
  and (_01412_, _41508_, _41506_);
  and (_41509_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_41510_, _40417_, _40974_);
  or (_41511_, _41510_, _41509_);
  and (_41512_, _41511_, _40613_);
  or (_41513_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_41514_, _40417_, _40998_);
  and (_41515_, _41514_, _41513_);
  and (_41516_, _41515_, _40757_);
  or (_41517_, _41516_, _41512_);
  or (_41518_, _41517_, _40740_);
  and (_41519_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_41520_, _40417_, _41063_);
  or (_41521_, _41520_, _41519_);
  and (_41522_, _41521_, _40613_);
  or (_41523_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_41524_, _40417_, _41085_);
  and (_41525_, _41524_, _41523_);
  and (_41526_, _41525_, _40757_);
  or (_41527_, _41526_, _41522_);
  or (_41528_, _41527_, _40502_);
  and (_41529_, _41528_, _40781_);
  and (_41530_, _41529_, _41518_);
  and (_41531_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_41532_, _40417_, _41152_);
  or (_41533_, _41532_, _41531_);
  and (_41534_, _41533_, _40613_);
  or (_41535_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_41536_, _40417_, _41174_);
  and (_41537_, _41536_, _41535_);
  and (_41538_, _41537_, _40757_);
  or (_41539_, _41538_, _41534_);
  or (_41540_, _41539_, _40740_);
  and (_41541_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_41542_, _40417_, _41267_);
  or (_41543_, _41542_, _41541_);
  and (_41544_, _41543_, _40613_);
  or (_41545_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_41546_, _40417_, _41289_);
  and (_41547_, _41546_, _41545_);
  and (_41548_, _41547_, _40757_);
  or (_41549_, _41548_, _41544_);
  or (_41550_, _41549_, _40502_);
  and (_41551_, _41550_, _40708_);
  and (_41552_, _41551_, _41540_);
  or (_41553_, _41552_, _41530_);
  or (_41554_, _41553_, _40734_);
  or (_41555_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_41556_, _41555_, _41806_);
  and (_01414_, _41556_, _41554_);
  and (_41557_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_41558_, _40417_, _40978_);
  or (_41559_, _41558_, _41557_);
  and (_41560_, _41559_, _40613_);
  or (_41561_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_41562_, _40417_, _41001_);
  and (_41563_, _41562_, _41561_);
  and (_41564_, _41563_, _40757_);
  or (_41565_, _41564_, _41560_);
  or (_41566_, _41565_, _40740_);
  and (_41567_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_41568_, _40417_, _41066_);
  or (_41569_, _41568_, _41567_);
  and (_41570_, _41569_, _40613_);
  or (_41571_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_41572_, _40417_, _41088_);
  and (_41573_, _41572_, _41571_);
  and (_41574_, _41573_, _40757_);
  or (_41575_, _41574_, _41570_);
  or (_41576_, _41575_, _40502_);
  and (_41577_, _41576_, _40781_);
  and (_41578_, _41577_, _41566_);
  and (_41579_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_41580_, _40417_, _41155_);
  or (_41581_, _41580_, _41579_);
  and (_41582_, _41581_, _40613_);
  or (_41583_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_41584_, _40417_, _41177_);
  and (_41585_, _41584_, _41583_);
  and (_41586_, _41585_, _40757_);
  or (_41587_, _41586_, _41582_);
  or (_41588_, _41587_, _40740_);
  and (_41589_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_41590_, _40417_, _41270_);
  or (_41591_, _41590_, _41589_);
  and (_41592_, _41591_, _40613_);
  or (_41593_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_41594_, _40417_, _41292_);
  and (_41595_, _41594_, _41593_);
  and (_41596_, _41595_, _40757_);
  or (_41597_, _41596_, _41592_);
  or (_41598_, _41597_, _40502_);
  and (_41599_, _41598_, _40708_);
  and (_41600_, _41599_, _41588_);
  or (_41601_, _41600_, _41578_);
  or (_41602_, _41601_, _40734_);
  or (_41603_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_41604_, _41603_, _41806_);
  and (_01416_, _41604_, _41602_);
  and (_41605_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_41606_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_41607_, _41606_, _41605_);
  and (_41608_, _41607_, _40613_);
  and (_41609_, _40745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_41610_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_41611_, _41610_, _41609_);
  and (_41612_, _41611_, _40757_);
  or (_41613_, _41612_, _41608_);
  or (_41614_, _41613_, _40740_);
  and (_41615_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_41616_, _40417_, _41069_);
  or (_41617_, _41616_, _41615_);
  and (_41618_, _41617_, _40613_);
  or (_41619_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nand (_41620_, _40417_, _41091_);
  and (_41621_, _41620_, _41619_);
  and (_41622_, _41621_, _40757_);
  or (_41623_, _41622_, _41618_);
  or (_41624_, _41623_, _40502_);
  and (_41625_, _41624_, _40781_);
  and (_41626_, _41625_, _41614_);
  nand (_41627_, _40417_, _41137_);
  or (_41628_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_41629_, _41628_, _41627_);
  and (_41630_, _41629_, _40613_);
  or (_41631_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_41632_, _40417_, _41180_);
  and (_41633_, _41632_, _41631_);
  and (_41634_, _41633_, _40757_);
  or (_41635_, _41634_, _41630_);
  or (_41636_, _41635_, _40740_);
  nand (_41637_, _40417_, _41248_);
  or (_41638_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_41639_, _41638_, _41637_);
  and (_41640_, _41639_, _40613_);
  or (_41641_, _40417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_41642_, _40417_, _41295_);
  and (_41643_, _41642_, _41641_);
  and (_41644_, _41643_, _40757_);
  or (_41645_, _41644_, _41640_);
  or (_41646_, _41645_, _40502_);
  and (_41647_, _41646_, _40708_);
  and (_41648_, _41647_, _41636_);
  or (_41649_, _41648_, _41626_);
  or (_41650_, _41649_, _40734_);
  or (_41651_, _40852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_41652_, _41651_, _41806_);
  and (_01418_, _41652_, _41650_);
  or (_41653_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_41654_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_41655_, _41654_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_41656_, _41655_, _41653_);
  nand (_41657_, _41656_, _41806_);
  or (_41658_, \oc8051_gm_cxrom_1.cell0.data [7], _41806_);
  and (_01426_, _41658_, _41657_);
  or (_41659_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41660_, \oc8051_gm_cxrom_1.cell0.data [0], _41654_);
  nand (_41661_, _41660_, _41659_);
  nand (_41662_, _41661_, _41806_);
  or (_41663_, \oc8051_gm_cxrom_1.cell0.data [0], _41806_);
  and (_01433_, _41663_, _41662_);
  or (_41664_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41665_, \oc8051_gm_cxrom_1.cell0.data [1], _41654_);
  nand (_41666_, _41665_, _41664_);
  nand (_41667_, _41666_, _41806_);
  or (_41668_, \oc8051_gm_cxrom_1.cell0.data [1], _41806_);
  and (_01437_, _41668_, _41667_);
  or (_41669_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41670_, \oc8051_gm_cxrom_1.cell0.data [2], _41654_);
  nand (_41671_, _41670_, _41669_);
  nand (_41672_, _41671_, _41806_);
  or (_41673_, \oc8051_gm_cxrom_1.cell0.data [2], _41806_);
  and (_01441_, _41673_, _41672_);
  or (_41674_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41675_, \oc8051_gm_cxrom_1.cell0.data [3], _41654_);
  nand (_41676_, _41675_, _41674_);
  nand (_41677_, _41676_, _41806_);
  or (_41678_, \oc8051_gm_cxrom_1.cell0.data [3], _41806_);
  and (_01444_, _41678_, _41677_);
  or (_41679_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41680_, \oc8051_gm_cxrom_1.cell0.data [4], _41654_);
  nand (_41681_, _41680_, _41679_);
  nand (_41682_, _41681_, _41806_);
  or (_41683_, \oc8051_gm_cxrom_1.cell0.data [4], _41806_);
  and (_01448_, _41683_, _41682_);
  or (_41684_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41685_, \oc8051_gm_cxrom_1.cell0.data [5], _41654_);
  nand (_41686_, _41685_, _41684_);
  nand (_41687_, _41686_, _41806_);
  or (_41688_, \oc8051_gm_cxrom_1.cell0.data [5], _41806_);
  and (_01452_, _41688_, _41687_);
  or (_41689_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41690_, \oc8051_gm_cxrom_1.cell0.data [6], _41654_);
  nand (_41691_, _41690_, _41689_);
  nand (_41692_, _41691_, _41806_);
  or (_41693_, \oc8051_gm_cxrom_1.cell0.data [6], _41806_);
  and (_01456_, _41693_, _41692_);
  or (_41694_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_41695_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_41696_, _41695_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_41697_, _41696_, _41694_);
  nand (_41698_, _41697_, _41806_);
  or (_41699_, \oc8051_gm_cxrom_1.cell1.data [7], _41806_);
  and (_01477_, _41699_, _41698_);
  or (_41700_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41701_, \oc8051_gm_cxrom_1.cell1.data [0], _41695_);
  nand (_41702_, _41701_, _41700_);
  nand (_41703_, _41702_, _41806_);
  or (_41704_, \oc8051_gm_cxrom_1.cell1.data [0], _41806_);
  and (_01484_, _41704_, _41703_);
  or (_41705_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41706_, \oc8051_gm_cxrom_1.cell1.data [1], _41695_);
  nand (_41707_, _41706_, _41705_);
  nand (_41708_, _41707_, _41806_);
  or (_41709_, \oc8051_gm_cxrom_1.cell1.data [1], _41806_);
  and (_01488_, _41709_, _41708_);
  or (_41710_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41711_, \oc8051_gm_cxrom_1.cell1.data [2], _41695_);
  nand (_41712_, _41711_, _41710_);
  nand (_41713_, _41712_, _41806_);
  or (_41714_, \oc8051_gm_cxrom_1.cell1.data [2], _41806_);
  and (_01492_, _41714_, _41713_);
  or (_41715_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41716_, \oc8051_gm_cxrom_1.cell1.data [3], _41695_);
  nand (_41717_, _41716_, _41715_);
  nand (_41718_, _41717_, _41806_);
  or (_41719_, \oc8051_gm_cxrom_1.cell1.data [3], _41806_);
  and (_01496_, _41719_, _41718_);
  or (_41720_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41721_, \oc8051_gm_cxrom_1.cell1.data [4], _41695_);
  nand (_41722_, _41721_, _41720_);
  nand (_41723_, _41722_, _41806_);
  or (_41724_, \oc8051_gm_cxrom_1.cell1.data [4], _41806_);
  and (_01500_, _41724_, _41723_);
  or (_41725_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41726_, \oc8051_gm_cxrom_1.cell1.data [5], _41695_);
  nand (_41727_, _41726_, _41725_);
  nand (_41728_, _41727_, _41806_);
  or (_41729_, \oc8051_gm_cxrom_1.cell1.data [5], _41806_);
  and (_01504_, _41729_, _41728_);
  or (_41730_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41731_, \oc8051_gm_cxrom_1.cell1.data [6], _41695_);
  nand (_41732_, _41731_, _41730_);
  nand (_41733_, _41732_, _41806_);
  or (_41734_, \oc8051_gm_cxrom_1.cell1.data [6], _41806_);
  and (_01508_, _41734_, _41733_);
  or (_41735_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_41736_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_41737_, _41736_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_41738_, _41737_, _41735_);
  nand (_41739_, _41738_, _41806_);
  or (_41740_, \oc8051_gm_cxrom_1.cell2.data [7], _41806_);
  and (_01529_, _41740_, _41739_);
  or (_41741_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41742_, \oc8051_gm_cxrom_1.cell2.data [0], _41736_);
  nand (_41743_, _41742_, _41741_);
  nand (_41744_, _41743_, _41806_);
  or (_41745_, \oc8051_gm_cxrom_1.cell2.data [0], _41806_);
  and (_01536_, _41745_, _41744_);
  or (_41746_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41747_, \oc8051_gm_cxrom_1.cell2.data [1], _41736_);
  nand (_41749_, _41747_, _41746_);
  nand (_41750_, _41749_, _41806_);
  or (_41752_, \oc8051_gm_cxrom_1.cell2.data [1], _41806_);
  and (_01540_, _41752_, _41750_);
  or (_41754_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41756_, \oc8051_gm_cxrom_1.cell2.data [2], _41736_);
  nand (_41758_, _41756_, _41754_);
  nand (_41760_, _41758_, _41806_);
  or (_41762_, \oc8051_gm_cxrom_1.cell2.data [2], _41806_);
  and (_01544_, _41762_, _41760_);
  or (_41763_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41764_, \oc8051_gm_cxrom_1.cell2.data [3], _41736_);
  nand (_41765_, _41764_, _41763_);
  nand (_41766_, _41765_, _41806_);
  or (_41767_, \oc8051_gm_cxrom_1.cell2.data [3], _41806_);
  and (_01548_, _41767_, _41766_);
  or (_41768_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41769_, \oc8051_gm_cxrom_1.cell2.data [4], _41736_);
  nand (_41770_, _41769_, _41768_);
  nand (_41771_, _41770_, _41806_);
  or (_41772_, \oc8051_gm_cxrom_1.cell2.data [4], _41806_);
  and (_01552_, _41772_, _41771_);
  or (_41773_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41774_, \oc8051_gm_cxrom_1.cell2.data [5], _41736_);
  nand (_41775_, _41774_, _41773_);
  nand (_41776_, _41775_, _41806_);
  or (_41777_, \oc8051_gm_cxrom_1.cell2.data [5], _41806_);
  and (_01555_, _41777_, _41776_);
  or (_41778_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41779_, \oc8051_gm_cxrom_1.cell2.data [6], _41736_);
  nand (_41780_, _41779_, _41778_);
  nand (_41781_, _41780_, _41806_);
  or (_41782_, \oc8051_gm_cxrom_1.cell2.data [6], _41806_);
  and (_01559_, _41782_, _41781_);
  or (_41783_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_41784_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_41785_, _41784_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_41786_, _41785_, _41783_);
  nand (_41787_, _41786_, _41806_);
  or (_41788_, \oc8051_gm_cxrom_1.cell3.data [7], _41806_);
  and (_01581_, _41788_, _41787_);
  or (_41789_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41790_, \oc8051_gm_cxrom_1.cell3.data [0], _41784_);
  nand (_41791_, _41790_, _41789_);
  nand (_41792_, _41791_, _41806_);
  or (_41794_, \oc8051_gm_cxrom_1.cell3.data [0], _41806_);
  and (_01588_, _41794_, _41792_);
  or (_41797_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41799_, \oc8051_gm_cxrom_1.cell3.data [1], _41784_);
  nand (_41801_, _41799_, _41797_);
  nand (_41803_, _41801_, _41806_);
  or (_41805_, \oc8051_gm_cxrom_1.cell3.data [1], _41806_);
  and (_01591_, _41805_, _41803_);
  or (_41807_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41808_, \oc8051_gm_cxrom_1.cell3.data [2], _41784_);
  nand (_41809_, _41808_, _41807_);
  nand (_41810_, _41809_, _41806_);
  or (_41811_, \oc8051_gm_cxrom_1.cell3.data [2], _41806_);
  and (_01595_, _41811_, _41810_);
  or (_41812_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41813_, \oc8051_gm_cxrom_1.cell3.data [3], _41784_);
  nand (_41814_, _41813_, _41812_);
  nand (_41815_, _41814_, _41806_);
  or (_41816_, \oc8051_gm_cxrom_1.cell3.data [3], _41806_);
  and (_01599_, _41816_, _41815_);
  or (_41817_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41818_, \oc8051_gm_cxrom_1.cell3.data [4], _41784_);
  nand (_41819_, _41818_, _41817_);
  nand (_41820_, _41819_, _41806_);
  or (_41821_, \oc8051_gm_cxrom_1.cell3.data [4], _41806_);
  and (_01603_, _41821_, _41820_);
  or (_41822_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41823_, \oc8051_gm_cxrom_1.cell3.data [5], _41784_);
  nand (_41824_, _41823_, _41822_);
  nand (_41825_, _41824_, _41806_);
  or (_41826_, \oc8051_gm_cxrom_1.cell3.data [5], _41806_);
  and (_01607_, _41826_, _41825_);
  or (_41827_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_41828_, \oc8051_gm_cxrom_1.cell3.data [6], _41784_);
  nand (_41829_, _41828_, _41827_);
  nand (_41830_, _41829_, _41806_);
  or (_41831_, \oc8051_gm_cxrom_1.cell3.data [6], _41806_);
  and (_01611_, _41831_, _41830_);
  or (_41832_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_41833_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_41834_, _41833_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_41835_, _41834_, _41832_);
  nand (_41836_, _41835_, _41806_);
  or (_41837_, \oc8051_gm_cxrom_1.cell4.data [7], _41806_);
  and (_01628_, _41837_, _41836_);
  or (_41838_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41839_, \oc8051_gm_cxrom_1.cell4.data [0], _41833_);
  nand (_41840_, _41839_, _41838_);
  nand (_41841_, _41840_, _41806_);
  or (_41842_, \oc8051_gm_cxrom_1.cell4.data [0], _41806_);
  and (_01630_, _41842_, _41841_);
  or (_41843_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41844_, \oc8051_gm_cxrom_1.cell4.data [1], _41833_);
  nand (_41845_, _41844_, _41843_);
  nand (_41846_, _41845_, _41806_);
  or (_41847_, \oc8051_gm_cxrom_1.cell4.data [1], _41806_);
  and (_01631_, _41847_, _41846_);
  or (_41848_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41849_, \oc8051_gm_cxrom_1.cell4.data [2], _41833_);
  nand (_41850_, _41849_, _41848_);
  nand (_41851_, _41850_, _41806_);
  or (_41852_, \oc8051_gm_cxrom_1.cell4.data [2], _41806_);
  and (_01634_, _41852_, _41851_);
  or (_41853_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41854_, \oc8051_gm_cxrom_1.cell4.data [3], _41833_);
  nand (_41855_, _41854_, _41853_);
  nand (_41856_, _41855_, _41806_);
  or (_41857_, \oc8051_gm_cxrom_1.cell4.data [3], _41806_);
  and (_01638_, _41857_, _41856_);
  or (_41858_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41859_, \oc8051_gm_cxrom_1.cell4.data [4], _41833_);
  nand (_41860_, _41859_, _41858_);
  nand (_41861_, _41860_, _41806_);
  or (_41862_, \oc8051_gm_cxrom_1.cell4.data [4], _41806_);
  and (_01642_, _41862_, _41861_);
  or (_41863_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41864_, \oc8051_gm_cxrom_1.cell4.data [5], _41833_);
  nand (_41865_, _41864_, _41863_);
  nand (_41866_, _41865_, _41806_);
  or (_41867_, \oc8051_gm_cxrom_1.cell4.data [5], _41806_);
  and (_01646_, _41867_, _41866_);
  or (_41868_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_41869_, \oc8051_gm_cxrom_1.cell4.data [6], _41833_);
  nand (_41870_, _41869_, _41868_);
  nand (_41871_, _41870_, _41806_);
  or (_41872_, \oc8051_gm_cxrom_1.cell4.data [6], _41806_);
  and (_01650_, _41872_, _41871_);
  or (_41873_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_41874_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_41875_, _41874_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_41876_, _41875_, _41873_);
  nand (_41877_, _41876_, _41806_);
  or (_41878_, \oc8051_gm_cxrom_1.cell5.data [7], _41806_);
  and (_01672_, _41878_, _41877_);
  or (_41879_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41880_, \oc8051_gm_cxrom_1.cell5.data [0], _41874_);
  nand (_41881_, _41880_, _41879_);
  nand (_41882_, _41881_, _41806_);
  or (_41883_, \oc8051_gm_cxrom_1.cell5.data [0], _41806_);
  and (_01679_, _41883_, _41882_);
  or (_41884_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41885_, \oc8051_gm_cxrom_1.cell5.data [1], _41874_);
  nand (_41886_, _41885_, _41884_);
  nand (_41887_, _41886_, _41806_);
  or (_41888_, \oc8051_gm_cxrom_1.cell5.data [1], _41806_);
  and (_01683_, _41888_, _41887_);
  or (_41889_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41890_, \oc8051_gm_cxrom_1.cell5.data [2], _41874_);
  nand (_41891_, _41890_, _41889_);
  nand (_41892_, _41891_, _41806_);
  or (_41893_, \oc8051_gm_cxrom_1.cell5.data [2], _41806_);
  and (_01687_, _41893_, _41892_);
  or (_41894_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41895_, \oc8051_gm_cxrom_1.cell5.data [3], _41874_);
  nand (_41896_, _41895_, _41894_);
  nand (_41897_, _41896_, _41806_);
  or (_41898_, \oc8051_gm_cxrom_1.cell5.data [3], _41806_);
  and (_01691_, _41898_, _41897_);
  or (_41899_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41900_, \oc8051_gm_cxrom_1.cell5.data [4], _41874_);
  nand (_41901_, _41900_, _41899_);
  nand (_41902_, _41901_, _41806_);
  or (_41903_, \oc8051_gm_cxrom_1.cell5.data [4], _41806_);
  and (_01695_, _41903_, _41902_);
  or (_41904_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41905_, \oc8051_gm_cxrom_1.cell5.data [5], _41874_);
  nand (_41906_, _41905_, _41904_);
  nand (_41907_, _41906_, _41806_);
  or (_41908_, \oc8051_gm_cxrom_1.cell5.data [5], _41806_);
  and (_01699_, _41908_, _41907_);
  or (_41909_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_41910_, \oc8051_gm_cxrom_1.cell5.data [6], _41874_);
  nand (_41911_, _41910_, _41909_);
  nand (_41912_, _41911_, _41806_);
  or (_41913_, \oc8051_gm_cxrom_1.cell5.data [6], _41806_);
  and (_01703_, _41913_, _41912_);
  or (_41914_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_41915_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_41916_, _41915_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_41917_, _41916_, _41914_);
  nand (_41918_, _41917_, _41806_);
  or (_41919_, \oc8051_gm_cxrom_1.cell6.data [7], _41806_);
  and (_01725_, _41919_, _41918_);
  or (_41920_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41921_, \oc8051_gm_cxrom_1.cell6.data [0], _41915_);
  nand (_41922_, _41921_, _41920_);
  nand (_41923_, _41922_, _41806_);
  or (_41924_, \oc8051_gm_cxrom_1.cell6.data [0], _41806_);
  and (_01732_, _41924_, _41923_);
  or (_41925_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41926_, \oc8051_gm_cxrom_1.cell6.data [1], _41915_);
  nand (_41927_, _41926_, _41925_);
  nand (_41928_, _41927_, _41806_);
  or (_41929_, \oc8051_gm_cxrom_1.cell6.data [1], _41806_);
  and (_01736_, _41929_, _41928_);
  or (_41930_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41931_, \oc8051_gm_cxrom_1.cell6.data [2], _41915_);
  nand (_41932_, _41931_, _41930_);
  nand (_41933_, _41932_, _41806_);
  or (_41934_, \oc8051_gm_cxrom_1.cell6.data [2], _41806_);
  and (_01740_, _41934_, _41933_);
  or (_41935_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41936_, \oc8051_gm_cxrom_1.cell6.data [3], _41915_);
  nand (_41937_, _41936_, _41935_);
  nand (_41938_, _41937_, _41806_);
  or (_41939_, \oc8051_gm_cxrom_1.cell6.data [3], _41806_);
  and (_01743_, _41939_, _41938_);
  or (_41940_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41941_, \oc8051_gm_cxrom_1.cell6.data [4], _41915_);
  nand (_41942_, _41941_, _41940_);
  nand (_41943_, _41942_, _41806_);
  or (_41944_, \oc8051_gm_cxrom_1.cell6.data [4], _41806_);
  and (_01747_, _41944_, _41943_);
  or (_41945_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41946_, \oc8051_gm_cxrom_1.cell6.data [5], _41915_);
  nand (_41947_, _41946_, _41945_);
  nand (_41948_, _41947_, _41806_);
  or (_41949_, \oc8051_gm_cxrom_1.cell6.data [5], _41806_);
  and (_01751_, _41949_, _41948_);
  or (_41950_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_41951_, \oc8051_gm_cxrom_1.cell6.data [6], _41915_);
  nand (_41952_, _41951_, _41950_);
  nand (_41953_, _41952_, _41806_);
  or (_41954_, \oc8051_gm_cxrom_1.cell6.data [6], _41806_);
  and (_01755_, _41954_, _41953_);
  or (_41955_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_41956_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_41957_, _41956_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_41958_, _41957_, _41955_);
  nand (_41959_, _41958_, _41806_);
  or (_41960_, \oc8051_gm_cxrom_1.cell7.data [7], _41806_);
  and (_01777_, _41960_, _41959_);
  or (_41961_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41962_, \oc8051_gm_cxrom_1.cell7.data [0], _41956_);
  nand (_41963_, _41962_, _41961_);
  nand (_41964_, _41963_, _41806_);
  or (_41965_, \oc8051_gm_cxrom_1.cell7.data [0], _41806_);
  and (_01783_, _41965_, _41964_);
  or (_41966_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41967_, \oc8051_gm_cxrom_1.cell7.data [1], _41956_);
  nand (_41968_, _41967_, _41966_);
  nand (_41969_, _41968_, _41806_);
  or (_41970_, \oc8051_gm_cxrom_1.cell7.data [1], _41806_);
  and (_01787_, _41970_, _41969_);
  or (_41971_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41972_, \oc8051_gm_cxrom_1.cell7.data [2], _41956_);
  nand (_41973_, _41972_, _41971_);
  nand (_41974_, _41973_, _41806_);
  or (_41975_, \oc8051_gm_cxrom_1.cell7.data [2], _41806_);
  and (_01791_, _41975_, _41974_);
  or (_41976_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41977_, \oc8051_gm_cxrom_1.cell7.data [3], _41956_);
  nand (_41978_, _41977_, _41976_);
  nand (_41979_, _41978_, _41806_);
  or (_41980_, \oc8051_gm_cxrom_1.cell7.data [3], _41806_);
  and (_01795_, _41980_, _41979_);
  or (_41981_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41982_, \oc8051_gm_cxrom_1.cell7.data [4], _41956_);
  nand (_41983_, _41982_, _41981_);
  nand (_41984_, _41983_, _41806_);
  or (_41985_, \oc8051_gm_cxrom_1.cell7.data [4], _41806_);
  and (_01799_, _41985_, _41984_);
  or (_41986_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41987_, \oc8051_gm_cxrom_1.cell7.data [5], _41956_);
  nand (_41988_, _41987_, _41986_);
  nand (_41989_, _41988_, _41806_);
  or (_41990_, \oc8051_gm_cxrom_1.cell7.data [5], _41806_);
  and (_01803_, _41990_, _41989_);
  or (_41991_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_41992_, \oc8051_gm_cxrom_1.cell7.data [6], _41956_);
  nand (_41993_, _41992_, _41991_);
  nand (_41994_, _41993_, _41806_);
  or (_41995_, \oc8051_gm_cxrom_1.cell7.data [6], _41806_);
  and (_01807_, _41995_, _41994_);
  or (_41996_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_41997_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_41998_, _41997_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_41999_, _41998_, _41996_);
  nand (_42000_, _41999_, _41806_);
  or (_42001_, \oc8051_gm_cxrom_1.cell8.data [7], _41806_);
  and (_01828_, _42001_, _42000_);
  or (_42002_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42003_, \oc8051_gm_cxrom_1.cell8.data [0], _41997_);
  nand (_42004_, _42003_, _42002_);
  nand (_42005_, _42004_, _41806_);
  or (_42006_, \oc8051_gm_cxrom_1.cell8.data [0], _41806_);
  and (_01835_, _42006_, _42005_);
  or (_42007_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42008_, \oc8051_gm_cxrom_1.cell8.data [1], _41997_);
  nand (_42009_, _42008_, _42007_);
  nand (_42010_, _42009_, _41806_);
  or (_42011_, \oc8051_gm_cxrom_1.cell8.data [1], _41806_);
  and (_01839_, _42011_, _42010_);
  or (_42012_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42013_, \oc8051_gm_cxrom_1.cell8.data [2], _41997_);
  nand (_42014_, _42013_, _42012_);
  nand (_42015_, _42014_, _41806_);
  or (_42016_, \oc8051_gm_cxrom_1.cell8.data [2], _41806_);
  and (_01843_, _42016_, _42015_);
  or (_42017_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42018_, \oc8051_gm_cxrom_1.cell8.data [3], _41997_);
  nand (_42019_, _42018_, _42017_);
  nand (_42020_, _42019_, _41806_);
  or (_42021_, \oc8051_gm_cxrom_1.cell8.data [3], _41806_);
  and (_01847_, _42021_, _42020_);
  or (_42022_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42023_, \oc8051_gm_cxrom_1.cell8.data [4], _41997_);
  nand (_42024_, _42023_, _42022_);
  nand (_42025_, _42024_, _41806_);
  or (_42026_, \oc8051_gm_cxrom_1.cell8.data [4], _41806_);
  and (_01851_, _42026_, _42025_);
  or (_42027_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42028_, \oc8051_gm_cxrom_1.cell8.data [5], _41997_);
  nand (_42029_, _42028_, _42027_);
  nand (_42030_, _42029_, _41806_);
  or (_42031_, \oc8051_gm_cxrom_1.cell8.data [5], _41806_);
  and (_01854_, _42031_, _42030_);
  or (_42032_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42033_, \oc8051_gm_cxrom_1.cell8.data [6], _41997_);
  nand (_42034_, _42033_, _42032_);
  nand (_42035_, _42034_, _41806_);
  or (_42036_, \oc8051_gm_cxrom_1.cell8.data [6], _41806_);
  and (_01858_, _42036_, _42035_);
  or (_42037_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_42038_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_42039_, _42038_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_42040_, _42039_, _42037_);
  nand (_42041_, _42040_, _41806_);
  or (_42042_, \oc8051_gm_cxrom_1.cell9.data [7], _41806_);
  and (_01880_, _42042_, _42041_);
  or (_42043_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42044_, \oc8051_gm_cxrom_1.cell9.data [0], _42038_);
  nand (_42045_, _42044_, _42043_);
  nand (_42046_, _42045_, _41806_);
  or (_42047_, \oc8051_gm_cxrom_1.cell9.data [0], _41806_);
  and (_01887_, _42047_, _42046_);
  or (_42048_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42049_, \oc8051_gm_cxrom_1.cell9.data [1], _42038_);
  nand (_42050_, _42049_, _42048_);
  nand (_42051_, _42050_, _41806_);
  or (_42052_, \oc8051_gm_cxrom_1.cell9.data [1], _41806_);
  and (_01891_, _42052_, _42051_);
  or (_42053_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42054_, \oc8051_gm_cxrom_1.cell9.data [2], _42038_);
  nand (_42055_, _42054_, _42053_);
  nand (_42056_, _42055_, _41806_);
  or (_42057_, \oc8051_gm_cxrom_1.cell9.data [2], _41806_);
  and (_01895_, _42057_, _42056_);
  or (_42058_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42059_, \oc8051_gm_cxrom_1.cell9.data [3], _42038_);
  nand (_42060_, _42059_, _42058_);
  nand (_42061_, _42060_, _41806_);
  or (_42062_, \oc8051_gm_cxrom_1.cell9.data [3], _41806_);
  and (_01899_, _42062_, _42061_);
  or (_42063_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42064_, \oc8051_gm_cxrom_1.cell9.data [4], _42038_);
  nand (_42065_, _42064_, _42063_);
  nand (_42066_, _42065_, _41806_);
  or (_42067_, \oc8051_gm_cxrom_1.cell9.data [4], _41806_);
  and (_01903_, _42067_, _42066_);
  or (_42068_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42069_, \oc8051_gm_cxrom_1.cell9.data [5], _42038_);
  nand (_42070_, _42069_, _42068_);
  nand (_42071_, _42070_, _41806_);
  or (_42072_, \oc8051_gm_cxrom_1.cell9.data [5], _41806_);
  and (_01907_, _42072_, _42071_);
  or (_42073_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42074_, \oc8051_gm_cxrom_1.cell9.data [6], _42038_);
  nand (_42075_, _42074_, _42073_);
  nand (_42076_, _42075_, _41806_);
  or (_42077_, \oc8051_gm_cxrom_1.cell9.data [6], _41806_);
  and (_01910_, _42077_, _42076_);
  or (_42078_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_42079_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_42080_, _42079_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_42081_, _42080_, _42078_);
  nand (_42082_, _42081_, _41806_);
  or (_42083_, \oc8051_gm_cxrom_1.cell10.data [7], _41806_);
  and (_01932_, _42083_, _42082_);
  or (_42084_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42085_, \oc8051_gm_cxrom_1.cell10.data [0], _42079_);
  nand (_42086_, _42085_, _42084_);
  nand (_42087_, _42086_, _41806_);
  or (_42088_, \oc8051_gm_cxrom_1.cell10.data [0], _41806_);
  and (_01939_, _42088_, _42087_);
  or (_42089_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42090_, \oc8051_gm_cxrom_1.cell10.data [1], _42079_);
  nand (_42091_, _42090_, _42089_);
  nand (_42092_, _42091_, _41806_);
  or (_42093_, \oc8051_gm_cxrom_1.cell10.data [1], _41806_);
  and (_01943_, _42093_, _42092_);
  or (_42094_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42095_, \oc8051_gm_cxrom_1.cell10.data [2], _42079_);
  nand (_42096_, _42095_, _42094_);
  nand (_42097_, _42096_, _41806_);
  or (_42098_, \oc8051_gm_cxrom_1.cell10.data [2], _41806_);
  and (_01947_, _42098_, _42097_);
  or (_42099_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42100_, \oc8051_gm_cxrom_1.cell10.data [3], _42079_);
  nand (_42101_, _42100_, _42099_);
  nand (_42102_, _42101_, _41806_);
  or (_42103_, \oc8051_gm_cxrom_1.cell10.data [3], _41806_);
  and (_01951_, _42103_, _42102_);
  or (_42104_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42105_, \oc8051_gm_cxrom_1.cell10.data [4], _42079_);
  nand (_42106_, _42105_, _42104_);
  nand (_42107_, _42106_, _41806_);
  or (_42108_, \oc8051_gm_cxrom_1.cell10.data [4], _41806_);
  and (_01955_, _42108_, _42107_);
  or (_42109_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42110_, \oc8051_gm_cxrom_1.cell10.data [5], _42079_);
  nand (_42111_, _42110_, _42109_);
  nand (_42112_, _42111_, _41806_);
  or (_42113_, \oc8051_gm_cxrom_1.cell10.data [5], _41806_);
  and (_01959_, _42113_, _42112_);
  or (_42114_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42115_, \oc8051_gm_cxrom_1.cell10.data [6], _42079_);
  nand (_42116_, _42115_, _42114_);
  nand (_42117_, _42116_, _41806_);
  or (_42118_, \oc8051_gm_cxrom_1.cell10.data [6], _41806_);
  and (_01963_, _42118_, _42117_);
  or (_42119_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_42120_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_42121_, _42120_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_42122_, _42121_, _42119_);
  nand (_42123_, _42122_, _41806_);
  or (_42124_, \oc8051_gm_cxrom_1.cell11.data [7], _41806_);
  and (_01984_, _42124_, _42123_);
  or (_42125_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42126_, \oc8051_gm_cxrom_1.cell11.data [0], _42120_);
  nand (_42127_, _42126_, _42125_);
  nand (_42128_, _42127_, _41806_);
  or (_42129_, \oc8051_gm_cxrom_1.cell11.data [0], _41806_);
  and (_01991_, _42129_, _42128_);
  or (_42130_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42131_, \oc8051_gm_cxrom_1.cell11.data [1], _42120_);
  nand (_42132_, _42131_, _42130_);
  nand (_42133_, _42132_, _41806_);
  or (_42134_, \oc8051_gm_cxrom_1.cell11.data [1], _41806_);
  and (_01995_, _42134_, _42133_);
  or (_42135_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42136_, \oc8051_gm_cxrom_1.cell11.data [2], _42120_);
  nand (_42137_, _42136_, _42135_);
  nand (_42138_, _42137_, _41806_);
  or (_42139_, \oc8051_gm_cxrom_1.cell11.data [2], _41806_);
  and (_01999_, _42139_, _42138_);
  or (_42140_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42141_, \oc8051_gm_cxrom_1.cell11.data [3], _42120_);
  nand (_42142_, _42141_, _42140_);
  nand (_42143_, _42142_, _41806_);
  or (_42144_, \oc8051_gm_cxrom_1.cell11.data [3], _41806_);
  and (_02003_, _42144_, _42143_);
  or (_42145_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42146_, \oc8051_gm_cxrom_1.cell11.data [4], _42120_);
  nand (_42147_, _42146_, _42145_);
  nand (_42148_, _42147_, _41806_);
  or (_42149_, \oc8051_gm_cxrom_1.cell11.data [4], _41806_);
  and (_02007_, _42149_, _42148_);
  or (_42150_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42151_, \oc8051_gm_cxrom_1.cell11.data [5], _42120_);
  nand (_42152_, _42151_, _42150_);
  nand (_42153_, _42152_, _41806_);
  or (_42154_, \oc8051_gm_cxrom_1.cell11.data [5], _41806_);
  and (_02011_, _42154_, _42153_);
  or (_42155_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42156_, \oc8051_gm_cxrom_1.cell11.data [6], _42120_);
  nand (_42157_, _42156_, _42155_);
  nand (_42158_, _42157_, _41806_);
  or (_42159_, \oc8051_gm_cxrom_1.cell11.data [6], _41806_);
  and (_02015_, _42159_, _42158_);
  or (_42160_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_42161_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_42162_, _42161_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_42163_, _42162_, _42160_);
  nand (_42164_, _42163_, _41806_);
  or (_42165_, \oc8051_gm_cxrom_1.cell12.data [7], _41806_);
  and (_02036_, _42165_, _42164_);
  or (_42166_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42167_, \oc8051_gm_cxrom_1.cell12.data [0], _42161_);
  nand (_42168_, _42167_, _42166_);
  nand (_42169_, _42168_, _41806_);
  or (_42170_, \oc8051_gm_cxrom_1.cell12.data [0], _41806_);
  and (_02043_, _42170_, _42169_);
  or (_42171_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42172_, \oc8051_gm_cxrom_1.cell12.data [1], _42161_);
  nand (_42173_, _42172_, _42171_);
  nand (_42174_, _42173_, _41806_);
  or (_42175_, \oc8051_gm_cxrom_1.cell12.data [1], _41806_);
  and (_02047_, _42175_, _42174_);
  or (_42176_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42177_, \oc8051_gm_cxrom_1.cell12.data [2], _42161_);
  nand (_42178_, _42177_, _42176_);
  nand (_42179_, _42178_, _41806_);
  or (_42180_, \oc8051_gm_cxrom_1.cell12.data [2], _41806_);
  and (_02051_, _42180_, _42179_);
  or (_42181_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42182_, \oc8051_gm_cxrom_1.cell12.data [3], _42161_);
  nand (_42183_, _42182_, _42181_);
  nand (_42184_, _42183_, _41806_);
  or (_42185_, \oc8051_gm_cxrom_1.cell12.data [3], _41806_);
  and (_02055_, _42185_, _42184_);
  or (_42186_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42187_, \oc8051_gm_cxrom_1.cell12.data [4], _42161_);
  nand (_42188_, _42187_, _42186_);
  nand (_42189_, _42188_, _41806_);
  or (_42190_, \oc8051_gm_cxrom_1.cell12.data [4], _41806_);
  and (_02059_, _42190_, _42189_);
  or (_42191_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42192_, \oc8051_gm_cxrom_1.cell12.data [5], _42161_);
  nand (_42193_, _42192_, _42191_);
  nand (_42194_, _42193_, _41806_);
  or (_42195_, \oc8051_gm_cxrom_1.cell12.data [5], _41806_);
  and (_02063_, _42195_, _42194_);
  or (_42196_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42197_, \oc8051_gm_cxrom_1.cell12.data [6], _42161_);
  nand (_42198_, _42197_, _42196_);
  nand (_42199_, _42198_, _41806_);
  or (_42200_, \oc8051_gm_cxrom_1.cell12.data [6], _41806_);
  and (_02067_, _42200_, _42199_);
  or (_42201_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_42202_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_42203_, _42202_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_42204_, _42203_, _42201_);
  nand (_42205_, _42204_, _41806_);
  or (_42206_, \oc8051_gm_cxrom_1.cell13.data [7], _41806_);
  and (_02088_, _42206_, _42205_);
  or (_42207_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42208_, \oc8051_gm_cxrom_1.cell13.data [0], _42202_);
  nand (_42209_, _42208_, _42207_);
  nand (_42210_, _42209_, _41806_);
  or (_42211_, \oc8051_gm_cxrom_1.cell13.data [0], _41806_);
  and (_02095_, _42211_, _42210_);
  or (_42212_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42213_, \oc8051_gm_cxrom_1.cell13.data [1], _42202_);
  nand (_42214_, _42213_, _42212_);
  nand (_42215_, _42214_, _41806_);
  or (_42216_, \oc8051_gm_cxrom_1.cell13.data [1], _41806_);
  and (_02099_, _42216_, _42215_);
  or (_42217_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42218_, \oc8051_gm_cxrom_1.cell13.data [2], _42202_);
  nand (_42219_, _42218_, _42217_);
  nand (_42220_, _42219_, _41806_);
  or (_42221_, \oc8051_gm_cxrom_1.cell13.data [2], _41806_);
  and (_02103_, _42221_, _42220_);
  or (_42222_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42223_, \oc8051_gm_cxrom_1.cell13.data [3], _42202_);
  nand (_42224_, _42223_, _42222_);
  nand (_42225_, _42224_, _41806_);
  or (_42226_, \oc8051_gm_cxrom_1.cell13.data [3], _41806_);
  and (_02107_, _42226_, _42225_);
  or (_42227_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42228_, \oc8051_gm_cxrom_1.cell13.data [4], _42202_);
  nand (_42229_, _42228_, _42227_);
  nand (_42230_, _42229_, _41806_);
  or (_42231_, \oc8051_gm_cxrom_1.cell13.data [4], _41806_);
  and (_02111_, _42231_, _42230_);
  or (_42232_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42233_, \oc8051_gm_cxrom_1.cell13.data [5], _42202_);
  nand (_42234_, _42233_, _42232_);
  nand (_42235_, _42234_, _41806_);
  or (_42236_, \oc8051_gm_cxrom_1.cell13.data [5], _41806_);
  and (_02115_, _42236_, _42235_);
  or (_42237_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42238_, \oc8051_gm_cxrom_1.cell13.data [6], _42202_);
  nand (_42239_, _42238_, _42237_);
  nand (_42240_, _42239_, _41806_);
  or (_42241_, \oc8051_gm_cxrom_1.cell13.data [6], _41806_);
  and (_02119_, _42241_, _42240_);
  or (_42242_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_42243_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_42244_, _42243_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_42245_, _42244_, _42242_);
  nand (_42246_, _42245_, _41806_);
  or (_42247_, \oc8051_gm_cxrom_1.cell14.data [7], _41806_);
  and (_02140_, _42247_, _42246_);
  or (_42248_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42249_, \oc8051_gm_cxrom_1.cell14.data [0], _42243_);
  nand (_42250_, _42249_, _42248_);
  nand (_42251_, _42250_, _41806_);
  or (_42252_, \oc8051_gm_cxrom_1.cell14.data [0], _41806_);
  and (_02147_, _42252_, _42251_);
  or (_42253_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42254_, \oc8051_gm_cxrom_1.cell14.data [1], _42243_);
  nand (_42255_, _42254_, _42253_);
  nand (_42256_, _42255_, _41806_);
  or (_42257_, \oc8051_gm_cxrom_1.cell14.data [1], _41806_);
  and (_02151_, _42257_, _42256_);
  or (_42258_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42259_, \oc8051_gm_cxrom_1.cell14.data [2], _42243_);
  nand (_42260_, _42259_, _42258_);
  nand (_42261_, _42260_, _41806_);
  or (_42262_, \oc8051_gm_cxrom_1.cell14.data [2], _41806_);
  and (_02155_, _42262_, _42261_);
  or (_42263_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42264_, \oc8051_gm_cxrom_1.cell14.data [3], _42243_);
  nand (_42265_, _42264_, _42263_);
  nand (_42266_, _42265_, _41806_);
  or (_42267_, \oc8051_gm_cxrom_1.cell14.data [3], _41806_);
  and (_02159_, _42267_, _42266_);
  or (_42268_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42269_, \oc8051_gm_cxrom_1.cell14.data [4], _42243_);
  nand (_42270_, _42269_, _42268_);
  nand (_42271_, _42270_, _41806_);
  or (_42272_, \oc8051_gm_cxrom_1.cell14.data [4], _41806_);
  and (_02163_, _42272_, _42271_);
  or (_42273_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42274_, \oc8051_gm_cxrom_1.cell14.data [5], _42243_);
  nand (_42275_, _42274_, _42273_);
  nand (_42276_, _42275_, _41806_);
  or (_42277_, \oc8051_gm_cxrom_1.cell14.data [5], _41806_);
  and (_02167_, _42277_, _42276_);
  or (_42278_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42279_, \oc8051_gm_cxrom_1.cell14.data [6], _42243_);
  nand (_42280_, _42279_, _42278_);
  nand (_42281_, _42280_, _41806_);
  or (_42282_, \oc8051_gm_cxrom_1.cell14.data [6], _41806_);
  and (_02171_, _42282_, _42281_);
  or (_42283_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_42284_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_42285_, _42284_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_42286_, _42285_, _42283_);
  nand (_42287_, _42286_, _41806_);
  or (_42288_, \oc8051_gm_cxrom_1.cell15.data [7], _41806_);
  and (_02192_, _42288_, _42287_);
  or (_42289_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42290_, \oc8051_gm_cxrom_1.cell15.data [0], _42284_);
  nand (_42291_, _42290_, _42289_);
  nand (_42292_, _42291_, _41806_);
  or (_42293_, \oc8051_gm_cxrom_1.cell15.data [0], _41806_);
  and (_02199_, _42293_, _42292_);
  or (_42294_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42295_, \oc8051_gm_cxrom_1.cell15.data [1], _42284_);
  nand (_42296_, _42295_, _42294_);
  nand (_42297_, _42296_, _41806_);
  or (_42298_, \oc8051_gm_cxrom_1.cell15.data [1], _41806_);
  and (_02203_, _42298_, _42297_);
  or (_42299_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42300_, \oc8051_gm_cxrom_1.cell15.data [2], _42284_);
  nand (_42301_, _42300_, _42299_);
  nand (_42302_, _42301_, _41806_);
  or (_42303_, \oc8051_gm_cxrom_1.cell15.data [2], _41806_);
  and (_02207_, _42303_, _42302_);
  or (_42304_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42305_, \oc8051_gm_cxrom_1.cell15.data [3], _42284_);
  nand (_42306_, _42305_, _42304_);
  nand (_42307_, _42306_, _41806_);
  or (_42308_, \oc8051_gm_cxrom_1.cell15.data [3], _41806_);
  and (_02211_, _42308_, _42307_);
  or (_42309_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42310_, \oc8051_gm_cxrom_1.cell15.data [4], _42284_);
  nand (_42311_, _42310_, _42309_);
  nand (_42312_, _42311_, _41806_);
  or (_42313_, \oc8051_gm_cxrom_1.cell15.data [4], _41806_);
  and (_02215_, _42313_, _42312_);
  or (_42314_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42315_, \oc8051_gm_cxrom_1.cell15.data [5], _42284_);
  nand (_42316_, _42315_, _42314_);
  nand (_42317_, _42316_, _41806_);
  or (_42318_, \oc8051_gm_cxrom_1.cell15.data [5], _41806_);
  and (_02219_, _42318_, _42317_);
  or (_42319_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42320_, \oc8051_gm_cxrom_1.cell15.data [6], _42284_);
  nand (_42321_, _42320_, _42319_);
  nand (_42322_, _42321_, _41806_);
  or (_42323_, \oc8051_gm_cxrom_1.cell15.data [6], _41806_);
  and (_02223_, _42323_, _42322_);
  nor (_05996_, _37932_, rst);
  and (_42324_, _33860_, _41806_);
  nand (_42325_, _42324_, _36091_);
  nor (_42326_, _36584_, _36453_);
  or (_05999_, _42326_, _42325_);
  and (_42327_, _35242_, _35012_);
  and (_42328_, _42327_, _35496_);
  not (_42329_, _34486_);
  nor (_42330_, _34727_, _34233_);
  and (_42331_, _42330_, _42329_);
  and (_42332_, _42331_, _42328_);
  not (_42333_, _34233_);
  and (_42334_, _34727_, _42333_);
  not (_42335_, _35751_);
  not (_42336_, _35242_);
  and (_42337_, _35496_, _42336_);
  not (_42338_, _35012_);
  and (_42339_, _36365_, _42338_);
  and (_42340_, _42339_, _42337_);
  and (_42341_, _42340_, _42335_);
  and (_42342_, _42341_, _42334_);
  and (_42343_, _42335_, _34486_);
  nor (_42344_, _42335_, _34486_);
  nor (_42345_, _42344_, _42343_);
  and (_42346_, _35496_, _35242_);
  and (_42347_, _42346_, _42339_);
  and (_42348_, _34727_, _34233_);
  and (_42349_, _42348_, _42347_);
  and (_42350_, _42349_, _42345_);
  or (_42351_, _42350_, _42342_);
  or (_42352_, _42351_, _42332_);
  not (_42353_, _34727_);
  and (_42354_, _42353_, _34233_);
  and (_42355_, _42354_, _42344_);
  not (_42356_, _36365_);
  and (_42357_, _42328_, _42356_);
  and (_42358_, _42357_, _42355_);
  and (_42359_, _42344_, _42334_);
  not (_42360_, _35496_);
  and (_42361_, _42336_, _35012_);
  nor (_42362_, _42361_, _42360_);
  not (_42363_, _42362_);
  and (_42364_, _42363_, _42359_);
  or (_42365_, _42364_, _42358_);
  and (_42366_, _35751_, _34486_);
  and (_42367_, _42366_, _42330_);
  and (_42368_, _42337_, _42338_);
  and (_42369_, _42368_, _42356_);
  and (_42370_, _42369_, _42367_);
  and (_42371_, _42348_, _42329_);
  and (_42372_, _42328_, _36365_);
  and (_42373_, _42372_, _42371_);
  or (_42374_, _42373_, _42370_);
  or (_42375_, _42374_, _42365_);
  and (_42376_, _42343_, _42334_);
  and (_42377_, _42347_, _42376_);
  and (_42378_, _42367_, _42360_);
  nor (_42379_, _42378_, _42377_);
  and (_42380_, _42354_, _35751_);
  and (_42381_, _42380_, _42347_);
  and (_42382_, _42348_, _34486_);
  and (_42383_, _42382_, _42372_);
  nor (_42384_, _42383_, _42381_);
  nand (_42385_, _42384_, _42379_);
  or (_42386_, _42385_, _42375_);
  nor (_42387_, _35751_, _34486_);
  and (_42388_, _42354_, _42387_);
  nor (_42389_, _42388_, _42356_);
  and (_42390_, _42346_, _42338_);
  not (_42391_, _42390_);
  nor (_42392_, _42391_, _42389_);
  not (_42393_, _42392_);
  and (_42394_, _42348_, _42344_);
  and (_42395_, _42394_, _42347_);
  and (_42396_, _42354_, _42343_);
  and (_42397_, _42396_, _42347_);
  nor (_42398_, _42397_, _42395_);
  and (_42399_, _42398_, _42393_);
  and (_42400_, _42359_, _42368_);
  and (_42401_, _42334_, _34486_);
  and (_42402_, _42357_, _42401_);
  and (_42403_, _42347_, _42331_);
  or (_42404_, _42403_, _42402_);
  nor (_42405_, _42404_, _42400_);
  nand (_42406_, _42405_, _42399_);
  or (_42407_, _42406_, _42386_);
  or (_42408_, _42407_, _42352_);
  and (_42409_, _42408_, _33881_);
  not (_42410_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_42411_, _33849_, _15636_);
  and (_42412_, _42411_, _36727_);
  nor (_42413_, _42412_, _42410_);
  or (_42414_, _42413_, rst);
  or (_06002_, _42414_, _42409_);
  nand (_42415_, _34233_, _33806_);
  or (_42416_, _33806_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_42417_, _42416_, _41806_);
  and (_06005_, _42417_, _42415_);
  and (_42418_, \oc8051_top_1.oc8051_sfr1.wait_data , _41806_);
  and (_42419_, _42418_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_42420_, _36464_, _36124_);
  and (_42421_, _37833_, _36935_);
  or (_42422_, _42421_, _42420_);
  and (_42423_, _36584_, _36124_);
  or (_42424_, _42423_, _37657_);
  or (_42425_, _42424_, _37340_);
  and (_42426_, _37102_, _36464_);
  and (_42427_, _36595_, _36453_);
  or (_42428_, _42427_, _42426_);
  or (_42429_, _42428_, _42425_);
  or (_42430_, _42429_, _37550_);
  or (_42431_, _42430_, _42422_);
  and (_42432_, _42431_, _42324_);
  or (_06008_, _42432_, _42419_);
  and (_42433_, _36584_, _36003_);
  or (_42434_, _42433_, _36485_);
  and (_42435_, _37023_, _36025_);
  or (_42436_, _42435_, _36036_);
  and (_42437_, _36880_, _35056_);
  and (_42438_, _42437_, _37102_);
  or (_42439_, _42438_, _42436_);
  or (_42440_, _42439_, _42434_);
  and (_42441_, _42440_, _33860_);
  and (_42442_, \oc8051_top_1.oc8051_decoder1.state [0], _15636_);
  and (_42443_, _42442_, _42410_);
  not (_42444_, _37866_);
  and (_42445_, _42444_, _42443_);
  and (_42446_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42447_, _42446_, _42445_);
  or (_42448_, _42447_, _42441_);
  and (_06011_, _42448_, _41806_);
  and (_42449_, _42418_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_42450_, _37833_, _37045_);
  not (_42451_, _36902_);
  nor (_42452_, _37045_, _36595_);
  nor (_42453_, _42452_, _42451_);
  or (_42454_, _42453_, _42450_);
  and (_42455_, _42437_, _37186_);
  or (_42456_, _42455_, _42454_);
  nor (_42457_, _42452_, _35542_);
  not (_42458_, _35542_);
  and (_42459_, _37186_, _42458_);
  or (_42460_, _42459_, _42457_);
  nor (_42461_, _35795_, _35542_);
  and (_42462_, _42461_, _35959_);
  and (_42463_, _37833_, _36913_);
  nor (_42464_, _42463_, _42462_);
  nand (_42465_, _42464_, _35981_);
  or (_42466_, _42465_, _42434_);
  or (_42467_, _42466_, _42460_);
  or (_42468_, _42467_, _42456_);
  and (_42469_, _42468_, _42324_);
  or (_06014_, _42469_, _42449_);
  and (_42470_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42471_, _37394_, _33860_);
  or (_42472_, _42471_, _42470_);
  or (_42473_, _42472_, _42445_);
  and (_06017_, _42473_, _41806_);
  and (_42474_, _36464_, _35992_);
  not (_42475_, _36935_);
  nor (_42476_, _42326_, _42475_);
  nor (_42477_, _42476_, _42474_);
  not (_42478_, _42477_);
  and (_42479_, _42478_, _42443_);
  and (_42480_, _37186_, _36628_);
  and (_42481_, _36891_, _36442_);
  and (_42482_, _42481_, _35806_);
  or (_42483_, _42482_, _42480_);
  or (_42484_, _42483_, _42420_);
  and (_42485_, _42484_, _36858_);
  or (_42486_, _42485_, _42479_);
  and (_42487_, _42483_, _36749_);
  or (_42488_, _42487_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42489_, _42488_, _42486_);
  or (_42490_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _15636_);
  and (_42491_, _42490_, _41806_);
  and (_06020_, _42491_, _42489_);
  and (_42492_, _42418_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_42493_, _42459_, _36485_);
  and (_42494_, _36595_, _42458_);
  or (_42495_, _42494_, _37263_);
  or (_42496_, _42495_, _42493_);
  and (_42497_, _36628_, _35959_);
  or (_42498_, _42455_, _42427_);
  or (_42499_, _42498_, _42497_);
  or (_42500_, _37186_, _37102_);
  and (_42501_, _42500_, _35850_);
  or (_42502_, _42435_, _37110_);
  or (_42503_, _42502_, _42501_);
  or (_42504_, _42503_, _42499_);
  or (_42505_, _42504_, _42496_);
  and (_42506_, _42505_, _42324_);
  or (_06023_, _42506_, _42492_);
  and (_42507_, _42418_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_42508_, _42438_, _37219_);
  and (_42509_, _36464_, _35860_);
  and (_42510_, _42437_, _36650_);
  or (_42511_, _42510_, _42509_);
  or (_42512_, _42511_, _42508_);
  or (_42513_, _42512_, _42460_);
  and (_42514_, _37833_, _37164_);
  or (_42515_, _37252_, _37175_);
  or (_42516_, _42515_, _42514_);
  and (_42517_, _36069_, _34782_);
  or (_42518_, _42517_, _36661_);
  and (_42519_, _36595_, _35850_);
  or (_42520_, _42519_, _42518_);
  or (_42521_, _42520_, _42516_);
  or (_42522_, _42521_, _42513_);
  and (_42523_, _37023_, _34782_);
  and (_42524_, _37023_, _36507_);
  or (_42525_, _42524_, _42523_);
  nor (_42526_, _37421_, _35926_);
  nand (_42527_, _42526_, _37318_);
  or (_42528_, _42527_, _42525_);
  or (_42529_, _42528_, _42456_);
  or (_42530_, _42529_, _42522_);
  and (_42531_, _42530_, _42324_);
  or (_06026_, _42531_, _42507_);
  and (_42532_, _42461_, _35992_);
  or (_42533_, _42532_, _35882_);
  and (_42534_, _42437_, _35871_);
  and (_42535_, _35871_, _42458_);
  or (_42536_, _42535_, _36014_);
  or (_42537_, _42536_, _42534_);
  or (_42538_, _42537_, _42533_);
  and (_42539_, _42437_, _36003_);
  or (_42540_, _42539_, _42538_);
  and (_42541_, _42540_, _33860_);
  and (_42542_, _37855_, _15636_);
  and (_42543_, _37844_, _15636_);
  or (_42544_, _42543_, _42542_);
  and (_42545_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_42546_, _42545_, _42544_);
  or (_42547_, _42546_, _42541_);
  and (_06029_, _42547_, _41806_);
  or (_42548_, _37133_, _37110_);
  not (_42549_, _37351_);
  or (_42550_, _42453_, _42549_);
  or (_42551_, _42550_, _42548_);
  and (_42552_, _36080_, _35806_);
  and (_42553_, _42552_, _36902_);
  or (_42554_, _42553_, _37197_);
  or (_42555_, _42554_, _37175_);
  or (_42556_, _42555_, _42480_);
  or (_42557_, _42556_, _37443_);
  or (_42558_, _42557_, _42551_);
  or (_42559_, _37034_, _36135_);
  or (_42560_, _42559_, _37464_);
  or (_42561_, _42560_, _42436_);
  and (_42562_, _42552_, _35850_);
  or (_42563_, _42562_, _35926_);
  or (_42564_, _42563_, _36957_);
  and (_42565_, _36124_, _42458_);
  and (_42566_, _42461_, _36080_);
  or (_42567_, _42566_, _42482_);
  or (_42568_, _42567_, _42565_);
  or (_42569_, _42568_, _42564_);
  or (_42570_, _42569_, _42561_);
  or (_42571_, _42570_, _42460_);
  or (_42572_, _42571_, _42558_);
  and (_42573_, _42572_, _33860_);
  and (_42574_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42575_, _42487_, _42445_);
  and (_42576_, _37712_, _36749_);
  or (_42577_, _42576_, _42575_);
  or (_42578_, _42577_, _42574_);
  or (_42579_, _42578_, _42573_);
  and (_06032_, _42579_, _41806_);
  nor (_06091_, _36814_, rst);
  nor (_06093_, _37778_, rst);
  nand (_06096_, _42478_, _42324_);
  and (_42580_, _36584_, _36091_);
  or (_42581_, _42580_, _42474_);
  nand (_06099_, _42581_, _42324_);
  or (_42582_, _42373_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_42583_, _42582_, _42402_);
  or (_42584_, _42583_, _42342_);
  and (_42585_, _42584_, _42412_);
  nor (_42586_, _42411_, _36727_);
  or (_42587_, _42586_, rst);
  or (_06102_, _42587_, _42585_);
  nand (_42588_, _36365_, _33806_);
  or (_42589_, _33806_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_42590_, _42589_, _41806_);
  and (_06105_, _42590_, _42588_);
  not (_42591_, _33806_);
  or (_42592_, _35012_, _42591_);
  or (_42593_, _33806_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_42594_, _42593_, _41806_);
  and (_06108_, _42594_, _42592_);
  nand (_42595_, _35242_, _33806_);
  or (_42596_, _33806_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_42597_, _42596_, _41806_);
  and (_06111_, _42597_, _42595_);
  nand (_42598_, _35496_, _33806_);
  or (_42599_, _33806_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_42600_, _42599_, _41806_);
  and (_06114_, _42600_, _42598_);
  or (_42601_, _35751_, _42591_);
  or (_42602_, _33806_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_42603_, _42602_, _41806_);
  and (_06117_, _42603_, _42601_);
  nand (_42604_, _34486_, _33806_);
  or (_42605_, _33806_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_42606_, _42605_, _41806_);
  and (_06120_, _42606_, _42604_);
  nand (_42607_, _34727_, _33806_);
  or (_42608_, _33806_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_42609_, _42608_, _41806_);
  and (_06123_, _42609_, _42607_);
  and (_42610_, _37023_, _34793_);
  or (_42611_, _42534_, _36014_);
  or (_42612_, _42611_, _42610_);
  or (_42613_, _36485_, _36113_);
  or (_42614_, _42613_, _42612_);
  and (_42615_, _42437_, _37164_);
  or (_42616_, _42615_, _42433_);
  or (_42617_, _36595_, _35915_);
  and (_42618_, _42617_, _37833_);
  or (_42619_, _42618_, _42616_);
  or (_42620_, _42619_, _42614_);
  or (_42621_, _42524_, _42509_);
  and (_42622_, _42437_, _36990_);
  or (_42623_, _42622_, _42533_);
  or (_42624_, _42623_, _42621_);
  or (_42625_, _36946_, _36661_);
  or (_42626_, _42510_, _42421_);
  or (_42627_, _42626_, _42625_);
  or (_42628_, _42627_, _42624_);
  and (_42629_, _37001_, _42458_);
  or (_42630_, _42629_, _42539_);
  and (_42631_, _36091_, _35806_);
  and (_42632_, _42631_, _37833_);
  or (_42633_, _42632_, _35839_);
  and (_42634_, _37833_, _36518_);
  and (_42635_, _37023_, _36091_);
  or (_42636_, _42635_, _42634_);
  or (_42637_, _42636_, _42633_);
  or (_42638_, _42637_, _42630_);
  or (_42639_, _42638_, _42628_);
  or (_42640_, _42639_, _42620_);
  and (_42641_, _42640_, _33860_);
  and (_42642_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42643_, _42642_, _42479_);
  or (_42644_, _42643_, _42641_);
  and (_30468_, _42644_, _41806_);
  and (_42645_, _42418_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_42646_, _37164_, _36650_);
  and (_42647_, _42646_, _36628_);
  or (_42648_, _42616_, _42525_);
  or (_42649_, _42648_, _42647_);
  nor (_42650_, _42462_, _35970_);
  not (_42651_, _42650_);
  or (_42652_, _42651_, _42463_);
  or (_42653_, _42652_, _37118_);
  or (_42654_, _42653_, _42422_);
  or (_42655_, _36650_, _37001_);
  and (_42656_, _42655_, _37833_);
  or (_42657_, _42656_, _42520_);
  or (_42658_, _42657_, _42654_);
  or (_42659_, _42658_, _42649_);
  and (_42660_, _42659_, _42324_);
  or (_30471_, _42660_, _42645_);
  or (_42661_, _42482_, _36135_);
  or (_42662_, _42661_, _42565_);
  or (_42663_, _42662_, _37464_);
  or (_42664_, _42663_, _42558_);
  and (_42665_, _42664_, _33860_);
  and (_42666_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42667_, _42666_, _42577_);
  or (_42668_, _42667_, _42665_);
  and (_30473_, _42668_, _41806_);
  and (_42669_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42670_, _37416_, _35795_);
  or (_42671_, _42670_, _36036_);
  or (_42672_, _42671_, _42564_);
  or (_42673_, _42672_, _42483_);
  and (_42674_, _42673_, _33860_);
  or (_42675_, _42674_, _42669_);
  or (_42676_, _42675_, _42575_);
  and (_30475_, _42676_, _41806_);
  and (_42677_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42678_, _42479_, _37910_);
  or (_42679_, _42678_, _42677_);
  and (_42680_, _42679_, _41806_);
  or (_42681_, _42474_, _37855_);
  and (_42682_, _42534_, _35806_);
  or (_42683_, _42682_, _42622_);
  or (_42684_, _42683_, _42681_);
  or (_42685_, _42684_, _42483_);
  or (_42686_, _42533_, _35839_);
  or (_42687_, _42646_, _36518_);
  and (_42688_, _42687_, _37833_);
  or (_42689_, _42688_, _42686_);
  or (_42690_, _42689_, _42685_);
  and (_42691_, _37833_, _37102_);
  or (_42692_, _42509_, _42691_);
  or (_42693_, _42692_, _42630_);
  and (_42694_, _42437_, _37208_);
  or (_42695_, _42694_, _42421_);
  or (_42696_, _42632_, _37844_);
  or (_42697_, _42696_, _42618_);
  or (_42698_, _42697_, _42695_);
  and (_42699_, _42631_, _36902_);
  or (_42700_, _42562_, _36014_);
  or (_42701_, _42700_, _42566_);
  or (_42702_, _42701_, _42699_);
  and (_42703_, _42534_, _35795_);
  or (_42704_, _42703_, _36529_);
  and (_42705_, _37464_, _36409_);
  or (_42706_, _42705_, _42704_);
  or (_42707_, _42706_, _42702_);
  or (_42708_, _42707_, _42698_);
  or (_42709_, _42708_, _42693_);
  or (_42710_, _42709_, _42690_);
  and (_42711_, _42710_, _42324_);
  or (_30477_, _42711_, _42680_);
  or (_42712_, _37855_, _36014_);
  or (_42713_, _42553_, _42433_);
  or (_42714_, _42713_, _42712_);
  or (_42715_, _35297_, _42458_);
  and (_42716_, _42715_, _42631_);
  or (_42717_, _42716_, _37464_);
  or (_42718_, _42717_, _42714_);
  or (_42719_, _37012_, _36551_);
  or (_42720_, _42719_, _42718_);
  or (_42721_, _37421_, _37175_);
  and (_42722_, _42721_, _36420_);
  or (_42723_, _42722_, _42686_);
  or (_42724_, _42723_, _42720_);
  or (_42725_, _42698_, _42693_);
  or (_42726_, _42725_, _42724_);
  and (_42727_, _42726_, _33860_);
  and (_42728_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42730_, _42728_, _42678_);
  or (_42732_, _42730_, _42727_);
  and (_30479_, _42732_, _41806_);
  and (_42735_, _42418_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_42737_, _40330_);
  or (_42739_, _42539_, _42737_);
  and (_42741_, _36464_, _35915_);
  and (_42743_, _42741_, _35806_);
  and (_42745_, _42427_, _36420_);
  or (_42747_, _42745_, _42743_);
  or (_42749_, _42747_, _42496_);
  or (_42751_, _42749_, _42739_);
  not (_42753_, _40329_);
  or (_42755_, _42501_, _42753_);
  and (_42757_, _37833_, _36595_);
  or (_42759_, _42757_, _42455_);
  or (_42761_, _42759_, _42548_);
  or (_42763_, _42761_, _42755_);
  and (_42765_, _36464_, _37208_);
  or (_42767_, _42532_, _42435_);
  and (_42769_, _35882_, _35806_);
  or (_42771_, _42769_, _42767_);
  or (_42773_, _42771_, _42765_);
  and (_42775_, _37507_, _42458_);
  or (_42777_, _42775_, _36014_);
  or (_42779_, _42777_, _37384_);
  and (_42781_, _37507_, _36464_);
  or (_42783_, _42682_, _42781_);
  or (_42785_, _42783_, _42779_);
  or (_42787_, _42785_, _42773_);
  or (_42789_, _42787_, _42763_);
  or (_42790_, _42789_, _42751_);
  and (_42791_, _42790_, _42324_);
  or (_30481_, _42791_, _42735_);
  or (_42792_, _42438_, _37307_);
  or (_42793_, _42519_, _42517_);
  or (_42794_, _42793_, _42792_);
  or (_42795_, _42794_, _42516_);
  or (_42796_, _42795_, _42684_);
  or (_42797_, _42757_, _42781_);
  or (_42798_, _42743_, _42704_);
  or (_42799_, _42798_, _42797_);
  or (_42800_, _42523_, _36485_);
  or (_42801_, _42800_, _35893_);
  or (_42802_, _42629_, _37475_);
  or (_42803_, _42802_, _42801_);
  or (_42804_, _42803_, _42799_);
  or (_42805_, _42804_, _42796_);
  and (_42806_, _42805_, _42324_);
  and (_42807_, _33817_, _41806_);
  and (_42808_, _42807_, _37855_);
  and (_42809_, _42418_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_42810_, _42809_, _42808_);
  or (_30483_, _42810_, _42806_);
  and (_42811_, _36464_, _35871_);
  or (_42812_, _42767_, _42438_);
  or (_42813_, _42812_, _42811_);
  or (_42814_, _42462_, _37296_);
  nor (_42815_, _42814_, _42539_);
  nand (_42816_, _42815_, _36058_);
  or (_42817_, _42816_, _42813_);
  not (_42818_, _37454_);
  nor (_42819_, _42622_, _37464_);
  and (_42820_, _42819_, _42818_);
  not (_42821_, _42820_);
  or (_42822_, _42821_, _42460_);
  or (_42823_, _42822_, _42817_);
  and (_42824_, _36453_, _37208_);
  or (_42825_, _42824_, _42632_);
  and (_42826_, _42461_, _34793_);
  or (_42827_, _42826_, _35839_);
  or (_42828_, _42827_, _42695_);
  or (_42829_, _42828_, _42825_);
  or (_42830_, _42829_, _42456_);
  or (_42831_, _42830_, _42823_);
  and (_42832_, _42831_, _33860_);
  and (_42833_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42834_, _42833_, _42542_);
  or (_42835_, _42834_, _42832_);
  and (_30485_, _42835_, _41806_);
  nor (_42836_, _42827_, _42825_);
  nand (_42837_, _42836_, _42819_);
  or (_42838_, _36036_, _35926_);
  nor (_42839_, _42838_, _42741_);
  nand (_42840_, _42839_, _40330_);
  or (_42841_, _42759_, _42502_);
  or (_42842_, _42841_, _42840_);
  or (_42843_, _42460_, _42454_);
  or (_42844_, _42843_, _42842_);
  or (_42845_, _42844_, _42837_);
  and (_42846_, _42845_, _33860_);
  and (_42847_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42848_, _42847_, _42543_);
  or (_42849_, _42848_, _42846_);
  and (_30487_, _42849_, _41806_);
  and (_42850_, _42418_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_42851_, _36442_);
  and (_42852_, _42851_, _37208_);
  or (_42853_, _42852_, _37125_);
  or (_42854_, _42765_, _42426_);
  or (_42855_, _42854_, _42853_);
  or (_42856_, _42797_, _42753_);
  or (_42857_, _42856_, _42855_);
  or (_42858_, _42747_, _42538_);
  or (_42859_, _42858_, _42739_);
  or (_42860_, _42859_, _42857_);
  and (_42861_, _42860_, _42324_);
  or (_30489_, _42861_, _42850_);
  nor (_38811_, _34233_, rst);
  nor (_38813_, _40321_, rst);
  and (_42862_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_42864_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_42865_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_42866_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_42867_, _42866_, _42865_);
  and (_42868_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_42869_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_42870_, _42869_, _42868_);
  and (_42871_, _42870_, _42867_);
  and (_42872_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_42873_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_42874_, _42873_, _42872_);
  and (_42876_, _42874_, _42871_);
  nor (_42877_, _42876_, _33915_);
  nor (_42878_, _42877_, _42864_);
  nor (_42879_, _42878_, _40305_);
  nor (_42880_, _42879_, _42862_);
  nor (_38814_, _42880_, rst);
  nor (_38825_, _36365_, rst);
  and (_38826_, _35012_, _41806_);
  nor (_38827_, _35242_, rst);
  nor (_38828_, _35496_, rst);
  and (_38829_, _35751_, _41806_);
  nor (_38830_, _34486_, rst);
  nor (_38831_, _34727_, rst);
  nor (_38832_, _40396_, rst);
  nor (_38834_, _40606_, rst);
  nor (_38835_, _40479_, rst);
  nor (_38836_, _40356_, rst);
  nor (_38837_, _40527_, rst);
  nor (_38838_, _40458_, rst);
  nor (_38840_, _40682_, rst);
  and (_42881_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_42882_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_42883_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_42884_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42885_, _42884_, _42883_);
  and (_42886_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42887_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_42888_, _42887_, _42886_);
  and (_42889_, _42888_, _42885_);
  and (_42890_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_42891_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_42892_, _42891_, _42890_);
  and (_42893_, _42892_, _42889_);
  nor (_42894_, _42893_, _33915_);
  nor (_42895_, _42894_, _42882_);
  nor (_42896_, _42895_, _40305_);
  nor (_42897_, _42896_, _42881_);
  nor (_38841_, _42897_, rst);
  and (_42898_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_42899_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_42900_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42901_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_42902_, _42901_, _42900_);
  and (_42903_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_42904_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_42905_, _42904_, _42903_);
  and (_42906_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_42907_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_42908_, _42907_, _42906_);
  and (_42909_, _42908_, _42905_);
  and (_42910_, _42909_, _42902_);
  nor (_42911_, _42910_, _33915_);
  nor (_42912_, _42911_, _42899_);
  nor (_42913_, _42912_, _40305_);
  nor (_42914_, _42913_, _42898_);
  nor (_38842_, _42914_, rst);
  and (_42915_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_42916_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_42917_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_42918_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_42919_, _42918_, _42917_);
  and (_42920_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_42921_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_42922_, _42921_, _42920_);
  and (_42923_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_42924_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_42925_, _42924_, _42923_);
  and (_42926_, _42925_, _42922_);
  and (_42927_, _42926_, _42919_);
  nor (_42928_, _42927_, _33915_);
  nor (_42929_, _42928_, _42916_);
  nor (_42930_, _42929_, _40305_);
  nor (_42931_, _42930_, _42915_);
  nor (_38843_, _42931_, rst);
  and (_42932_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_42933_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_42934_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_42935_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_42936_, _42935_, _42934_);
  and (_42937_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_42938_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_42939_, _42938_, _42937_);
  and (_42940_, _42939_, _42936_);
  and (_42941_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_42942_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_42943_, _42942_, _42941_);
  and (_42944_, _42943_, _42940_);
  nor (_42945_, _42944_, _33915_);
  nor (_42946_, _42945_, _42933_);
  nor (_42947_, _42946_, _40305_);
  nor (_42948_, _42947_, _42932_);
  nor (_38844_, _42948_, rst);
  and (_42949_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_42950_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_42951_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_42952_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_42953_, _42952_, _42951_);
  and (_42954_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42955_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_42956_, _42955_, _42954_);
  and (_42957_, _42956_, _42953_);
  and (_42958_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_42959_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_42960_, _42959_, _42958_);
  and (_42961_, _42960_, _42957_);
  nor (_42962_, _42961_, _33915_);
  nor (_42963_, _42962_, _42950_);
  nor (_42964_, _42963_, _40305_);
  nor (_42965_, _42964_, _42949_);
  nor (_38846_, _42965_, rst);
  and (_42966_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_42967_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_42968_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_42969_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_42970_, _42969_, _42968_);
  and (_42971_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42972_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_42973_, _42972_, _42971_);
  and (_42974_, _42973_, _42970_);
  and (_42975_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_42976_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_42977_, _42976_, _42975_);
  and (_42978_, _42977_, _42974_);
  nor (_42979_, _42978_, _33915_);
  nor (_42980_, _42979_, _42967_);
  nor (_42981_, _42980_, _40305_);
  nor (_42982_, _42981_, _42966_);
  nor (_38847_, _42982_, rst);
  and (_42983_, _40305_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_42984_, _33915_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_42985_, _34047_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_42986_, _34003_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_42987_, _42986_, _42985_);
  and (_42988_, _34156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42989_, _34091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_42990_, _42989_, _42988_);
  and (_42991_, _42990_, _42987_);
  and (_42992_, _33959_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_42993_, _34124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42994_, _42993_, _42992_);
  and (_42995_, _42994_, _42991_);
  nor (_42996_, _42995_, _33915_);
  nor (_42997_, _42996_, _42984_);
  nor (_42998_, _42997_, _40305_);
  nor (_42999_, _42998_, _42983_);
  nor (_38848_, _42999_, rst);
  and (_43000_, _33881_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_43001_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_43002_, _43000_, _38571_);
  and (_43003_, _43002_, _41806_);
  and (_38872_, _43003_, _43001_);
  not (_43004_, _43000_);
  or (_43005_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _43000_, _41806_);
  and (_43006_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _41806_);
  or (_43007_, _43006_, _00000_);
  and (_38874_, _43007_, _43005_);
  nor (_38911_, _40327_, rst);
  and (_38913_, _40544_, _41806_);
  nor (_38914_, _40300_, rst);
  nor (_43008_, _40327_, _24949_);
  and (_43009_, _40327_, _24949_);
  nor (_43010_, _43009_, _43008_);
  nor (_43011_, _40703_, _24665_);
  and (_43012_, _40703_, _24665_);
  nor (_43013_, _43012_, _43011_);
  nor (_43014_, _43013_, _43010_);
  nor (_43015_, _40380_, _25112_);
  and (_43016_, _40380_, _25112_);
  nor (_43017_, _43016_, _43015_);
  not (_43018_, _43017_);
  and (_43019_, _40547_, _40614_);
  nor (_43020_, _40547_, _40614_);
  nor (_43021_, _43020_, _43019_);
  nor (_43022_, _40463_, _24796_);
  and (_43023_, _40463_, _24796_);
  nor (_43024_, _43023_, _43022_);
  nor (_43025_, _43024_, _43021_);
  and (_43026_, _43025_, _43018_);
  and (_43027_, _43026_, _43014_);
  nor (_43028_, _37539_, _42442_);
  and (_43029_, _38853_, _28087_);
  and (_43030_, _43029_, _43028_);
  and (_43031_, _43030_, _43027_);
  nor (_43032_, _25984_, _25593_);
  and (_43033_, _43032_, _28872_);
  and (_43034_, _43033_, _30240_);
  nand (_43035_, _43034_, _30914_);
  nor (_43036_, _43035_, _31652_);
  and (_43037_, _43036_, _32393_);
  nor (_43038_, _43028_, _37668_);
  and (_43039_, _43038_, _43037_);
  and (_43040_, _43039_, _26604_);
  and (_43041_, _43028_, _26354_);
  not (_43042_, _37668_);
  nor (_43043_, _43028_, _34530_);
  nor (_43044_, _43043_, _43042_);
  and (_43045_, _43044_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_43046_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_43047_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_43048_, _43047_, _43046_);
  nor (_43049_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_43050_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_43051_, _43050_, _43049_);
  and (_43052_, _43051_, _43048_);
  and (_43053_, _43052_, _36771_);
  or (_43054_, _43053_, _43045_);
  or (_43055_, _43054_, _43041_);
  nor (_43056_, _43055_, _43040_);
  not (_43057_, _42494_);
  nor (_43058_, _42694_, _37263_);
  and (_43059_, _43058_, _43057_);
  or (_43060_, _37507_, _36518_);
  or (_43061_, _43060_, _36990_);
  and (_43062_, _43061_, _36584_);
  nor (_43063_, _43062_, _42651_);
  nand (_43064_, _43063_, _43059_);
  and (_43065_, _43064_, _43056_);
  nand (_43066_, _37657_, _35795_);
  and (_43067_, _43066_, _37723_);
  or (_43068_, _43067_, _43056_);
  nor (_43069_, _42423_, _36529_);
  nand (_43070_, _43069_, _43068_);
  or (_43071_, _43070_, _43065_);
  and (_43072_, _43071_, _36749_);
  and (_43073_, _36628_, _35915_);
  nor (_43074_, _43073_, _42481_);
  nor (_43075_, _43074_, _33817_);
  nor (_43076_, _43075_, _36781_);
  not (_43077_, _43076_);
  nor (_43078_, _43077_, _43072_);
  nor (_43079_, _38955_, _38823_);
  and (_43080_, _43079_, _38860_);
  not (_43081_, _43080_);
  and (_43082_, _43081_, _43044_);
  not (_43083_, _39080_);
  and (_43084_, _43083_, _36771_);
  nor (_43085_, _43084_, _43082_);
  not (_43086_, _43085_);
  nor (_43087_, _43086_, _43078_);
  not (_43088_, _43087_);
  nor (_43089_, _43088_, _43031_);
  and (_43090_, _40611_, _30686_);
  nor (_43091_, _40611_, _30686_);
  or (_43092_, _43091_, _43090_);
  nand (_43093_, _43018_, _28076_);
  nor (_43094_, _40415_, _24434_);
  and (_43095_, _40415_, _24434_);
  nor (_43096_, _43095_, _43094_);
  nor (_43097_, _40500_, _24197_);
  and (_43098_, _40500_, _24197_);
  nor (_43099_, _43098_, _43097_);
  or (_43100_, _43099_, _43096_);
  or (_43101_, _43100_, _43093_);
  nor (_43102_, _43101_, _43092_);
  and (_43103_, _43102_, _43025_);
  and (_43104_, _43103_, _43014_);
  nor (_43105_, _24949_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_43106_, _43105_, _43104_);
  not (_43107_, _43106_);
  and (_43108_, _43107_, _43089_);
  and (_43109_, _43108_, _37635_);
  and (_38918_, _43109_, _41806_);
  and (_38919_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _41806_);
  and (_38920_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _41806_);
  nor (_43110_, _37635_, _28011_);
  and (_43111_, _36749_, _36529_);
  not (_43112_, _43111_);
  nor (_43113_, _43112_, _38582_);
  and (_43114_, _43073_, _36858_);
  and (_43115_, _43114_, _40322_);
  and (_43116_, _42650_, _37539_);
  and (_43117_, _43116_, _43058_);
  nor (_43118_, _43117_, _37679_);
  nor (_43119_, _43114_, _37624_);
  not (_43120_, _43119_);
  nor (_43121_, _43120_, _43118_);
  nor (_43122_, _43111_, _43075_);
  and (_43123_, _43122_, _43121_);
  and (_43124_, _36584_, _36858_);
  and (_43125_, _43124_, _35871_);
  not (_43126_, _37657_);
  and (_43127_, _43069_, _43126_);
  and (_43128_, _43127_, _43059_);
  and (_43129_, _43128_, _43116_);
  nor (_43130_, _43129_, _37679_);
  nor (_43131_, _43130_, _43125_);
  and (_43132_, _43131_, _43123_);
  and (_43134_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_43135_, _43134_, _43115_);
  or (_43136_, _43135_, _43113_);
  or (_43137_, _43136_, _43110_);
  not (_43138_, _42880_);
  and (_43140_, _37485_, _36858_);
  not (_43141_, _43140_);
  and (_43142_, _43141_, _43121_);
  nor (_43143_, _43142_, _43138_);
  and (_43144_, _43142_, _40321_);
  nor (_43146_, _43144_, _43143_);
  and (_43147_, _43146_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_43148_, _43147_);
  nor (_43149_, _43146_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_43150_, _43149_, _43147_);
  not (_43152_, _42999_);
  nor (_43153_, _43142_, _43152_);
  and (_43154_, _43142_, _40682_);
  nor (_43155_, _43154_, _43153_);
  and (_43156_, _43155_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_43158_, _43155_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_43159_, _43158_, _43156_);
  not (_43160_, _42982_);
  nor (_43161_, _43142_, _43160_);
  and (_43162_, _43142_, _40458_);
  nor (_43164_, _43162_, _43161_);
  and (_43165_, _43164_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_43166_, _43164_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_43167_, _42965_);
  nor (_43168_, _43142_, _43167_);
  and (_43170_, _43142_, _40527_);
  nor (_43171_, _43170_, _43168_);
  nand (_43173_, _43171_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_43174_, _42948_);
  nor (_43175_, _43142_, _43174_);
  and (_43176_, _43142_, _40356_);
  nor (_43177_, _43176_, _43175_);
  and (_43178_, _43177_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_43179_, _43177_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_43181_, _42931_);
  nor (_43182_, _43142_, _43181_);
  and (_43183_, _43142_, _40479_);
  nor (_43185_, _43183_, _43182_);
  and (_43186_, _43185_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_43187_, _42914_);
  nor (_43189_, _43142_, _43187_);
  and (_43190_, _43142_, _40606_);
  nor (_43191_, _43190_, _43189_);
  and (_43193_, _43191_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_43194_, _42897_);
  nor (_43195_, _43142_, _43194_);
  and (_43197_, _43142_, _40396_);
  nor (_43198_, _43197_, _43195_);
  and (_43199_, _43198_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_43201_, _43191_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_43202_, _43201_, _43193_);
  and (_43203_, _43202_, _43199_);
  nor (_43205_, _43203_, _43193_);
  not (_43206_, _43205_);
  nor (_43208_, _43185_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_43209_, _43208_, _43186_);
  and (_43210_, _43209_, _43206_);
  nor (_43211_, _43210_, _43186_);
  nor (_43212_, _43211_, _43179_);
  or (_43213_, _43212_, _43178_);
  or (_43214_, _43171_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43216_, _43214_, _43173_);
  nand (_43217_, _43216_, _43213_);
  and (_43218_, _43217_, _43173_);
  nor (_43220_, _43218_, _43166_);
  or (_43221_, _43220_, _43165_);
  and (_43222_, _43221_, _43159_);
  nor (_43224_, _43222_, _43156_);
  not (_43225_, _43224_);
  nand (_43226_, _43225_, _43150_);
  and (_43228_, _43226_, _43148_);
  nor (_43229_, _43228_, _38543_);
  and (_43230_, _43229_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_43232_, _43230_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_43233_, _43232_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43234_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43236_, _43234_, _43233_);
  nor (_43237_, _43236_, _43146_);
  not (_43238_, _43146_);
  and (_43240_, _43228_, _38543_);
  and (_43241_, _43240_, _38549_);
  and (_43243_, _43241_, _38554_);
  and (_43244_, _43243_, _38539_);
  nor (_43245_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43246_, _43245_, _43244_);
  nor (_43247_, _43246_, _43238_);
  nor (_43249_, _43247_, _43237_);
  or (_43250_, _43146_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43251_, _43146_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_43253_, _43251_, _43250_);
  and (_43254_, _43253_, _43249_);
  or (_43255_, _43254_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_43257_, _43254_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_43258_, _43122_);
  and (_43259_, _43258_, _43142_);
  nor (_43261_, _43131_, _43259_);
  and (_43262_, _43261_, _43257_);
  and (_43263_, _43262_, _43255_);
  or (_43265_, _43263_, _43137_);
  and (_43266_, _43121_, _43075_);
  and (_43267_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43269_, _43267_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_43270_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43271_, _43270_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_43273_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43274_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_43276_, _43274_, _43273_);
  and (_43277_, _43276_, _43271_);
  and (_43278_, _43277_, _43269_);
  and (_43279_, _43278_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43280_, _43279_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43281_, _43280_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_43282_, _43281_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43284_, _43282_, _38571_);
  or (_43285_, _43282_, _38571_);
  and (_43286_, _43285_, _43284_);
  nand (_43288_, _43286_, _43266_);
  nand (_43289_, _43288_, _43108_);
  or (_43290_, _43289_, _43265_);
  not (_43292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43293_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_43294_, _43293_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_43296_, _43294_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_43297_, _43296_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_43298_, _43297_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_43300_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_43301_, _43300_, _43298_);
  and (_43302_, _43301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_43304_, _43302_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_43305_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_43306_, _34036_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43308_, _43306_, _40305_);
  nor (_43309_, _43308_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_43311_, _43309_);
  and (_43312_, _43311_, _43305_);
  and (_43313_, _43312_, _43304_);
  nand (_43314_, _43313_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_43316_, _43314_, _43292_);
  or (_43317_, _43314_, _43292_);
  and (_43318_, _43317_, _43316_);
  or (_43320_, _43318_, _43108_);
  and (_43321_, _43320_, _41806_);
  and (_38922_, _43321_, _43290_);
  and (_43323_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _41806_);
  and (_43324_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_43325_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_43327_, _33860_, _43325_);
  not (_43328_, _43327_);
  not (_43329_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_43331_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_43332_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_43333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_43335_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_43336_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_43337_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_43339_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_43340_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_43342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43343_, _43342_, _43340_);
  and (_43344_, _43343_, _43339_);
  and (_43345_, _43344_, _43337_);
  and (_43347_, _43345_, _43336_);
  and (_43348_, _43347_, _43335_);
  and (_43349_, _43348_, _43333_);
  and (_43351_, _43349_, _43332_);
  and (_43352_, _43351_, _43331_);
  and (_43353_, _43352_, _43329_);
  nor (_43355_, _43353_, _43292_);
  and (_43356_, _43353_, _43292_);
  nor (_43357_, _43356_, _43355_);
  nor (_43359_, _43352_, _43329_);
  or (_43360_, _43359_, _43353_);
  and (_43361_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_43363_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_43364_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43365_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_43367_, _43365_, _43363_);
  and (_43368_, _43367_, _43364_);
  nor (_43369_, _43368_, _43363_);
  nor (_43371_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43372_, _43371_, _43361_);
  not (_43374_, _43372_);
  nor (_43375_, _43374_, _43369_);
  nor (_43376_, _43375_, _43361_);
  not (_43377_, _43376_);
  and (_43379_, _43377_, _43349_);
  and (_43380_, _43379_, _43332_);
  and (_43381_, _43380_, _43331_);
  and (_43383_, _43381_, _43360_);
  nor (_43384_, _43381_, _43360_);
  or (_43385_, _43384_, _43383_);
  not (_43387_, _43385_);
  and (_43388_, _43376_, _43352_);
  and (_43389_, _43376_, _43351_);
  nor (_43391_, _43389_, _43331_);
  nor (_43392_, _43391_, _43388_);
  not (_43393_, _43392_);
  and (_43395_, _43376_, _43349_);
  nor (_43396_, _43395_, _43332_);
  nor (_43397_, _43396_, _43389_);
  not (_43399_, _43397_);
  and (_43400_, _43376_, _43347_);
  and (_43401_, _43400_, _43335_);
  nor (_43403_, _43401_, _43333_);
  nor (_43404_, _43403_, _43395_);
  not (_43406_, _43404_);
  nor (_43407_, _43400_, _43335_);
  nor (_43408_, _43407_, _43401_);
  not (_43409_, _43408_);
  not (_43410_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_43411_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_43412_, _43376_, _43345_);
  and (_43414_, _43412_, _43411_);
  nor (_43415_, _43414_, _43410_);
  nor (_43416_, _43415_, _43400_);
  not (_43418_, _43416_);
  and (_43419_, _43376_, _43343_);
  and (_43420_, _43419_, _43339_);
  nor (_43422_, _43420_, _43337_);
  nor (_43423_, _43422_, _43412_);
  not (_43424_, _43423_);
  nor (_43426_, _43419_, _43339_);
  nor (_43427_, _43426_, _43420_);
  not (_43428_, _43427_);
  and (_43430_, _43376_, _43342_);
  nor (_43431_, _43430_, _43340_);
  nor (_43432_, _43431_, _43419_);
  not (_43434_, _43432_);
  not (_43435_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43436_, _43376_, _43435_);
  nor (_43438_, _43376_, _43435_);
  nor (_43439_, _43438_, _43436_);
  not (_43441_, _43439_);
  nor (_43442_, _42372_, _42340_);
  not (_43443_, _42372_);
  nor (_43444_, _42367_, _42355_);
  nor (_43446_, _43444_, _43443_);
  nor (_43447_, _43446_, _42396_);
  or (_43448_, _43447_, _43442_);
  and (_43450_, _42354_, _42366_);
  not (_43451_, _43450_);
  nor (_43452_, _42372_, _42368_);
  nor (_43454_, _43452_, _43451_);
  not (_43455_, _42369_);
  and (_43456_, _42387_, _42330_);
  nor (_43458_, _43456_, _42348_);
  nor (_43459_, _43458_, _43455_);
  nor (_43460_, _43459_, _43454_);
  and (_43462_, _43460_, _43448_);
  and (_43463_, _42343_, _42330_);
  nor (_43464_, _43463_, _42359_);
  nor (_43466_, _43464_, _43443_);
  and (_43467_, _42372_, _42334_);
  and (_43468_, _43467_, _42345_);
  nor (_43470_, _43468_, _43466_);
  and (_43471_, _42396_, _42357_);
  nor (_43473_, _43471_, _42364_);
  not (_43474_, _43473_);
  not (_43475_, _42361_);
  and (_43476_, _42335_, _35496_);
  and (_43478_, _43476_, _42334_);
  and (_43479_, _42354_, _42329_);
  and (_43483_, _35751_, _35496_);
  and (_43489_, _43483_, _43479_);
  nor (_43490_, _43489_, _43478_);
  nor (_43503_, _43490_, _43475_);
  nor (_43508_, _43503_, _43474_);
  and (_43509_, _43508_, _43470_);
  and (_43523_, _43509_, _43462_);
  and (_43528_, _42359_, _42340_);
  not (_43529_, _43528_);
  nor (_43541_, _42370_, _42350_);
  and (_43548_, _43541_, _43529_);
  nor (_43549_, _42355_, _42376_);
  nor (_43559_, _43549_, _43455_);
  not (_43568_, _43559_);
  not (_43569_, _42368_);
  and (_43577_, _42366_, _42334_);
  nor (_43586_, _43577_, _42388_);
  nor (_43587_, _43586_, _43569_);
  not (_43597_, _42347_);
  and (_43598_, _42387_, _42334_);
  and (_43605_, _42330_, _34486_);
  nor (_43616_, _43605_, _43598_);
  nor (_43622_, _43616_, _43597_);
  nor (_43623_, _43622_, _43587_);
  and (_43636_, _43623_, _43568_);
  and (_43641_, _43636_, _43548_);
  and (_43642_, _43641_, _43523_);
  not (_43656_, _43598_);
  and (_43661_, _43549_, _43656_);
  nor (_43662_, _43661_, _35496_);
  not (_43668_, _43662_);
  and (_43680_, _42344_, _42330_);
  not (_43681_, _43680_);
  nor (_43693_, _43463_, _42396_);
  and (_43700_, _43693_, _43681_);
  nor (_43701_, _43700_, _43455_);
  not (_43711_, _43701_);
  and (_43720_, _43711_, _42399_);
  and (_43721_, _43720_, _43668_);
  and (_43722_, _43467_, _42343_);
  not (_43724_, _43722_);
  and (_43725_, _43724_, _42379_);
  and (_43727_, _42369_, _42359_);
  and (_43728_, _43450_, _42357_);
  nor (_43729_, _43728_, _43727_);
  and (_43730_, _42371_, _42341_);
  not (_43731_, _43730_);
  and (_43733_, _43731_, _43729_);
  and (_43734_, _43733_, _43725_);
  and (_43735_, _42394_, _42340_);
  not (_43737_, _43735_);
  and (_43738_, _42388_, _42328_);
  and (_43739_, _42355_, _42340_);
  nor (_43741_, _43739_, _43738_);
  and (_43742_, _43741_, _43737_);
  and (_43743_, _43577_, _42347_);
  and (_43745_, _42359_, _42347_);
  nor (_43746_, _43745_, _43743_);
  and (_43747_, _43746_, _42384_);
  and (_43749_, _43747_, _43742_);
  and (_43750_, _43749_, _43734_);
  and (_43751_, _43750_, _43721_);
  and (_43753_, _43751_, _43642_);
  nor (_43754_, _43367_, _43364_);
  nor (_43755_, _43754_, _43368_);
  not (_43757_, _43755_);
  nor (_43758_, _43757_, _43753_);
  and (_43760_, _43729_, _43548_);
  nor (_43761_, _42383_, _42364_);
  and (_43762_, _43761_, _43568_);
  nor (_43763_, _43471_, _42395_);
  and (_43765_, _42388_, _42357_);
  nor (_43766_, _43765_, _43743_);
  and (_43767_, _43766_, _43763_);
  and (_43769_, _43767_, _43762_);
  and (_43770_, _43769_, _43760_);
  not (_43771_, _43770_);
  nor (_43773_, _43771_, _43753_);
  not (_43774_, _43773_);
  nor (_43775_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43777_, _43775_, _43364_);
  and (_43778_, _43777_, _43774_);
  and (_43779_, _43757_, _43753_);
  nor (_43781_, _43779_, _43758_);
  and (_43782_, _43781_, _43778_);
  nor (_43783_, _43782_, _43758_);
  not (_43785_, _43783_);
  and (_43786_, _43374_, _43369_);
  nor (_43787_, _43786_, _43375_);
  and (_43789_, _43787_, _43785_);
  and (_43790_, _43789_, _43441_);
  not (_43792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_43793_, _43436_, _43792_);
  or (_43794_, _43793_, _43430_);
  and (_43795_, _43794_, _43790_);
  and (_43797_, _43795_, _43434_);
  and (_43798_, _43797_, _43428_);
  and (_43799_, _43798_, _43424_);
  nor (_43801_, _43412_, _43411_);
  or (_43802_, _43801_, _43414_);
  and (_43803_, _43802_, _43799_);
  and (_43805_, _43803_, _43418_);
  and (_43806_, _43805_, _43409_);
  and (_43807_, _43806_, _43406_);
  and (_43809_, _43807_, _43399_);
  and (_43810_, _43809_, _43393_);
  and (_43811_, _43810_, _43387_);
  or (_43813_, _43811_, _43383_);
  nor (_43814_, _43813_, _43357_);
  and (_43815_, _43813_, _43357_);
  or (_43817_, _43815_, _43814_);
  or (_43818_, _43817_, _43328_);
  or (_43819_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_43821_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_43822_, _43821_, _43819_);
  and (_43824_, _43822_, _43818_);
  or (_38923_, _43824_, _43324_);
  nor (_43825_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_38924_, _43825_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_38925_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _41806_);
  nor (_43827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_43828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_43830_, _43828_, _43827_);
  nor (_43831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_43832_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_43834_, _43832_, _43831_);
  and (_43835_, _43834_, _43830_);
  nor (_43836_, _43835_, rst);
  and (_43838_, \oc8051_top_1.oc8051_rom1.ea_int , _33828_);
  nand (_43839_, _43838_, _33860_);
  and (_43840_, _43839_, _38925_);
  or (_38927_, _43840_, _43836_);
  and (_43842_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_43843_, _43842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_38928_, _43843_, _41806_);
  nor (_43845_, _43309_, _40305_);
  nor (_43846_, _43753_, _33981_);
  nor (_43848_, _43773_, _34069_);
  and (_43849_, _43753_, _33981_);
  nor (_43850_, _43849_, _43846_);
  and (_43851_, _43850_, _43848_);
  nor (_43852_, _43851_, _43846_);
  nor (_43853_, _43852_, _40305_);
  and (_43854_, _43853_, _33937_);
  nor (_43855_, _43853_, _33937_);
  nor (_43856_, _43855_, _43854_);
  nor (_43857_, _43856_, _43845_);
  and (_43858_, _33992_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_43859_, _43858_, _43845_);
  nor (_43860_, _43859_, _43770_);
  or (_43861_, _43860_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_43862_, _43861_, _43857_);
  and (_38929_, _43862_, _41806_);
  not (_43863_, _34935_);
  and (_43864_, _34190_, _43863_);
  not (_43865_, _35685_);
  and (_43866_, _43865_, _34683_);
  and (_43867_, _43866_, _43864_);
  and (_43868_, _33881_, _41806_);
  nand (_43869_, _43868_, _35199_);
  nor (_43870_, _43869_, _35451_);
  not (_43871_, _34442_);
  nor (_43872_, _36321_, _43871_);
  and (_43873_, _43872_, _43870_);
  and (_38932_, _43873_, _43867_);
  nor (_43874_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_43875_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_43876_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_38935_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _41806_);
  and (_43877_, _38935_, _43876_);
  or (_38934_, _43877_, _43875_);
  not (_43878_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_43879_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43880_, _43879_, _43878_);
  and (_43881_, _43879_, _43878_);
  nor (_43882_, _43881_, _43880_);
  not (_43883_, _43882_);
  and (_43884_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_43885_, _43884_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43886_, _43884_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_43887_, _43886_, _43885_);
  or (_43888_, _43887_, _43879_);
  and (_43889_, _43888_, _43883_);
  nor (_43890_, _43880_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_43891_, _43880_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_43892_, _43891_, _43890_);
  or (_43893_, _43885_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_38937_, _43893_, _41806_);
  and (_43894_, _38937_, _43892_);
  and (_38936_, _43894_, _43889_);
  not (_43895_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_43896_, _43309_, _43895_);
  and (_43897_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_43898_, _43896_);
  and (_43899_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_43900_, _43899_, _43897_);
  and (_38938_, _43900_, _41806_);
  and (_43901_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_43902_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_43903_, _43902_, _43901_);
  and (_38939_, _43903_, _41806_);
  and (_43904_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_43905_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_43906_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _43905_);
  and (_43907_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_43908_, _43907_, _43904_);
  and (_38940_, _43908_, _41806_);
  and (_43909_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_43910_, _43909_, _43906_);
  and (_38941_, _43910_, _41806_);
  or (_43911_, _43905_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_38942_, _43911_, _41806_);
  not (_43912_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_43913_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_43914_, _43913_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_43915_, _43905_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_43916_, _43915_, _41806_);
  and (_38943_, _43916_, _43914_);
  or (_43917_, _43905_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_38944_, _43917_, _41806_);
  nor (_43918_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_43919_, _43918_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_43920_, _43919_, _41806_);
  and (_43921_, _38935_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_38945_, _43921_, _43920_);
  and (_43922_, _43895_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_43923_, _43922_, _43919_);
  and (_38946_, _43923_, _41806_);
  nand (_43924_, _43919_, _38582_);
  or (_43925_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_43926_, _43925_, _41806_);
  and (_38947_, _43926_, _43924_);
  and (_38948_, _37965_, _40269_);
  or (_43927_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_43928_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _41806_);
  or (_43929_, _43928_, _00000_);
  and (_38985_, _43929_, _43927_);
  or (_43930_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_43931_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_43932_, _43000_, _43931_);
  and (_43933_, _43932_, _41806_);
  and (_38986_, _43933_, _43930_);
  or (_43934_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_43935_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_43936_, _43000_, _43935_);
  and (_43937_, _43936_, _41806_);
  and (_38987_, _43937_, _43934_);
  or (_43938_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_43939_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_43940_, _43000_, _43939_);
  and (_43941_, _43940_, _41806_);
  and (_38989_, _43941_, _43938_);
  or (_43942_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_43943_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_43944_, _43000_, _43943_);
  and (_43945_, _43944_, _41806_);
  and (_38990_, _43945_, _43942_);
  or (_43946_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_43947_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_43948_, _43000_, _43947_);
  and (_43949_, _43948_, _41806_);
  and (_38991_, _43949_, _43946_);
  or (_43950_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_43951_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_43952_, _43000_, _43951_);
  and (_43953_, _43952_, _41806_);
  and (_38992_, _43953_, _43950_);
  or (_43954_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_43955_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_43956_, _43000_, _43955_);
  and (_43957_, _43956_, _41806_);
  and (_38993_, _43957_, _43954_);
  or (_43958_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_43959_, _43000_, _38543_);
  and (_43960_, _43959_, _41806_);
  and (_38994_, _43960_, _43958_);
  or (_43961_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_43962_, _43000_, _38549_);
  and (_43963_, _43962_, _41806_);
  and (_38995_, _43963_, _43961_);
  or (_43964_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_43965_, _43000_, _38554_);
  and (_43966_, _43965_, _41806_);
  and (_38996_, _43966_, _43964_);
  or (_43967_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_43968_, _43000_, _38539_);
  and (_43969_, _43968_, _41806_);
  and (_38997_, _43969_, _43967_);
  or (_43970_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_43971_, _43000_, _38560_);
  and (_43972_, _43971_, _41806_);
  and (_38998_, _43972_, _43970_);
  or (_43973_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_43974_, _43000_, _38535_);
  and (_43975_, _43974_, _41806_);
  and (_39000_, _43975_, _43973_);
  or (_43976_, _43000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_43977_, _43000_, _38566_);
  and (_43978_, _43977_, _41806_);
  and (_39001_, _43978_, _43976_);
  or (_43979_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_43980_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _41806_);
  or (_43981_, _43980_, _00000_);
  and (_39005_, _43981_, _43979_);
  or (_43982_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_43983_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _41806_);
  or (_43984_, _43983_, _00000_);
  and (_39006_, _43984_, _43982_);
  or (_43985_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_43986_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _41806_);
  or (_43987_, _43986_, _00000_);
  and (_39007_, _43987_, _43985_);
  or (_43988_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_43989_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _41806_);
  or (_43990_, _43989_, _00000_);
  and (_39008_, _43990_, _43988_);
  or (_43991_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_43992_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _41806_);
  or (_43993_, _43992_, _00000_);
  and (_39009_, _43993_, _43991_);
  or (_43994_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_43995_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _41806_);
  or (_43996_, _43995_, _00000_);
  and (_39010_, _43996_, _43994_);
  or (_43997_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_43998_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _41806_);
  or (_43999_, _43998_, _00000_);
  and (_39011_, _43999_, _43997_);
  or (_44000_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_44001_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _41806_);
  or (_44002_, _44001_, _00000_);
  and (_39012_, _44002_, _44000_);
  or (_44003_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_44004_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _41806_);
  or (_44005_, _44004_, _00000_);
  and (_39013_, _44005_, _44003_);
  or (_44006_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_44007_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _41806_);
  or (_44008_, _44007_, _00000_);
  and (_39014_, _44008_, _44006_);
  or (_44009_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_44010_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _41806_);
  or (_44011_, _44010_, _00000_);
  and (_39015_, _44011_, _44009_);
  or (_44012_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_44013_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _41806_);
  or (_44014_, _44013_, _00000_);
  and (_39016_, _44014_, _44012_);
  or (_44015_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_44016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _41806_);
  or (_44017_, _44016_, _00000_);
  and (_39017_, _44017_, _44015_);
  or (_44018_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_44019_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _41806_);
  or (_44020_, _44019_, _00000_);
  and (_39018_, _44020_, _44018_);
  or (_44021_, _43004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_44022_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _41806_);
  or (_44023_, _44022_, _00000_);
  and (_39019_, _44023_, _44021_);
  and (_44024_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_44025_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_44026_, _44025_, _44024_);
  and (_39197_, _44026_, _41806_);
  and (_44027_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_44028_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_44029_, _44028_, _44027_);
  and (_39198_, _44029_, _41806_);
  and (_44030_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_44031_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_44032_, _44031_, _44030_);
  and (_39199_, _44032_, _41806_);
  and (_44033_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_44034_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_44035_, _44034_, _43896_);
  or (_44036_, _44035_, _44033_);
  and (_39200_, _44036_, _41806_);
  and (_44037_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_44038_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_44039_, _44038_, _44037_);
  and (_39201_, _44039_, _41806_);
  and (_44040_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_44041_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_44042_, _44041_, _44040_);
  and (_39202_, _44042_, _41806_);
  and (_44043_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_44044_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_44045_, _44044_, _43896_);
  or (_44046_, _44045_, _44043_);
  and (_39204_, _44046_, _41806_);
  and (_44047_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_44048_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_44049_, _44048_, _44047_);
  and (_39205_, _44049_, _41806_);
  and (_44050_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_44051_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_44052_, _44051_, _44050_);
  and (_39206_, _44052_, _41806_);
  and (_44053_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_44054_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_44055_, _44054_, _44053_);
  and (_39207_, _44055_, _41806_);
  and (_44056_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_44057_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_44058_, _44057_, _44056_);
  and (_39208_, _44058_, _41806_);
  and (_44059_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_44060_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_00008_, _44060_, _44059_);
  and (_39209_, _00008_, _41806_);
  and (_00009_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_00010_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_00011_, _00010_, _00009_);
  and (_39210_, _00011_, _41806_);
  and (_00012_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_00013_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_00014_, _00013_, _00012_);
  and (_39211_, _00014_, _41806_);
  and (_00015_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_00016_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_00017_, _00016_, _00015_);
  and (_39212_, _00017_, _41806_);
  and (_00018_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_00019_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_00020_, _00019_, _00018_);
  and (_39213_, _00020_, _41806_);
  and (_00021_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_00022_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_00023_, _00022_, _00021_);
  and (_39215_, _00023_, _41806_);
  and (_00024_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_00025_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_00026_, _00025_, _00024_);
  and (_39216_, _00026_, _41806_);
  and (_00027_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_00028_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_00029_, _00028_, _00027_);
  and (_39217_, _00029_, _41806_);
  and (_00030_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_00031_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_00032_, _00031_, _00030_);
  and (_39218_, _00032_, _41806_);
  and (_00033_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_00034_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_00035_, _00034_, _00033_);
  and (_39219_, _00035_, _41806_);
  and (_00036_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_00037_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_00038_, _00037_, _00036_);
  and (_39220_, _00038_, _41806_);
  and (_00039_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_00040_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_00041_, _00040_, _00039_);
  and (_39221_, _00041_, _41806_);
  and (_00042_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_00043_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_00044_, _00043_, _00042_);
  and (_39222_, _00044_, _41806_);
  and (_00045_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_00046_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_00047_, _00046_, _00045_);
  and (_39223_, _00047_, _41806_);
  and (_00048_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_00049_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_00050_, _00049_, _00048_);
  and (_39224_, _00050_, _41806_);
  and (_00051_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_00052_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_00053_, _00052_, _00051_);
  and (_39226_, _00053_, _41806_);
  and (_00054_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_00055_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_00056_, _00055_, _00054_);
  and (_39227_, _00056_, _41806_);
  and (_00057_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_00058_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_00059_, _00058_, _00057_);
  and (_39228_, _00059_, _41806_);
  and (_00060_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_00061_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_00062_, _00061_, _00060_);
  and (_39229_, _00062_, _41806_);
  and (_00063_, _43896_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_00064_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_00065_, _00064_, _00063_);
  and (_39230_, _00065_, _41806_);
  nor (_39231_, _36409_, rst);
  nor (_39232_, _35056_, rst);
  nor (_39233_, _35286_, rst);
  nor (_39234_, _40279_, rst);
  nor (_39236_, _40408_, rst);
  nor (_39237_, _40564_, rst);
  nor (_39238_, _40492_, rst);
  nor (_39239_, _40370_, rst);
  and (_39240_, _40540_, _41806_);
  nor (_39242_, _40442_, rst);
  nor (_39243_, _40639_, rst);
  and (_39259_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _41806_);
  and (_39260_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _41806_);
  and (_39261_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _41806_);
  and (_39263_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _41806_);
  and (_39264_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _41806_);
  and (_39265_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _41806_);
  and (_39266_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _41806_);
  or (_00066_, _43132_, _43111_);
  and (_00067_, _00066_, _29242_);
  and (_00068_, _43266_, _40397_);
  and (_00069_, _43114_, _43194_);
  or (_00070_, _00069_, _00068_);
  and (_00071_, _37624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00072_, _00071_, _00070_);
  or (_00073_, _00072_, _00067_);
  nor (_00074_, _43198_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00075_, _00074_, _43199_);
  nand (_00076_, _00075_, _43261_);
  nand (_00077_, _00076_, _43108_);
  or (_00078_, _00077_, _00073_);
  or (_00079_, _43108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00080_, _00079_, _41806_);
  and (_39267_, _00080_, _00078_);
  not (_00081_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_00082_, _43109_, _00081_);
  and (_00083_, _43114_, _43187_);
  and (_00084_, _43266_, _40607_);
  or (_00085_, _00084_, _00083_);
  or (_00086_, _43202_, _43199_);
  not (_00087_, _43261_);
  nor (_00088_, _00087_, _43203_);
  and (_00089_, _00088_, _00086_);
  or (_00090_, _00089_, _00085_);
  and (_00091_, _00066_, _29904_);
  or (_00092_, _00091_, _00090_);
  and (_00093_, _00092_, _43108_);
  or (_00094_, _00093_, _00082_);
  and (_39268_, _00094_, _41806_);
  and (_00095_, _00066_, _30578_);
  and (_00096_, _43266_, _40480_);
  and (_00097_, _43114_, _43181_);
  or (_00098_, _00097_, _00096_);
  or (_00099_, _43209_, _43206_);
  nor (_00100_, _00087_, _43210_);
  and (_00101_, _00100_, _00099_);
  or (_00102_, _00101_, _00098_);
  and (_00103_, _37624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00104_, _00103_, _00102_);
  nand (_00105_, _00104_, _43108_);
  or (_00106_, _00105_, _00095_);
  not (_00107_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00108_, _43309_, _00107_);
  and (_00109_, _43309_, _00107_);
  nor (_00110_, _00109_, _00108_);
  or (_00111_, _00110_, _43108_);
  and (_00112_, _00111_, _41806_);
  and (_39269_, _00112_, _00106_);
  and (_00113_, _00066_, _31349_);
  and (_00114_, _43266_, _40357_);
  and (_00115_, _43114_, _43174_);
  or (_00116_, _00115_, _00114_);
  and (_00117_, _37624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_00118_, _00117_, _00116_);
  or (_00119_, _43179_, _43178_);
  or (_00120_, _00119_, _43211_);
  nand (_00121_, _00119_, _43211_);
  and (_00122_, _00121_, _00120_);
  and (_00123_, _00122_, _43261_);
  nor (_00124_, _00123_, _00118_);
  nand (_00125_, _00124_, _43108_);
  or (_00126_, _00125_, _00113_);
  and (_00127_, _00108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00128_, _00108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00129_, _00128_, _00127_);
  or (_00130_, _00129_, _43108_);
  and (_00131_, _00130_, _41806_);
  and (_39270_, _00131_, _00126_);
  and (_00132_, _00066_, _32055_);
  and (_00133_, _43266_, _40528_);
  and (_00134_, _43114_, _43167_);
  and (_00135_, _36792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00136_, _00135_, _00134_);
  or (_00137_, _00136_, _00133_);
  or (_00138_, _00137_, _00132_);
  or (_00139_, _43216_, _43213_);
  and (_00140_, _00139_, _43217_);
  nand (_00141_, _00140_, _43261_);
  nand (_00142_, _00141_, _43108_);
  or (_00143_, _00142_, _00138_);
  and (_00144_, _43294_, _43311_);
  nor (_00145_, _00127_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00146_, _00145_, _00144_);
  or (_00147_, _00146_, _43108_);
  and (_00148_, _00147_, _41806_);
  and (_39271_, _00148_, _00143_);
  and (_00149_, _00066_, _32864_);
  and (_00150_, _43266_, _40459_);
  and (_00151_, _43114_, _43160_);
  and (_00152_, _36792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00153_, _00152_, _00151_);
  or (_00154_, _00153_, _00150_);
  or (_00155_, _00154_, _00149_);
  or (_00156_, _43165_, _43166_);
  or (_00157_, _00156_, _43218_);
  nand (_00158_, _00156_, _43218_);
  and (_00159_, _00158_, _00157_);
  nand (_00160_, _00159_, _43261_);
  nand (_00161_, _00160_, _43108_);
  or (_00162_, _00161_, _00155_);
  and (_00163_, _43296_, _43311_);
  nor (_00164_, _00144_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00165_, _00164_, _00163_);
  or (_00166_, _00165_, _43108_);
  and (_00167_, _00166_, _41806_);
  and (_39272_, _00167_, _00162_);
  not (_00168_, _43108_);
  nor (_00169_, _43221_, _43159_);
  nor (_00170_, _00169_, _43222_);
  and (_00171_, _00170_, _43261_);
  and (_00172_, _00066_, _33609_);
  and (_00173_, _43266_, _40683_);
  and (_00174_, _43114_, _43152_);
  and (_00175_, _36792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00176_, _00175_, _00174_);
  or (_00177_, _00176_, _00173_);
  or (_00178_, _00177_, _00172_);
  or (_00179_, _00178_, _00171_);
  or (_00180_, _00179_, _00168_);
  and (_00181_, _00163_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00182_, _00163_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00183_, _00182_, _00181_);
  or (_00184_, _00183_, _43108_);
  and (_00185_, _00184_, _41806_);
  and (_39274_, _00185_, _00180_);
  and (_00186_, _00066_, _28022_);
  and (_00187_, _43266_, _40322_);
  and (_00188_, _43114_, _43138_);
  and (_00189_, _36792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_00190_, _00189_, _00188_);
  or (_00191_, _00190_, _00187_);
  or (_00192_, _43225_, _43150_);
  and (_00193_, _00192_, _43226_);
  and (_00194_, _00193_, _43261_);
  or (_00195_, _00194_, _00191_);
  or (_00196_, _00195_, _00186_);
  or (_00197_, _00196_, _00168_);
  and (_00198_, _00181_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00199_, _00181_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00200_, _00199_, _00198_);
  or (_00201_, _00200_, _43108_);
  and (_00202_, _00201_, _41806_);
  and (_39275_, _00202_, _00197_);
  nor (_00203_, _37635_, _29231_);
  nor (_00204_, _43112_, _38617_);
  and (_00205_, _43114_, _40397_);
  and (_00206_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00207_, _00206_, _00205_);
  and (_00208_, _43266_, _42329_);
  nor (_00209_, _43228_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00210_, _43228_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_00211_, _00210_, _00209_);
  or (_00212_, _00211_, _43238_);
  nand (_00213_, _00211_, _43238_);
  and (_00214_, _00213_, _43261_);
  and (_00215_, _00214_, _00212_);
  or (_00216_, _00215_, _00208_);
  or (_00217_, _00216_, _00207_);
  or (_00218_, _00217_, _00204_);
  or (_00219_, _00218_, _00203_);
  or (_00220_, _00219_, _00168_);
  and (_00221_, _00198_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00222_, _00198_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00223_, _00222_, _00221_);
  or (_00224_, _00223_, _43108_);
  and (_00225_, _00224_, _41806_);
  and (_39276_, _00225_, _00220_);
  nor (_00226_, _43112_, _38645_);
  and (_00227_, _43266_, _42353_);
  and (_00228_, _43114_, _40607_);
  and (_00229_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_00230_, _00229_, _00228_);
  or (_00231_, _00230_, _00227_);
  or (_00232_, _00231_, _00226_);
  nor (_00233_, _37635_, _29893_);
  or (_00234_, _00233_, _00232_);
  and (_00235_, _43240_, _43146_);
  and (_00236_, _43229_, _43238_);
  nor (_00237_, _00236_, _00235_);
  nor (_00238_, _00237_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00239_, _00237_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_00240_, _00239_, _00238_);
  and (_00241_, _00240_, _43261_);
  or (_00242_, _00241_, _00168_);
  or (_00243_, _00242_, _00234_);
  and (_00244_, _43301_, _43311_);
  nor (_00245_, _00221_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00246_, _00245_, _00244_);
  or (_00247_, _00246_, _43108_);
  and (_00248_, _00247_, _41806_);
  and (_39277_, _00248_, _00243_);
  or (_00249_, _37635_, _30567_);
  or (_00250_, _43112_, _38673_);
  nand (_00251_, _43114_, _40480_);
  nand (_00252_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00253_, _00252_, _00251_);
  and (_00254_, _00253_, _00250_);
  nand (_00255_, _43266_, _42333_);
  and (_00256_, _43241_, _43146_);
  and (_00257_, _43230_, _43238_);
  nor (_00258_, _00257_, _00256_);
  nor (_00259_, _00258_, _38554_);
  and (_00260_, _00258_, _38554_);
  or (_00261_, _00260_, _00087_);
  or (_00262_, _00261_, _00259_);
  and (_00263_, _00262_, _00255_);
  and (_00264_, _00263_, _00254_);
  and (_00265_, _00264_, _00249_);
  nand (_00266_, _00265_, _43108_);
  and (_00267_, _00244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00268_, _00244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00269_, _00268_, _00267_);
  or (_00270_, _00269_, _43108_);
  and (_00271_, _00270_, _41806_);
  and (_39278_, _00271_, _00266_);
  nor (_00272_, _43278_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00273_, _00272_, _43279_);
  and (_00274_, _00273_, _43266_);
  and (_00275_, _43232_, _43238_);
  and (_00276_, _43243_, _43146_);
  nor (_00277_, _00276_, _00275_);
  or (_00278_, _00277_, _38539_);
  nand (_00279_, _00277_, _38539_);
  and (_00280_, _00279_, _43261_);
  and (_00281_, _00280_, _00278_);
  nor (_00282_, _37635_, _31338_);
  nor (_00283_, _43112_, _38702_);
  and (_00284_, _43114_, _40357_);
  and (_00285_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_00286_, _00285_, _00284_);
  or (_00287_, _00286_, _00283_);
  or (_00288_, _00287_, _00282_);
  or (_00289_, _00288_, _00281_);
  or (_00290_, _00289_, _00274_);
  or (_00291_, _00290_, _00168_);
  and (_00292_, _00267_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00293_, _00267_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00294_, _00293_, _00292_);
  or (_00295_, _00294_, _43108_);
  and (_00296_, _00295_, _41806_);
  and (_39279_, _00296_, _00291_);
  and (_00297_, _43233_, _43238_);
  and (_00298_, _43244_, _43146_);
  nor (_00299_, _00298_, _00297_);
  or (_00300_, _00299_, _38560_);
  nand (_00301_, _00299_, _38560_);
  and (_00302_, _00301_, _43261_);
  and (_00303_, _00302_, _00300_);
  nor (_00304_, _43279_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00305_, _00304_, _43280_);
  and (_00306_, _00305_, _43266_);
  nor (_00307_, _37635_, _32044_);
  nor (_00308_, _43112_, _38731_);
  and (_00309_, _43114_, _40528_);
  and (_00310_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_00311_, _00310_, _00309_);
  or (_00312_, _00311_, _00308_);
  or (_00313_, _00312_, _00307_);
  or (_00314_, _00313_, _00306_);
  or (_00315_, _00314_, _00303_);
  or (_00316_, _00315_, _00168_);
  and (_00317_, _00292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00318_, _00292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00319_, _00318_, _00317_);
  or (_00320_, _00319_, _43108_);
  and (_00321_, _00320_, _41806_);
  and (_39280_, _00321_, _00316_);
  nor (_00322_, _37635_, _32853_);
  nor (_00323_, _43112_, _38760_);
  and (_00324_, _43114_, _40459_);
  and (_00325_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00326_, _00325_, _00324_);
  or (_00327_, _00326_, _00323_);
  or (_00328_, _00327_, _00322_);
  and (_00329_, _00297_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00330_, _00298_, _38560_);
  nor (_00331_, _00330_, _00329_);
  nand (_00332_, _00331_, _38535_);
  or (_00333_, _00331_, _38535_);
  and (_00334_, _00333_, _00332_);
  and (_00335_, _00334_, _43261_);
  or (_00336_, _00335_, _00328_);
  nor (_00337_, _43280_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00338_, _00337_, _43281_);
  nand (_00339_, _00338_, _43266_);
  nand (_00340_, _00339_, _43108_);
  or (_00341_, _00340_, _00336_);
  or (_00342_, _00317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_00343_, _00317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_00344_, _00343_, _00342_);
  or (_00345_, _00344_, _43108_);
  and (_00346_, _00345_, _41806_);
  and (_39281_, _00346_, _00341_);
  or (_00347_, _43281_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00348_, _00347_, _43282_);
  nand (_00349_, _00348_, _43266_);
  or (_00350_, _37635_, _33598_);
  or (_00351_, _43112_, _38787_);
  nand (_00352_, _43114_, _40683_);
  nand (_00353_, _43132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00354_, _00353_, _00352_);
  and (_00355_, _00354_, _00351_);
  and (_00356_, _00355_, _00350_);
  or (_00357_, _43249_, _38566_);
  nand (_00358_, _43249_, _38566_);
  and (_00359_, _00358_, _00357_);
  or (_00360_, _00359_, _00087_);
  and (_00361_, _00360_, _00356_);
  and (_00362_, _00361_, _00349_);
  nand (_00363_, _00362_, _43108_);
  or (_00364_, _43313_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00365_, _00364_, _43314_);
  or (_00366_, _00365_, _43108_);
  and (_00367_, _00366_, _41806_);
  and (_39282_, _00367_, _00363_);
  and (_00368_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_00369_, _43777_, _43774_);
  nor (_00370_, _00369_, _43778_);
  or (_00371_, _00370_, _43328_);
  or (_00372_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00373_, _00372_, _43821_);
  and (_00374_, _00373_, _00371_);
  or (_39283_, _00374_, _00368_);
  nor (_00375_, _43781_, _43778_);
  nor (_00376_, _00375_, _43782_);
  or (_00377_, _00376_, _43328_);
  or (_00378_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00379_, _00378_, _43821_);
  and (_00380_, _00379_, _00377_);
  and (_00381_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39285_, _00381_, _00380_);
  and (_00382_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00383_, _43787_, _43785_);
  nor (_00384_, _00383_, _43789_);
  or (_00385_, _00384_, _43328_);
  or (_00386_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00387_, _00386_, _43821_);
  and (_00388_, _00387_, _00385_);
  or (_39286_, _00388_, _00382_);
  and (_00389_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00390_, _43789_, _43441_);
  nor (_00391_, _00390_, _43790_);
  or (_00392_, _00391_, _43328_);
  or (_00393_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00394_, _00393_, _43821_);
  and (_00395_, _00394_, _00392_);
  or (_39287_, _00395_, _00389_);
  and (_00396_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00397_, _43794_, _43790_);
  nor (_00398_, _00397_, _43795_);
  or (_00399_, _00398_, _43328_);
  or (_00400_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00401_, _00400_, _43821_);
  and (_00402_, _00401_, _00399_);
  or (_39288_, _00402_, _00396_);
  and (_00403_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00404_, _43795_, _43434_);
  nor (_00405_, _00404_, _43797_);
  or (_00406_, _00405_, _43328_);
  or (_00407_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_00408_, _00407_, _43821_);
  and (_00409_, _00408_, _00406_);
  or (_39289_, _00409_, _00403_);
  nor (_00410_, _43797_, _43428_);
  nor (_00411_, _00410_, _43798_);
  or (_00412_, _00411_, _43328_);
  or (_00413_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00414_, _00413_, _43821_);
  and (_00415_, _00414_, _00412_);
  and (_00416_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39290_, _00416_, _00415_);
  and (_00417_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00418_, _43798_, _43424_);
  nor (_00419_, _00418_, _43799_);
  or (_00420_, _00419_, _43328_);
  or (_00421_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_00422_, _00421_, _43821_);
  and (_00423_, _00422_, _00420_);
  or (_39291_, _00423_, _00417_);
  nor (_00424_, _43802_, _43799_);
  nor (_00425_, _00424_, _43803_);
  or (_00426_, _00425_, _43328_);
  or (_00427_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00428_, _00427_, _43821_);
  and (_00429_, _00428_, _00426_);
  and (_00430_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_39292_, _00430_, _00429_);
  nor (_00431_, _43803_, _43418_);
  nor (_00432_, _00431_, _43805_);
  or (_00433_, _00432_, _43328_);
  or (_00434_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00435_, _00434_, _43821_);
  and (_00436_, _00435_, _00433_);
  and (_00437_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39293_, _00437_, _00436_);
  nor (_00438_, _43805_, _43409_);
  nor (_00439_, _00438_, _43806_);
  or (_00440_, _00439_, _43328_);
  or (_00441_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00442_, _00441_, _43821_);
  and (_00443_, _00442_, _00440_);
  and (_00444_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_39294_, _00444_, _00443_);
  nor (_00445_, _43806_, _43406_);
  nor (_00446_, _00445_, _43807_);
  or (_00447_, _00446_, _43328_);
  or (_00448_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00449_, _00448_, _43821_);
  and (_00450_, _00449_, _00447_);
  and (_00451_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39296_, _00451_, _00450_);
  nor (_00452_, _43807_, _43399_);
  nor (_00453_, _00452_, _43809_);
  or (_00454_, _00453_, _43328_);
  or (_00455_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00456_, _00455_, _43821_);
  and (_00457_, _00456_, _00454_);
  and (_00458_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_39297_, _00458_, _00457_);
  nor (_00459_, _43809_, _43393_);
  nor (_00460_, _00459_, _43810_);
  or (_00461_, _00460_, _43328_);
  or (_00462_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00463_, _00462_, _43821_);
  and (_00464_, _00463_, _00461_);
  and (_00465_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_39298_, _00465_, _00464_);
  nor (_00466_, _43810_, _43387_);
  nor (_00467_, _00466_, _43811_);
  or (_00468_, _00467_, _43328_);
  or (_00469_, _43327_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00470_, _00469_, _43821_);
  and (_00471_, _00470_, _00468_);
  and (_00472_, _43323_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_39299_, _00472_, _00471_);
  and (_00473_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_00474_, _00473_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39300_, _00474_, _41806_);
  and (_00475_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_00476_, _00475_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39301_, _00476_, _41806_);
  and (_00477_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_00478_, _00477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39302_, _00478_, _41806_);
  and (_00479_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_00480_, _00479_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39303_, _00480_, _41806_);
  and (_00481_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_00482_, _00481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39304_, _00482_, _41806_);
  and (_00483_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_00484_, _00483_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39305_, _00484_, _41806_);
  and (_00485_, _43835_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_00486_, _00485_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39307_, _00486_, _41806_);
  nor (_00487_, _43773_, _40305_);
  nand (_00488_, _00487_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00489_, _00487_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00490_, _00489_, _43821_);
  and (_39308_, _00490_, _00488_);
  nor (_00491_, _43850_, _43848_);
  nor (_00492_, _00491_, _43851_);
  or (_00493_, _00492_, _40305_);
  or (_00494_, _33860_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00495_, _00494_, _43821_);
  and (_39309_, _00495_, _00493_);
  and (_00496_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_00497_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_00498_, _00497_, _38935_);
  or (_39324_, _00498_, _00496_);
  and (_00499_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00500_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00501_, _00500_, _38935_);
  or (_39325_, _00501_, _00499_);
  and (_00502_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00503_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00504_, _00503_, _38935_);
  or (_39326_, _00504_, _00502_);
  and (_00505_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00506_, _44034_, _38935_);
  or (_39328_, _00506_, _00505_);
  and (_00507_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00508_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_00509_, _00508_, _38935_);
  or (_39329_, _00509_, _00507_);
  and (_00510_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00511_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_00512_, _00511_, _38935_);
  or (_39330_, _00512_, _00510_);
  and (_00513_, _43874_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00514_, _44044_, _38935_);
  or (_39331_, _00514_, _00513_);
  and (_39332_, _43882_, _41806_);
  nor (_39333_, _43892_, rst);
  and (_39334_, _43888_, _41806_);
  and (_00515_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00516_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00517_, _00516_, _00515_);
  and (_39335_, _00517_, _41806_);
  and (_00518_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00519_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00520_, _00519_, _00518_);
  and (_39336_, _00520_, _41806_);
  and (_00521_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00522_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00523_, _00522_, _00521_);
  and (_39337_, _00523_, _41806_);
  and (_00524_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00525_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00526_, _00525_, _00524_);
  and (_39339_, _00526_, _41806_);
  and (_00527_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00528_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00529_, _00528_, _00527_);
  and (_39340_, _00529_, _41806_);
  and (_00530_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00531_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00532_, _00531_, _00530_);
  and (_39341_, _00532_, _41806_);
  and (_00533_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00534_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00535_, _00534_, _00533_);
  and (_39342_, _00535_, _41806_);
  and (_00536_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00537_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00538_, _00537_, _00536_);
  and (_39343_, _00538_, _41806_);
  and (_00539_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00540_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00541_, _00540_, _00539_);
  and (_39344_, _00541_, _41806_);
  and (_00542_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00543_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00544_, _00543_, _00542_);
  and (_39345_, _00544_, _41806_);
  and (_00545_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00546_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00547_, _00546_, _00545_);
  and (_39346_, _00547_, _41806_);
  and (_00548_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00549_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00550_, _00549_, _00548_);
  and (_39347_, _00550_, _41806_);
  and (_00551_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00552_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00553_, _00552_, _00551_);
  and (_39348_, _00553_, _41806_);
  and (_00554_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00555_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00556_, _00555_, _00554_);
  and (_39350_, _00556_, _41806_);
  and (_00557_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00558_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00559_, _00558_, _00557_);
  and (_39351_, _00559_, _41806_);
  and (_00560_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00561_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00562_, _00561_, _00560_);
  and (_39352_, _00562_, _41806_);
  and (_00563_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00564_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00565_, _00564_, _00563_);
  and (_39353_, _00565_, _41806_);
  and (_00566_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00567_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00568_, _00567_, _00566_);
  and (_39354_, _00568_, _41806_);
  and (_00569_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00570_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00571_, _00570_, _00569_);
  and (_39355_, _00571_, _41806_);
  and (_00572_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00573_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00574_, _00573_, _00572_);
  and (_39356_, _00574_, _41806_);
  and (_00575_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00576_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00577_, _00576_, _00575_);
  and (_39357_, _00577_, _41806_);
  and (_00578_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00579_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00580_, _00579_, _00578_);
  and (_39358_, _00580_, _41806_);
  and (_00581_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00582_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00583_, _00582_, _00581_);
  and (_39359_, _00583_, _41806_);
  and (_00584_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00585_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00586_, _00585_, _00584_);
  and (_39361_, _00586_, _41806_);
  and (_00587_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00588_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00589_, _00588_, _00587_);
  and (_39362_, _00589_, _41806_);
  and (_00590_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00591_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00592_, _00591_, _00590_);
  and (_39363_, _00592_, _41806_);
  and (_00593_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00594_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00595_, _00594_, _00593_);
  and (_39364_, _00595_, _41806_);
  and (_00596_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00597_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00598_, _00597_, _00596_);
  and (_39365_, _00598_, _41806_);
  and (_00599_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00600_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00601_, _00600_, _00599_);
  and (_39366_, _00601_, _41806_);
  and (_00602_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00603_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00604_, _00603_, _00602_);
  and (_39367_, _00604_, _41806_);
  and (_00605_, _43896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00606_, _43898_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00607_, _00606_, _00605_);
  and (_39368_, _00607_, _41806_);
  and (_00608_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00609_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00610_, _00609_, _00608_);
  and (_39369_, _00610_, _41806_);
  and (_00611_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00612_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00613_, _00612_, _00611_);
  and (_39370_, _00613_, _41806_);
  and (_00614_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00615_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00616_, _00615_, _00614_);
  and (_39372_, _00616_, _41806_);
  and (_00617_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00618_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00619_, _00618_, _00617_);
  and (_39373_, _00619_, _41806_);
  and (_00620_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00621_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00622_, _00621_, _00620_);
  and (_39374_, _00622_, _41806_);
  and (_00623_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00624_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00625_, _00624_, _00623_);
  and (_39375_, _00625_, _41806_);
  and (_00626_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00627_, _43906_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00628_, _00627_, _00626_);
  and (_39376_, _00628_, _41806_);
  and (_00629_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00630_, _40408_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00631_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00632_, _00631_, _43905_);
  and (_00633_, _00632_, _00630_);
  or (_00634_, _00633_, _00629_);
  and (_39377_, _00634_, _41806_);
  and (_00635_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00636_, _40564_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00637_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00638_, _00637_, _43905_);
  and (_00639_, _00638_, _00636_);
  or (_00640_, _00639_, _00635_);
  and (_39378_, _00640_, _41806_);
  and (_00641_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00642_, _40492_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00643_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00644_, _00643_, _43905_);
  and (_00645_, _00644_, _00642_);
  or (_00646_, _00645_, _00641_);
  and (_39379_, _00646_, _41806_);
  and (_00647_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00648_, _40370_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00649_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00650_, _00649_, _43905_);
  and (_00651_, _00650_, _00648_);
  or (_00652_, _00651_, _00647_);
  and (_39380_, _00652_, _41806_);
  and (_00653_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00654_, _40540_, _43912_);
  or (_00655_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00656_, _00655_, _43905_);
  and (_00657_, _00656_, _00654_);
  or (_00658_, _00657_, _00653_);
  and (_39381_, _00658_, _41806_);
  and (_00659_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00660_, _40442_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00661_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00662_, _00661_, _43905_);
  and (_00663_, _00662_, _00660_);
  or (_00664_, _00663_, _00659_);
  and (_39383_, _00664_, _41806_);
  and (_00665_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00666_, _40639_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00667_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00668_, _00667_, _43905_);
  and (_00669_, _00668_, _00666_);
  or (_00670_, _00669_, _00665_);
  and (_39384_, _00670_, _41806_);
  and (_00671_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00672_, _40300_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00673_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00674_, _00673_, _43905_);
  and (_00675_, _00674_, _00672_);
  or (_00676_, _00675_, _00671_);
  and (_39385_, _00676_, _41806_);
  and (_00677_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00678_, _00677_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00679_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _43905_);
  and (_00680_, _00679_, _41806_);
  and (_39386_, _00680_, _00678_);
  and (_00681_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00682_, _00681_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00683_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _43905_);
  and (_00684_, _00683_, _41806_);
  and (_39387_, _00684_, _00682_);
  and (_00685_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00686_, _00685_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00687_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _43905_);
  and (_00688_, _00687_, _41806_);
  and (_39388_, _00688_, _00686_);
  and (_00689_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00690_, _00689_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00691_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _43905_);
  and (_00692_, _00691_, _41806_);
  and (_39389_, _00692_, _00690_);
  and (_00693_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00694_, _00693_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00695_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _43905_);
  and (_00696_, _00695_, _41806_);
  and (_39390_, _00696_, _00694_);
  and (_00697_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_00698_, _00697_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00699_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _43905_);
  and (_00700_, _00699_, _41806_);
  and (_39391_, _00700_, _00698_);
  and (_00701_, _43912_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_00702_, _00701_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00703_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _43905_);
  and (_00704_, _00703_, _41806_);
  and (_39392_, _00704_, _00702_);
  nand (_00705_, _43919_, _29231_);
  or (_00706_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00707_, _00706_, _41806_);
  and (_39394_, _00707_, _00705_);
  nand (_00708_, _43919_, _29893_);
  or (_00709_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00710_, _00709_, _41806_);
  and (_39395_, _00710_, _00708_);
  nand (_00711_, _43919_, _30567_);
  or (_00712_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00713_, _00712_, _41806_);
  and (_39396_, _00713_, _00711_);
  nand (_00714_, _43919_, _31338_);
  or (_00715_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00716_, _00715_, _41806_);
  and (_39397_, _00716_, _00714_);
  nand (_00717_, _43919_, _32044_);
  or (_00718_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00719_, _00718_, _41806_);
  and (_39398_, _00719_, _00717_);
  nand (_00720_, _43919_, _32853_);
  or (_00721_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00722_, _00721_, _41806_);
  and (_39399_, _00722_, _00720_);
  nand (_00723_, _43919_, _33598_);
  or (_00724_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00725_, _00724_, _41806_);
  and (_39400_, _00725_, _00723_);
  nand (_00726_, _43919_, _28011_);
  or (_00727_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00728_, _00727_, _41806_);
  and (_39401_, _00728_, _00726_);
  nand (_00729_, _43919_, _38617_);
  or (_00730_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00731_, _00730_, _41806_);
  and (_39402_, _00731_, _00729_);
  nand (_00732_, _43919_, _38645_);
  or (_00733_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00734_, _00733_, _41806_);
  and (_39403_, _00734_, _00732_);
  nand (_00735_, _43919_, _38673_);
  or (_00736_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00737_, _00736_, _41806_);
  and (_39405_, _00737_, _00735_);
  nand (_00738_, _43919_, _38702_);
  or (_00739_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00740_, _00739_, _41806_);
  and (_39406_, _00740_, _00738_);
  nand (_00741_, _43919_, _38731_);
  or (_00742_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00743_, _00742_, _41806_);
  and (_39407_, _00743_, _00741_);
  nand (_00744_, _43919_, _38760_);
  or (_00745_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00746_, _00745_, _41806_);
  and (_39408_, _00746_, _00744_);
  nand (_00747_, _43919_, _38787_);
  or (_00748_, _43919_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00749_, _00748_, _41806_);
  and (_39409_, _00749_, _00747_);
  nor (_39617_, _40339_, rst);
  nor (_00750_, _40703_, _40463_);
  nor (_00751_, _40547_, _40327_);
  and (_00752_, _00751_, _40380_);
  and (_00753_, _00752_, _00750_);
  not (_00754_, _00753_);
  nor (_00755_, _00754_, _39024_);
  and (_00756_, _40380_, _40547_);
  and (_00757_, _00756_, _40463_);
  nor (_00758_, _40703_, _40327_);
  and (_00759_, _00758_, _00757_);
  not (_00760_, _40500_);
  nor (_00761_, _39128_, _39116_);
  and (_00762_, _39128_, _39116_);
  nor (_00763_, _00762_, _00761_);
  nor (_00764_, _39140_, _39048_);
  and (_00765_, _39140_, _39048_);
  nor (_00766_, _00765_, _00764_);
  and (_00767_, _00766_, _00763_);
  nor (_00768_, _00766_, _00763_);
  or (_00769_, _00768_, _00767_);
  and (_00770_, _39073_, _39060_);
  nor (_00771_, _39073_, _39060_);
  or (_00772_, _00771_, _00770_);
  not (_00773_, _00772_);
  nor (_00774_, _39104_, _39093_);
  and (_00775_, _39104_, _39093_);
  or (_00776_, _00775_, _00774_);
  and (_00777_, _00776_, _00773_);
  nor (_00778_, _00776_, _00773_);
  nor (_00779_, _00778_, _00777_);
  nor (_00780_, _00779_, _00769_);
  and (_00781_, _00779_, _00769_);
  nor (_00782_, _00781_, _00780_);
  nor (_00783_, _00782_, _00760_);
  and (_00784_, _40415_, _40611_);
  nand (_00785_, _00760_, _38964_);
  nand (_00786_, _00785_, _00784_);
  or (_00787_, _00786_, _00783_);
  not (_00788_, _40415_);
  and (_00789_, _00788_, _40611_);
  not (_00790_, _00789_);
  and (_00791_, _00760_, _38971_);
  and (_00792_, _40500_, _38870_);
  nor (_00793_, _00792_, _00791_);
  or (_00794_, _00793_, _00790_);
  nor (_00795_, _40415_, _40611_);
  not (_00796_, _00795_);
  and (_00797_, _00760_, _38862_);
  and (_00798_, _40500_, _38933_);
  or (_00799_, _00798_, _00797_);
  or (_00800_, _00799_, _00796_);
  and (_00801_, _00800_, _00794_);
  nor (_00802_, _00760_, _38907_);
  nor (_00803_, _00788_, _40611_);
  nand (_00804_, _00760_, _39004_);
  nand (_00805_, _00804_, _00803_);
  or (_00806_, _00805_, _00802_);
  and (_00807_, _00806_, _00801_);
  nand (_00808_, _00807_, _00787_);
  and (_00809_, _00808_, _00759_);
  and (_00810_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_00811_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_00812_, _00811_, _00810_);
  and (_00813_, _00812_, _00803_);
  or (_00814_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_00815_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_00816_, _00815_, _00789_);
  and (_00817_, _00816_, _00814_);
  and (_00818_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_00819_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_00820_, _00819_, _00818_);
  and (_00821_, _00820_, _00795_);
  nand (_00822_, _40500_, _39870_);
  or (_00823_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_00824_, _00823_, _00784_);
  and (_00825_, _00824_, _00822_);
  or (_00826_, _00825_, _00821_);
  or (_00827_, _00826_, _00817_);
  or (_00828_, _00827_, _00813_);
  and (_00829_, _40703_, _40463_);
  and (_00830_, _00751_, _40381_);
  and (_00831_, _00830_, _00829_);
  and (_00832_, _00831_, _00828_);
  and (_00833_, _40703_, _40464_);
  and (_00834_, _00830_, _00833_);
  and (_00835_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_00836_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00837_, _00836_, _00835_);
  and (_00838_, _00837_, _00803_);
  or (_00839_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_00840_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_00841_, _00840_, _00789_);
  and (_00842_, _00841_, _00839_);
  nor (_00843_, _40500_, _39908_);
  and (_00844_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_00845_, _00844_, _00843_);
  and (_00846_, _00845_, _00795_);
  or (_00847_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_00848_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_00849_, _00848_, _00784_);
  and (_00850_, _00849_, _00847_);
  or (_00851_, _00850_, _00846_);
  or (_00852_, _00851_, _00842_);
  or (_00853_, _00852_, _00838_);
  and (_00854_, _00853_, _00834_);
  nor (_00855_, _00854_, _00832_);
  nor (_00856_, _42622_, _37475_);
  and (_00857_, _36069_, _37646_);
  or (_00858_, _00857_, _37095_);
  nor (_00859_, _00858_, _35839_);
  and (_00860_, _42461_, _35915_);
  and (_00861_, _34793_, _42458_);
  or (_00863_, _00861_, _00860_);
  or (_00864_, _00863_, _42524_);
  nor (_00865_, _00864_, _37133_);
  and (_00866_, _00865_, _00859_);
  nor (_00867_, _42457_, _37056_);
  and (_00868_, _00867_, _42526_);
  and (_00869_, _00868_, _00866_);
  and (_00870_, _00869_, _37373_);
  and (_00871_, _00870_, _00856_);
  nor (_00872_, _00871_, _33817_);
  and (_00873_, _43004_, p2in_reg[2]);
  and (_00874_, _43000_, p2_in[2]);
  nor (_00875_, _00874_, _00873_);
  nor (_00876_, _00875_, _00872_);
  and (_00877_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_00878_, _00877_, _00876_);
  nor (_00879_, _00878_, _00760_);
  and (_00880_, _43004_, p2in_reg[6]);
  and (_00881_, _43000_, p2_in[6]);
  nor (_00882_, _00881_, _00880_);
  nor (_00883_, _00882_, _00872_);
  and (_00884_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_00885_, _00884_, _00883_);
  or (_00886_, _00885_, _40500_);
  nand (_00887_, _00886_, _00803_);
  or (_00888_, _00887_, _00879_);
  not (_00889_, _00784_);
  and (_00890_, _43004_, p2in_reg[4]);
  and (_00891_, _43000_, p2_in[4]);
  nor (_00892_, _00891_, _00890_);
  nor (_00894_, _00892_, _00872_);
  and (_00895_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_00896_, _00895_, _00894_);
  nand (_00897_, _00896_, _00760_);
  and (_00898_, _43004_, p2in_reg[0]);
  and (_00899_, _43000_, p2_in[0]);
  nor (_00900_, _00899_, _00898_);
  nor (_00901_, _00900_, _00872_);
  and (_00902_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_00903_, _00902_, _00901_);
  nand (_00904_, _00903_, _40500_);
  and (_00905_, _00904_, _00897_);
  or (_00906_, _00905_, _00889_);
  and (_00907_, _43004_, p2in_reg[7]);
  and (_00908_, _43000_, p2_in[7]);
  nor (_00909_, _00908_, _00907_);
  nor (_00910_, _00909_, _00872_);
  and (_00911_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_00912_, _00911_, _00910_);
  nand (_00913_, _00912_, _00760_);
  and (_00915_, _43004_, p2in_reg[3]);
  and (_00916_, _43000_, p2_in[3]);
  nor (_00917_, _00916_, _00915_);
  nor (_00918_, _00917_, _00872_);
  and (_00919_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_00920_, _00919_, _00918_);
  nand (_00921_, _00920_, _40500_);
  and (_00922_, _00921_, _00913_);
  or (_00923_, _00922_, _00796_);
  and (_00924_, _00923_, _00906_);
  and (_00925_, _43004_, p2in_reg[1]);
  and (_00926_, _43000_, p2_in[1]);
  nor (_00927_, _00926_, _00925_);
  nor (_00928_, _00927_, _00872_);
  and (_00929_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_00930_, _00929_, _00928_);
  nor (_00931_, _00930_, _00760_);
  and (_00932_, _43004_, p2in_reg[5]);
  and (_00933_, _43000_, p2_in[5]);
  nor (_00934_, _00933_, _00932_);
  nor (_00935_, _00934_, _00872_);
  and (_00936_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_00937_, _00936_, _00935_);
  or (_00938_, _00937_, _40500_);
  nand (_00939_, _00938_, _00789_);
  or (_00940_, _00939_, _00931_);
  and (_00941_, _00940_, _00924_);
  and (_00942_, _00941_, _00888_);
  nand (_00943_, _00833_, _00752_);
  or (_00944_, _00943_, _00942_);
  and (_00945_, _00944_, _00855_);
  not (_00946_, _40327_);
  and (_00947_, _00756_, _00946_);
  and (_00948_, _00947_, _00750_);
  nand (_00949_, _40500_, _29264_);
  or (_00950_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_00951_, _00950_, _00784_);
  and (_00952_, _00951_, _00949_);
  nor (_00953_, _40500_, _28098_);
  and (_00954_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00955_, _00954_, _00953_);
  and (_00956_, _00955_, _00795_);
  nor (_00957_, _40500_, _33631_);
  and (_00958_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00959_, _00958_, _00957_);
  and (_00960_, _00959_, _00803_);
  nand (_00961_, _40500_, _29926_);
  or (_00962_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_00963_, _00962_, _00789_);
  and (_00964_, _00963_, _00961_);
  or (_00965_, _00964_, _00960_);
  or (_00966_, _00965_, _00956_);
  or (_00967_, _00966_, _00952_);
  and (_00968_, _00967_, _00948_);
  nor (_00969_, _40380_, _40327_);
  and (_00970_, _40703_, _40547_);
  and (_00971_, _00970_, _00969_);
  and (_00972_, _00971_, _40464_);
  nand (_00973_, _40500_, _39920_);
  or (_00974_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_00975_, _00974_, _00784_);
  and (_00976_, _00975_, _00973_);
  and (_00977_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_00978_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_00979_, _00978_, _00977_);
  and (_00980_, _00979_, _00795_);
  and (_00981_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_00982_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_00983_, _00982_, _00981_);
  and (_00984_, _00983_, _00803_);
  nand (_00985_, _40500_, _39922_);
  or (_00986_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_00987_, _00986_, _00789_);
  and (_00988_, _00987_, _00985_);
  or (_00989_, _00988_, _00984_);
  or (_00990_, _00989_, _00980_);
  or (_00991_, _00990_, _00976_);
  and (_00992_, _00991_, _00972_);
  nor (_00993_, _00992_, _00968_);
  nand (_00994_, _00947_, _00833_);
  and (_00995_, _43004_, p3in_reg[2]);
  and (_00996_, _43000_, p3_in[2]);
  nor (_00997_, _00996_, _00995_);
  nor (_00998_, _00997_, _00872_);
  and (_00999_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_01000_, _00999_, _00998_);
  nor (_01001_, _01000_, _00760_);
  and (_01002_, _43004_, p3in_reg[6]);
  and (_01003_, _43000_, p3_in[6]);
  nor (_01004_, _01003_, _01002_);
  nor (_01005_, _01004_, _00872_);
  and (_01006_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_01007_, _01006_, _01005_);
  or (_01008_, _01007_, _40500_);
  nand (_01009_, _01008_, _00803_);
  or (_01010_, _01009_, _01001_);
  and (_01011_, _43004_, p3in_reg[4]);
  and (_01012_, _43000_, p3_in[4]);
  nor (_01013_, _01012_, _01011_);
  nor (_01014_, _01013_, _00872_);
  and (_01015_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_01016_, _01015_, _01014_);
  nand (_01017_, _01016_, _00760_);
  and (_01018_, _43004_, p3in_reg[0]);
  and (_01019_, _43000_, p3_in[0]);
  nor (_01020_, _01019_, _01018_);
  nor (_01021_, _01020_, _00872_);
  and (_01022_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_01023_, _01022_, _01021_);
  nand (_01024_, _01023_, _40500_);
  and (_01025_, _01024_, _01017_);
  or (_01026_, _01025_, _00889_);
  and (_01027_, _43004_, p3in_reg[7]);
  and (_01028_, _43000_, p3_in[7]);
  nor (_01029_, _01028_, _01027_);
  nor (_01030_, _01029_, _00872_);
  and (_01031_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_01032_, _01031_, _01030_);
  nand (_01033_, _01032_, _00760_);
  and (_01034_, _43004_, p3in_reg[3]);
  and (_01035_, _43000_, p3_in[3]);
  nor (_01036_, _01035_, _01034_);
  nor (_01037_, _01036_, _00872_);
  and (_01038_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_01039_, _01038_, _01037_);
  nand (_01040_, _01039_, _40500_);
  and (_01041_, _01040_, _01033_);
  or (_01042_, _01041_, _00796_);
  and (_01043_, _01042_, _01026_);
  and (_01044_, _43004_, p3in_reg[1]);
  and (_01045_, _43000_, p3_in[1]);
  nor (_01046_, _01045_, _01044_);
  nor (_01047_, _01046_, _00872_);
  and (_01048_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_01049_, _01048_, _01047_);
  nor (_01050_, _01049_, _00760_);
  and (_01051_, _43004_, p3in_reg[5]);
  and (_01052_, _43000_, p3_in[5]);
  nor (_01053_, _01052_, _01051_);
  nor (_01054_, _01053_, _00872_);
  and (_01055_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_01056_, _01055_, _01054_);
  or (_01057_, _01056_, _40500_);
  nand (_01058_, _01057_, _00789_);
  or (_01059_, _01058_, _01050_);
  and (_01060_, _01059_, _01043_);
  and (_01061_, _01060_, _01010_);
  or (_01062_, _01061_, _00994_);
  and (_01063_, _01062_, _00993_);
  and (_01064_, _00830_, _40703_);
  or (_01065_, _01064_, _00948_);
  nor (_01066_, _01065_, _00759_);
  nor (_01067_, _40381_, _40327_);
  and (_01068_, _01067_, _40703_);
  nor (_01069_, _01068_, _00971_);
  and (_01070_, _01069_, _00754_);
  and (_01071_, _01070_, _01066_);
  nand (_01072_, _43104_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_01073_, _01072_, _01071_);
  nand (_01074_, _00947_, _00829_);
  and (_01075_, _43004_, p1in_reg[5]);
  and (_01076_, _43000_, p1_in[5]);
  nor (_01077_, _01076_, _01075_);
  nor (_01078_, _01077_, _00872_);
  and (_01079_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_01080_, _01079_, _01078_);
  nand (_01081_, _01080_, _00760_);
  and (_01082_, _43004_, p1in_reg[1]);
  and (_01083_, _43000_, p1_in[1]);
  nor (_01084_, _01083_, _01082_);
  nor (_01085_, _01084_, _00872_);
  and (_01086_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_01087_, _01086_, _01085_);
  nand (_01088_, _01087_, _40500_);
  and (_01089_, _01088_, _01081_);
  or (_01090_, _01089_, _00790_);
  and (_01091_, _43004_, p1in_reg[7]);
  and (_01092_, _43000_, p1_in[7]);
  nor (_01093_, _01092_, _01091_);
  nor (_01094_, _01093_, _00872_);
  and (_01095_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_01096_, _01095_, _01094_);
  nand (_01097_, _01096_, _00760_);
  and (_01098_, _43004_, p1in_reg[3]);
  and (_01099_, _43000_, p1_in[3]);
  nor (_01100_, _01099_, _01098_);
  nor (_01101_, _01100_, _00872_);
  and (_01102_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_01103_, _01102_, _01101_);
  nand (_01104_, _01103_, _40500_);
  and (_01105_, _01104_, _01097_);
  or (_01106_, _01105_, _00796_);
  and (_01107_, _01106_, _01090_);
  not (_01108_, _00803_);
  and (_01109_, _43004_, p1in_reg[6]);
  and (_01110_, _43000_, p1_in[6]);
  nor (_01111_, _01110_, _01109_);
  nor (_01112_, _01111_, _00872_);
  and (_01113_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_01114_, _01113_, _01112_);
  nand (_01115_, _01114_, _00760_);
  and (_01116_, _43004_, p1in_reg[2]);
  and (_01117_, _43000_, p1_in[2]);
  nor (_01118_, _01117_, _01116_);
  nor (_01119_, _01118_, _00872_);
  and (_01120_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_01121_, _01120_, _01119_);
  nand (_01122_, _01121_, _40500_);
  and (_01123_, _01122_, _01115_);
  or (_01124_, _01123_, _01108_);
  and (_01125_, _43004_, p1in_reg[4]);
  and (_01126_, _43000_, p1_in[4]);
  nor (_01127_, _01126_, _01125_);
  nor (_01128_, _01127_, _00872_);
  and (_01129_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_01130_, _01129_, _01128_);
  nand (_01131_, _01130_, _00760_);
  and (_01132_, _43004_, p1in_reg[0]);
  and (_01133_, _43000_, p1_in[0]);
  nor (_01134_, _01133_, _01132_);
  nor (_01135_, _01134_, _00872_);
  and (_01136_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_01137_, _01136_, _01135_);
  nand (_01138_, _01137_, _40500_);
  and (_01139_, _01138_, _01131_);
  or (_01140_, _01139_, _00889_);
  and (_01141_, _01140_, _01124_);
  and (_01142_, _01141_, _01107_);
  or (_01143_, _01142_, _01074_);
  and (_01144_, _00829_, _00752_);
  and (_01145_, _43004_, p0in_reg[5]);
  and (_01146_, _43000_, p0_in[5]);
  nor (_01147_, _01146_, _01145_);
  nor (_01148_, _01147_, _00872_);
  and (_01149_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_01150_, _01149_, _01148_);
  nand (_01151_, _01150_, _00760_);
  and (_01152_, _43004_, p0in_reg[1]);
  and (_01153_, _43000_, p0_in[1]);
  nor (_01154_, _01153_, _01152_);
  nor (_01155_, _01154_, _00872_);
  and (_01156_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_01157_, _01156_, _01155_);
  nand (_01158_, _01157_, _40500_);
  and (_01159_, _01158_, _01151_);
  or (_01160_, _01159_, _00790_);
  and (_01161_, _43004_, p0in_reg[4]);
  and (_01162_, _43000_, p0_in[4]);
  nor (_01163_, _01162_, _01161_);
  nor (_01164_, _01163_, _00872_);
  and (_01165_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_01166_, _01165_, _01164_);
  nand (_01167_, _01166_, _00760_);
  and (_01168_, _43004_, p0in_reg[0]);
  and (_01169_, _43000_, p0_in[0]);
  nor (_01170_, _01169_, _01168_);
  nor (_01171_, _01170_, _00872_);
  and (_01172_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_01173_, _01172_, _01171_);
  nand (_01174_, _01173_, _40500_);
  and (_01175_, _01174_, _01167_);
  or (_01176_, _01175_, _00889_);
  and (_01177_, _01176_, _01160_);
  and (_01178_, _43004_, p0in_reg[6]);
  and (_01179_, _43000_, p0_in[6]);
  nor (_01180_, _01179_, _01178_);
  nor (_01181_, _01180_, _00872_);
  and (_01182_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_01183_, _01182_, _01181_);
  nand (_01184_, _01183_, _00760_);
  and (_01185_, _43004_, p0in_reg[2]);
  and (_01186_, _43000_, p0_in[2]);
  nor (_01187_, _01186_, _01185_);
  nor (_01188_, _01187_, _00872_);
  and (_01189_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_01190_, _01189_, _01188_);
  nand (_01191_, _01190_, _40500_);
  and (_01192_, _01191_, _01184_);
  or (_01193_, _01192_, _01108_);
  and (_01194_, _43004_, p0in_reg[7]);
  and (_01195_, _43000_, p0_in[7]);
  nor (_01196_, _01195_, _01194_);
  nor (_01197_, _01196_, _00872_);
  and (_01198_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_01199_, _01198_, _01197_);
  nand (_01200_, _01199_, _00760_);
  and (_01201_, _43004_, p0in_reg[3]);
  and (_01202_, _43000_, p0_in[3]);
  nor (_01203_, _01202_, _01201_);
  nor (_01204_, _01203_, _00872_);
  and (_01205_, _00872_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_01206_, _01205_, _01204_);
  nand (_01207_, _01206_, _40500_);
  and (_01208_, _01207_, _01200_);
  or (_01209_, _01208_, _00796_);
  and (_01210_, _01209_, _01193_);
  nand (_01211_, _01210_, _01177_);
  nand (_01212_, _01211_, _01144_);
  and (_01213_, _01212_, _01143_);
  and (_01214_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01215_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_01216_, _01215_, _01214_);
  and (_01217_, _01216_, _00784_);
  or (_01218_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_01219_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01220_, _01219_, _00795_);
  and (_01221_, _01220_, _01218_);
  and (_01222_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01223_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_01224_, _01223_, _01222_);
  and (_01225_, _01224_, _00789_);
  nand (_01226_, _40500_, _39082_);
  or (_01227_, _40500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01228_, _01227_, _00803_);
  and (_01229_, _01228_, _01226_);
  or (_01230_, _01229_, _01225_);
  or (_01231_, _01230_, _01221_);
  or (_01232_, _01231_, _01217_);
  nand (_01233_, _01232_, _00753_);
  and (_01234_, _01233_, _01213_);
  and (_01235_, _01234_, _01073_);
  and (_01236_, _01235_, _01063_);
  nand (_01237_, _01236_, _00945_);
  or (_01238_, _01237_, _00809_);
  or (_01239_, _01073_, _29318_);
  and (_01240_, _01239_, _01238_);
  or (_01241_, _01240_, _00755_);
  and (_01242_, _00789_, _39073_);
  and (_01243_, _00784_, _39060_);
  or (_01244_, _01243_, _01242_);
  nor (_01245_, _00796_, _39104_);
  nor (_01246_, _01108_, _39093_);
  or (_01247_, _01246_, _01245_);
  or (_01248_, _01247_, _01244_);
  and (_01249_, _01248_, _40500_);
  and (_01250_, _00789_, _39128_);
  and (_01251_, _00795_, _39048_);
  or (_01252_, _01251_, _01250_);
  and (_01253_, _00784_, _39116_);
  and (_01254_, _00803_, _39140_);
  or (_01255_, _01254_, _01253_);
  or (_01256_, _01255_, _01252_);
  nand (_01257_, _01256_, _00760_);
  nand (_01258_, _01257_, _00755_);
  or (_01259_, _01258_, _01249_);
  and (_01260_, _01259_, _01241_);
  not (_01261_, _38817_);
  not (_01262_, _00872_);
  and (_01263_, _01068_, _01262_);
  nor (_01264_, _01263_, _01261_);
  and (_01265_, _01264_, _43027_);
  not (_01266_, _01265_);
  nor (_01267_, _01266_, _01071_);
  or (_01268_, _01267_, _01260_);
  and (_01269_, _00803_, _40633_);
  and (_01270_, _00784_, _40538_);
  or (_01271_, _01270_, _40500_);
  or (_01272_, _01271_, _01269_);
  and (_01273_, _00803_, _40482_);
  and (_01274_, _00784_, _38426_);
  or (_01275_, _01274_, _00760_);
  or (_01276_, _01275_, _01273_);
  and (_01277_, _01276_, _01272_);
  and (_01278_, _40500_, _38418_);
  nor (_01279_, _40500_, _38366_);
  or (_01280_, _01279_, _01278_);
  and (_01281_, _01280_, _00789_);
  and (_01282_, _40500_, _40360_);
  nor (_01283_, _40500_, _38162_);
  or (_01284_, _01283_, _01282_);
  and (_01285_, _01284_, _00795_);
  or (_01286_, _01285_, _01281_);
  nor (_01287_, _01286_, _01277_);
  nand (_01288_, _01287_, _01267_);
  and (_01289_, _01288_, _41806_);
  and (_39648_, _01289_, _01268_);
  and (_01290_, _40547_, _40463_);
  and (_01291_, _40380_, _40500_);
  and (_01292_, _01291_, _00784_);
  and (_01293_, _01292_, _01290_);
  and (_01294_, _01293_, _00758_);
  and (_01295_, _01294_, _38823_);
  and (_01296_, _00829_, _00751_);
  and (_01297_, _01291_, _00795_);
  and (_01298_, _01297_, _01296_);
  and (_01299_, _01298_, _38493_);
  nor (_01300_, _01299_, _01295_);
  nor (_01301_, _01300_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_01302_, _01301_);
  nand (_01303_, _39024_, _39022_);
  and (_01304_, _00784_, _40500_);
  and (_01305_, _01304_, _00753_);
  and (_01306_, _01305_, _01303_);
  and (_01307_, _00795_, _00760_);
  nor (_01308_, _01307_, _38954_);
  and (_01309_, _01308_, _43027_);
  nor (_01310_, _01309_, _01306_);
  and (_01311_, _01310_, _43107_);
  and (_01312_, _01311_, _01302_);
  and (_01313_, _01291_, _00803_);
  and (_01314_, _01313_, _01296_);
  and (_01315_, _01314_, _38493_);
  or (_01316_, _01315_, rst);
  nor (_39649_, _01316_, _01312_);
  not (_01317_, _01315_);
  and (_01318_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_01319_, _40703_, _00946_);
  and (_01320_, _40547_, _40464_);
  and (_01321_, _01320_, _01319_);
  and (_01322_, _01304_, _40381_);
  and (_01323_, _01322_, _01321_);
  and (_01324_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_01325_, _01324_, _01318_);
  and (_01326_, _01322_, _01296_);
  and (_01327_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_01328_, _00833_, _00751_);
  and (_01329_, _01328_, _01322_);
  and (_01330_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_01331_, _01330_, _01327_);
  or (_01332_, _01331_, _01325_);
  and (_01333_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_01334_, _01320_, _00758_);
  and (_01335_, _01334_, _01292_);
  and (_01336_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_01337_, _01336_, _01333_);
  and (_01338_, _01291_, _00789_);
  and (_01339_, _01338_, _01296_);
  and (_01340_, _01339_, _40266_);
  and (_01341_, _01292_, _01321_);
  and (_01342_, _01341_, _01032_);
  or (_01343_, _01342_, _01340_);
  or (_01344_, _01343_, _01337_);
  or (_01345_, _01344_, _01332_);
  and (_01346_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01347_, _01328_, _01292_);
  and (_01348_, _01347_, _00912_);
  and (_01349_, _01319_, _01290_);
  and (_01350_, _01349_, _01292_);
  and (_01351_, _01350_, _01096_);
  or (_01352_, _01351_, _01348_);
  and (_01353_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01354_, _01296_, _01292_);
  and (_01355_, _01354_, _01199_);
  or (_01356_, _01355_, _01353_);
  or (_01357_, _01356_, _01352_);
  or (_01358_, _01357_, _01346_);
  or (_01359_, _01358_, _01345_);
  and (_01360_, _01359_, _01312_);
  nor (_01361_, _01312_, _17497_);
  or (_01362_, _01361_, _01360_);
  and (_01363_, _01362_, _01317_);
  nor (_01364_, _01317_, _28011_);
  or (_01365_, _01364_, _01363_);
  and (_39650_, _01365_, _41806_);
  and (_01366_, _01294_, _00782_);
  and (_01367_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_01368_, _01304_, _01144_);
  and (_01369_, _01368_, _01173_);
  and (_01370_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01371_, _01293_, _01319_);
  and (_01372_, _01371_, _01137_);
  or (_01373_, _01372_, _01370_);
  or (_01374_, _01373_, _01369_);
  or (_01375_, _01374_, _01367_);
  and (_01376_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01377_, _01341_, _01023_);
  or (_01378_, _01377_, _01376_);
  and (_01379_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_01380_, _01339_, _40411_);
  or (_01381_, _01380_, _01379_);
  or (_01382_, _01381_, _01378_);
  and (_01383_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_01384_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_01385_, _01384_, _01383_);
  and (_01386_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_01387_, _01347_, _00903_);
  or (_01388_, _01387_, _01386_);
  or (_01389_, _01388_, _01385_);
  or (_01390_, _01389_, _01382_);
  nor (_01391_, _01390_, _01375_);
  nand (_01392_, _01391_, _01312_);
  or (_01393_, _01392_, _01366_);
  or (_01394_, _01312_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_01395_, _01394_, _01393_);
  or (_01396_, _01395_, _01315_);
  nand (_01397_, _01315_, _29231_);
  and (_01398_, _01397_, _41806_);
  and (_39713_, _01398_, _01396_);
  and (_01399_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_01400_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_01401_, _01400_, _01399_);
  and (_01402_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_01403_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_01404_, _01403_, _01402_);
  or (_01405_, _01404_, _01401_);
  and (_01407_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_01409_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_01411_, _01409_, _01407_);
  and (_01413_, _01341_, _01049_);
  and (_01415_, _01339_, _40550_);
  or (_01417_, _01415_, _01413_);
  or (_01419_, _01417_, _01411_);
  or (_01420_, _01419_, _01405_);
  and (_01421_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01422_, _01347_, _00930_);
  and (_01423_, _01350_, _01087_);
  or (_01424_, _01423_, _01422_);
  and (_01425_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_01427_, _01354_, _01157_);
  or (_01428_, _01427_, _01425_);
  or (_01430_, _01428_, _01424_);
  or (_01431_, _01430_, _01421_);
  or (_01432_, _01431_, _01420_);
  and (_01434_, _01432_, _01312_);
  nor (_01435_, _01312_, _17323_);
  or (_01436_, _01435_, _01434_);
  and (_01438_, _01436_, _01317_);
  nor (_01439_, _01317_, _29893_);
  or (_01440_, _01439_, _01438_);
  and (_39714_, _01440_, _41806_);
  and (_01442_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_01443_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01445_, _01443_, _01442_);
  and (_01446_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_01447_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_01449_, _01447_, _01446_);
  or (_01450_, _01449_, _01445_);
  and (_01451_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_01453_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_01454_, _01453_, _01451_);
  and (_01455_, _01339_, _40496_);
  and (_01457_, _01341_, _01000_);
  or (_01458_, _01457_, _01455_);
  or (_01459_, _01458_, _01454_);
  or (_01460_, _01459_, _01450_);
  and (_01461_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01462_, _01347_, _00878_);
  and (_01463_, _01350_, _01121_);
  or (_01464_, _01463_, _01462_);
  and (_01465_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_01466_, _01354_, _01190_);
  or (_01467_, _01466_, _01465_);
  or (_01468_, _01467_, _01464_);
  or (_01469_, _01468_, _01461_);
  or (_01470_, _01469_, _01460_);
  and (_01471_, _01470_, _01312_);
  nor (_01472_, _01312_, _15975_);
  or (_01473_, _01472_, _01471_);
  and (_01474_, _01473_, _01317_);
  nor (_01475_, _01317_, _30567_);
  or (_01476_, _01475_, _01474_);
  and (_39715_, _01476_, _41806_);
  and (_01478_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_01479_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_01481_, _01479_, _01478_);
  and (_01482_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_01483_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_01485_, _01483_, _01482_);
  or (_01486_, _01485_, _01481_);
  and (_01487_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_01489_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_01490_, _01489_, _01487_);
  and (_01491_, _01341_, _01039_);
  and (_01493_, _01339_, _40373_);
  or (_01494_, _01493_, _01491_);
  or (_01495_, _01494_, _01490_);
  or (_01497_, _01495_, _01486_);
  and (_01498_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01499_, _01347_, _00920_);
  and (_01501_, _01350_, _01103_);
  or (_01502_, _01501_, _01499_);
  and (_01503_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_01505_, _01354_, _01206_);
  or (_01506_, _01505_, _01503_);
  or (_01507_, _01506_, _01502_);
  or (_01509_, _01507_, _01498_);
  or (_01510_, _01509_, _01497_);
  and (_01511_, _01510_, _01312_);
  nor (_01512_, _01312_, _17007_);
  or (_01513_, _01512_, _01511_);
  and (_01514_, _01513_, _01317_);
  nor (_01515_, _01317_, _31338_);
  or (_01516_, _01515_, _01514_);
  and (_39716_, _01516_, _41806_);
  and (_01517_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_01518_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or (_01519_, _01518_, _01517_);
  and (_01520_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_01521_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01522_, _01521_, _01520_);
  or (_01523_, _01522_, _01519_);
  and (_01524_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_01525_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_01526_, _01525_, _01524_);
  and (_01527_, _01339_, _40511_);
  and (_01528_, _01341_, _01016_);
  or (_01530_, _01528_, _01527_);
  or (_01531_, _01530_, _01526_);
  or (_01533_, _01531_, _01523_);
  and (_01534_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01535_, _01347_, _00896_);
  and (_01537_, _01350_, _01130_);
  or (_01538_, _01537_, _01535_);
  and (_01539_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01541_, _01354_, _01166_);
  or (_01542_, _01541_, _01539_);
  or (_01543_, _01542_, _01538_);
  or (_01545_, _01543_, _01534_);
  or (_01546_, _01545_, _01533_);
  and (_01547_, _01546_, _01312_);
  nor (_01549_, _01312_, _16172_);
  or (_01550_, _01549_, _01547_);
  and (_01551_, _01550_, _01317_);
  nor (_01553_, _01317_, _32044_);
  or (_01554_, _01553_, _01551_);
  and (_39717_, _01554_, _41806_);
  and (_01556_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01557_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_01558_, _01557_, _01556_);
  and (_01560_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_01561_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01562_, _01561_, _01560_);
  or (_01563_, _01562_, _01558_);
  and (_01564_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_01565_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_01566_, _01565_, _01564_);
  and (_01567_, _01339_, _40427_);
  and (_01568_, _01341_, _01056_);
  or (_01569_, _01568_, _01567_);
  or (_01570_, _01569_, _01566_);
  or (_01571_, _01570_, _01563_);
  and (_01572_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01573_, _01347_, _00937_);
  and (_01574_, _01350_, _01080_);
  or (_01575_, _01574_, _01573_);
  and (_01576_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01577_, _01354_, _01150_);
  or (_01578_, _01577_, _01576_);
  or (_01579_, _01578_, _01575_);
  or (_01580_, _01579_, _01572_);
  or (_01582_, _01580_, _01571_);
  and (_01583_, _01582_, _01312_);
  nor (_01585_, _01312_, _17160_);
  or (_01586_, _01585_, _01583_);
  and (_01587_, _01586_, _01317_);
  nor (_01589_, _01317_, _32853_);
  or (_01590_, _01589_, _01587_);
  and (_39718_, _01590_, _41806_);
  and (_01592_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01593_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_01594_, _01593_, _01592_);
  and (_01596_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_01597_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_01598_, _01597_, _01596_);
  or (_01600_, _01598_, _01594_);
  and (_01601_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_01602_, _01335_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_01604_, _01602_, _01601_);
  and (_01605_, _01339_, _40695_);
  and (_01606_, _01341_, _01007_);
  or (_01608_, _01606_, _01605_);
  or (_01609_, _01608_, _01604_);
  or (_01610_, _01609_, _01600_);
  and (_01612_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01613_, _01347_, _00885_);
  and (_01614_, _01350_, _01114_);
  or (_01615_, _01614_, _01613_);
  and (_01616_, _01294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01617_, _01354_, _01183_);
  or (_01618_, _01617_, _01616_);
  or (_01619_, _01618_, _01615_);
  or (_01620_, _01619_, _01612_);
  or (_01621_, _01620_, _01610_);
  and (_01622_, _01621_, _01312_);
  nor (_01623_, _01312_, _16512_);
  or (_01624_, _01623_, _01622_);
  and (_01625_, _01624_, _01317_);
  nor (_01626_, _01317_, _33598_);
  or (_01627_, _01626_, _01625_);
  and (_39719_, _01627_, _41806_);
  and (_39764_, _40734_, _41806_);
  and (_39765_, _40870_, _41806_);
  nor (_39767_, _40500_, rst);
  and (_39783_, _40888_, _41806_);
  and (_39784_, _40901_, _41806_);
  and (_39785_, _40914_, _41806_);
  and (_39786_, _40922_, _41806_);
  and (_39787_, _40932_, _41806_);
  and (_39788_, _40942_, _41806_);
  and (_39789_, _40952_, _41806_);
  nor (_39790_, _40415_, rst);
  nor (_39791_, _40611_, rst);
  not (_01632_, _41697_);
  nor (_01633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01635_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01636_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01635_);
  nor (_01637_, _01636_, _01633_);
  nor (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01640_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01635_);
  nor (_01641_, _01640_, _01639_);
  not (_01643_, _01641_);
  nor (_01644_, _01643_, _01637_);
  nor (_01645_, _00129_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01647_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01635_);
  nor (_01648_, _01647_, _01645_);
  not (_01649_, _01648_);
  nor (_01651_, _01641_, _01637_);
  not (_01652_, _01651_);
  nor (_01653_, _00110_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01654_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01635_);
  nor (_01655_, _01654_, _01653_);
  and (_01656_, _01655_, _01652_);
  or (_01657_, _01656_, _01649_);
  nor (_01658_, _01655_, _01652_);
  or (_01659_, _01658_, _01648_);
  and (_01660_, _01659_, _01657_);
  and (_01661_, _01660_, _01644_);
  and (_01662_, _01661_, _01632_);
  not (_01663_, _41738_);
  and (_01664_, _01641_, _01637_);
  and (_01665_, _01660_, _01664_);
  and (_01666_, _01665_, _01663_);
  or (_01667_, _01666_, _01662_);
  not (_01668_, _41656_);
  and (_01669_, _01643_, _01637_);
  and (_01670_, _01669_, _01660_);
  and (_01671_, _01670_, _01668_);
  not (_01673_, _42040_);
  and (_01674_, _01649_, _01655_);
  and (_01676_, _01674_, _01644_);
  and (_01677_, _01676_, _01673_);
  not (_01678_, _42081_);
  and (_01680_, _01674_, _01664_);
  and (_01681_, _01680_, _01678_);
  or (_01682_, _01681_, _01677_);
  not (_01684_, _41999_);
  and (_01685_, _01669_, _01674_);
  and (_01686_, _01685_, _01684_);
  not (_01688_, _41786_);
  and (_01689_, _01658_, _01649_);
  and (_01690_, _01689_, _01688_);
  or (_01692_, _01690_, _01686_);
  or (_01693_, _01692_, _01682_);
  or (_01694_, _01693_, _01671_);
  or (_01696_, _01694_, _01667_);
  not (_01697_, _41917_);
  nor (_01698_, _01658_, _01656_);
  and (_01700_, _01698_, _01649_);
  and (_01701_, _01700_, _01664_);
  and (_01702_, _01701_, _01697_);
  not (_01704_, _42204_);
  and (_01705_, _01698_, _01648_);
  and (_01706_, _01705_, _01644_);
  and (_01707_, _01706_, _01704_);
  not (_01708_, _42163_);
  and (_01709_, _01705_, _01669_);
  and (_01710_, _01709_, _01708_);
  or (_01711_, _01710_, _01707_);
  or (_01712_, _01711_, _01702_);
  not (_01713_, _41876_);
  and (_01714_, _01700_, _01644_);
  and (_01715_, _01714_, _01713_);
  not (_01716_, _41958_);
  and (_01717_, _01674_, _01651_);
  and (_01718_, _01717_, _01716_);
  not (_01719_, _42286_);
  and (_01720_, _01655_, _01651_);
  and (_01721_, _01720_, _01648_);
  and (_01722_, _01721_, _01719_);
  not (_01723_, _42122_);
  and (_01724_, _01658_, _01648_);
  and (_01726_, _01724_, _01723_);
  or (_01727_, _01726_, _01722_);
  or (_01729_, _01727_, _01718_);
  or (_01730_, _01729_, _01715_);
  not (_01731_, _42245_);
  and (_01733_, _01705_, _01664_);
  and (_01734_, _01733_, _01731_);
  not (_01735_, _41835_);
  and (_01737_, _01700_, _01669_);
  and (_01738_, _01737_, _01735_);
  or (_01739_, _01738_, _01734_);
  or (_01741_, _01739_, _01730_);
  or (_01742_, _01741_, _01712_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01742_, _01696_);
  and (_01744_, _01661_, _01719_);
  and (_01745_, _01680_, _01684_);
  and (_01746_, _01676_, _01716_);
  or (_01748_, _01746_, _01745_);
  and (_01749_, _01689_, _01632_);
  and (_01750_, _01685_, _01697_);
  or (_01752_, _01750_, _01749_);
  or (_01753_, _01752_, _01748_);
  or (_01754_, _01753_, _01744_);
  and (_01756_, _01665_, _01668_);
  and (_01757_, _01670_, _01731_);
  or (_01758_, _01757_, _01756_);
  or (_01759_, _01758_, _01754_);
  and (_01760_, _01737_, _01663_);
  and (_01761_, _01714_, _01688_);
  and (_01762_, _01706_, _01723_);
  or (_01763_, _01762_, _01761_);
  or (_01764_, _01763_, _01760_);
  and (_01765_, _01709_, _01678_);
  and (_01766_, _01717_, _01713_);
  and (_01767_, _01724_, _01673_);
  and (_01768_, _01721_, _01704_);
  or (_01769_, _01768_, _01767_);
  or (_01770_, _01769_, _01766_);
  or (_01771_, _01770_, _01765_);
  and (_01772_, _01701_, _01735_);
  and (_01773_, _01733_, _01708_);
  or (_01774_, _01773_, _01772_);
  or (_01775_, _01774_, _01771_);
  or (_01776_, _01775_, _01764_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01776_, _01759_);
  and (_01778_, _01665_, _01632_);
  and (_01780_, _01717_, _01697_);
  and (_01781_, _01676_, _01684_);
  or (_01782_, _01781_, _01780_);
  and (_01784_, _01689_, _01663_);
  and (_01785_, _01680_, _01673_);
  or (_01786_, _01785_, _01784_);
  or (_01788_, _01786_, _01782_);
  or (_01789_, _01788_, _01778_);
  and (_01790_, _01670_, _01719_);
  and (_01792_, _01661_, _01668_);
  or (_01793_, _01792_, _01790_);
  or (_01794_, _01793_, _01789_);
  and (_01796_, _01714_, _01735_);
  and (_01797_, _01701_, _01713_);
  and (_01798_, _01709_, _01723_);
  or (_01800_, _01798_, _01797_);
  or (_01801_, _01800_, _01796_);
  and (_01802_, _01737_, _01688_);
  and (_01804_, _01685_, _01716_);
  and (_01805_, _01724_, _01678_);
  and (_01806_, _01721_, _01731_);
  or (_01808_, _01806_, _01805_);
  or (_01809_, _01808_, _01804_);
  or (_01810_, _01809_, _01802_);
  and (_01811_, _01733_, _01704_);
  and (_01812_, _01706_, _01708_);
  or (_01813_, _01812_, _01811_);
  or (_01814_, _01813_, _01810_);
  or (_01815_, _01814_, _01801_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01815_, _01794_);
  and (_01816_, _01665_, _01719_);
  and (_01817_, _01661_, _01731_);
  or (_01818_, _01817_, _01816_);
  and (_01819_, _01670_, _01704_);
  and (_01820_, _01676_, _01697_);
  and (_01821_, _01685_, _01713_);
  or (_01822_, _01821_, _01820_);
  and (_01823_, _01689_, _01668_);
  and (_01824_, _01717_, _01735_);
  or (_01825_, _01824_, _01823_);
  or (_01826_, _01825_, _01822_);
  or (_01827_, _01826_, _01819_);
  or (_01829_, _01827_, _01818_);
  and (_01830_, _01714_, _01663_);
  and (_01832_, _01733_, _01723_);
  and (_01833_, _01737_, _01632_);
  or (_01834_, _01833_, _01832_);
  or (_01836_, _01834_, _01830_);
  and (_01837_, _01709_, _01673_);
  and (_01838_, _01680_, _01716_);
  and (_01840_, _01721_, _01708_);
  and (_01841_, _01724_, _01684_);
  or (_01842_, _01841_, _01840_);
  or (_01844_, _01842_, _01838_);
  or (_01845_, _01844_, _01837_);
  and (_01846_, _01706_, _01678_);
  and (_01848_, _01701_, _01688_);
  or (_01849_, _01848_, _01846_);
  or (_01850_, _01849_, _01845_);
  or (_01852_, _01850_, _01836_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01852_, _01829_);
  not (_01853_, _41743_);
  and (_01855_, _01665_, _01853_);
  not (_01856_, _41791_);
  and (_01857_, _01689_, _01856_);
  not (_01859_, _42086_);
  and (_01860_, _01680_, _01859_);
  or (_01861_, _01860_, _01857_);
  not (_01862_, _42045_);
  and (_01863_, _01676_, _01862_);
  not (_01864_, _42004_);
  and (_01865_, _01685_, _01864_);
  or (_01866_, _01865_, _01863_);
  or (_01867_, _01866_, _01861_);
  or (_01868_, _01867_, _01855_);
  not (_01869_, _41661_);
  and (_01870_, _01670_, _01869_);
  not (_01871_, _41702_);
  and (_01872_, _01661_, _01871_);
  or (_01873_, _01872_, _01870_);
  or (_01874_, _01873_, _01868_);
  not (_01875_, _42168_);
  and (_01876_, _01709_, _01875_);
  not (_01877_, _41922_);
  and (_01878_, _01701_, _01877_);
  not (_01879_, _42209_);
  and (_01881_, _01706_, _01879_);
  or (_01882_, _01881_, _01878_);
  or (_01884_, _01882_, _01876_);
  not (_01885_, _41881_);
  and (_01886_, _01714_, _01885_);
  not (_01888_, _41963_);
  and (_01889_, _01717_, _01888_);
  not (_01890_, _42291_);
  and (_01892_, _01721_, _01890_);
  not (_01893_, _42127_);
  and (_01894_, _01724_, _01893_);
  or (_01896_, _01894_, _01892_);
  or (_01897_, _01896_, _01889_);
  or (_01898_, _01897_, _01886_);
  not (_01900_, _41840_);
  and (_01901_, _01737_, _01900_);
  not (_01902_, _42250_);
  and (_01904_, _01733_, _01902_);
  or (_01905_, _01904_, _01901_);
  or (_01906_, _01905_, _01898_);
  or (_01908_, _01906_, _01884_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01908_, _01874_);
  not (_01909_, _41749_);
  and (_01911_, _01665_, _01909_);
  not (_01912_, _42050_);
  and (_01913_, _01676_, _01912_);
  not (_01914_, _42091_);
  and (_01915_, _01680_, _01914_);
  or (_01916_, _01915_, _01913_);
  not (_01917_, _41968_);
  and (_01918_, _01717_, _01917_);
  not (_01919_, _42009_);
  and (_01920_, _01685_, _01919_);
  or (_01921_, _01920_, _01918_);
  or (_01922_, _01921_, _01916_);
  or (_01923_, _01922_, _01911_);
  not (_01924_, _41666_);
  and (_01925_, _01670_, _01924_);
  not (_01926_, _41707_);
  and (_01927_, _01661_, _01926_);
  or (_01928_, _01927_, _01925_);
  or (_01929_, _01928_, _01923_);
  not (_01930_, _41886_);
  and (_01931_, _01714_, _01930_);
  not (_01933_, _41927_);
  and (_01934_, _01701_, _01933_);
  or (_01936_, _01934_, _01931_);
  not (_01937_, _42214_);
  and (_01938_, _01706_, _01937_);
  or (_01940_, _01938_, _01936_);
  not (_01941_, _42173_);
  and (_01942_, _01709_, _01941_);
  not (_01944_, _41801_);
  and (_01945_, _01689_, _01944_);
  not (_01946_, _42296_);
  and (_01948_, _01721_, _01946_);
  not (_01949_, _42132_);
  and (_01950_, _01724_, _01949_);
  or (_01952_, _01950_, _01948_);
  or (_01953_, _01952_, _01945_);
  or (_01954_, _01953_, _01942_);
  not (_01956_, _41845_);
  and (_01957_, _01737_, _01956_);
  not (_01958_, _42255_);
  and (_01960_, _01733_, _01958_);
  or (_01961_, _01960_, _01957_);
  or (_01962_, _01961_, _01954_);
  or (_01964_, _01962_, _01940_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01964_, _01929_);
  not (_01965_, _41671_);
  and (_01966_, _01670_, _01965_);
  not (_01967_, _41758_);
  and (_01968_, _01665_, _01967_);
  or (_01969_, _01968_, _01966_);
  not (_01970_, _41712_);
  and (_01971_, _01661_, _01970_);
  not (_01972_, _42096_);
  and (_01973_, _01680_, _01972_);
  not (_01974_, _42055_);
  and (_01975_, _01676_, _01974_);
  or (_01976_, _01975_, _01973_);
  not (_01977_, _41973_);
  and (_01978_, _01717_, _01977_);
  not (_01979_, _41809_);
  and (_01980_, _01689_, _01979_);
  or (_01981_, _01980_, _01978_);
  or (_01982_, _01981_, _01976_);
  or (_01983_, _01982_, _01971_);
  or (_01985_, _01983_, _01969_);
  not (_01986_, _41891_);
  and (_01988_, _01714_, _01986_);
  not (_01989_, _42260_);
  and (_01990_, _01733_, _01989_);
  not (_01992_, _41932_);
  and (_01993_, _01701_, _01992_);
  or (_01994_, _01993_, _01990_);
  or (_01996_, _01994_, _01988_);
  not (_01997_, _42219_);
  and (_01998_, _01706_, _01997_);
  not (_02000_, _42014_);
  and (_02001_, _01685_, _02000_);
  not (_02002_, _42301_);
  and (_02004_, _01721_, _02002_);
  not (_02005_, _42137_);
  and (_02006_, _01724_, _02005_);
  or (_02008_, _02006_, _02004_);
  or (_02009_, _02008_, _02001_);
  or (_02010_, _02009_, _01998_);
  not (_02012_, _42178_);
  and (_02013_, _01709_, _02012_);
  not (_02014_, _41850_);
  and (_02016_, _01737_, _02014_);
  or (_02017_, _02016_, _02013_);
  or (_02018_, _02017_, _02010_);
  or (_02019_, _02018_, _01996_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _02019_, _01985_);
  not (_02020_, _41676_);
  and (_02021_, _01670_, _02020_);
  not (_02022_, _41765_);
  and (_02023_, _01665_, _02022_);
  or (_02024_, _02023_, _02021_);
  not (_02025_, _41978_);
  and (_02026_, _01717_, _02025_);
  not (_02027_, _42019_);
  and (_02028_, _01685_, _02027_);
  or (_02029_, _02028_, _02026_);
  not (_02030_, _42101_);
  and (_02031_, _01680_, _02030_);
  not (_02032_, _42060_);
  and (_02033_, _01676_, _02032_);
  or (_02034_, _02033_, _02031_);
  or (_02035_, _02034_, _02029_);
  not (_02037_, _41717_);
  and (_02038_, _01661_, _02037_);
  or (_02040_, _02038_, _02035_);
  or (_02041_, _02040_, _02024_);
  not (_02042_, _41937_);
  and (_02044_, _01701_, _02042_);
  not (_02045_, _42224_);
  and (_02046_, _01706_, _02045_);
  not (_02048_, _41896_);
  and (_02049_, _01714_, _02048_);
  or (_02050_, _02049_, _02046_);
  or (_02052_, _02050_, _02044_);
  not (_02053_, _41855_);
  and (_02054_, _01737_, _02053_);
  not (_02056_, _41814_);
  and (_02057_, _01689_, _02056_);
  not (_02058_, _42306_);
  and (_02060_, _01721_, _02058_);
  not (_02061_, _42142_);
  and (_02062_, _01724_, _02061_);
  or (_02064_, _02062_, _02060_);
  or (_02065_, _02064_, _02057_);
  or (_02066_, _02065_, _02054_);
  not (_02068_, _42265_);
  and (_02069_, _01733_, _02068_);
  not (_02070_, _42183_);
  and (_02071_, _01709_, _02070_);
  or (_02072_, _02071_, _02069_);
  or (_02073_, _02072_, _02066_);
  or (_02074_, _02073_, _02052_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _02074_, _02041_);
  not (_02075_, _41681_);
  and (_02076_, _01670_, _02075_);
  not (_02077_, _41770_);
  and (_02078_, _01665_, _02077_);
  or (_02079_, _02078_, _02076_);
  not (_02080_, _41722_);
  and (_02081_, _01661_, _02080_);
  not (_02082_, _42065_);
  and (_02083_, _01676_, _02082_);
  not (_02084_, _42106_);
  and (_02085_, _01680_, _02084_);
  or (_02086_, _02085_, _02083_);
  not (_02087_, _41983_);
  and (_02089_, _01717_, _02087_);
  not (_02090_, _42024_);
  and (_02092_, _01685_, _02090_);
  or (_02093_, _02092_, _02089_);
  or (_02094_, _02093_, _02086_);
  or (_02096_, _02094_, _02081_);
  or (_02097_, _02096_, _02079_);
  not (_02098_, _42270_);
  and (_02100_, _01733_, _02098_);
  not (_02101_, _41901_);
  and (_02102_, _01714_, _02101_);
  not (_02104_, _42229_);
  and (_02105_, _01706_, _02104_);
  or (_02106_, _02105_, _02102_);
  or (_02108_, _02106_, _02100_);
  not (_02109_, _42188_);
  and (_02110_, _01709_, _02109_);
  not (_02112_, _41819_);
  and (_02113_, _01689_, _02112_);
  not (_02114_, _42311_);
  and (_02116_, _01721_, _02114_);
  not (_02117_, _42147_);
  and (_02118_, _01724_, _02117_);
  or (_02120_, _02118_, _02116_);
  or (_02121_, _02120_, _02113_);
  or (_02122_, _02121_, _02110_);
  not (_02123_, _41942_);
  and (_02124_, _01701_, _02123_);
  not (_02125_, _41860_);
  and (_02126_, _01737_, _02125_);
  or (_02127_, _02126_, _02124_);
  or (_02128_, _02127_, _02122_);
  or (_02129_, _02128_, _02108_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _02129_, _02097_);
  not (_02130_, _41727_);
  and (_02131_, _01661_, _02130_);
  not (_02132_, _41775_);
  and (_02133_, _01665_, _02132_);
  or (_02134_, _02133_, _02131_);
  not (_02135_, _41686_);
  and (_02136_, _01670_, _02135_);
  not (_02137_, _42111_);
  and (_02138_, _01680_, _02137_);
  not (_02139_, _41824_);
  and (_02141_, _01689_, _02139_);
  or (_02142_, _02141_, _02138_);
  not (_02144_, _42070_);
  and (_02145_, _01676_, _02144_);
  not (_02146_, _41988_);
  and (_02148_, _01717_, _02146_);
  or (_02149_, _02148_, _02145_);
  or (_02150_, _02149_, _02142_);
  or (_02152_, _02150_, _02136_);
  or (_02153_, _02152_, _02134_);
  not (_02154_, _42275_);
  and (_02156_, _01733_, _02154_);
  not (_02157_, _42193_);
  and (_02158_, _01709_, _02157_);
  not (_02160_, _41947_);
  and (_02161_, _01701_, _02160_);
  or (_02162_, _02161_, _02158_);
  or (_02164_, _02162_, _02156_);
  not (_02165_, _42234_);
  and (_02166_, _01706_, _02165_);
  not (_02168_, _42029_);
  and (_02169_, _01685_, _02168_);
  not (_02170_, _42316_);
  and (_02172_, _01721_, _02170_);
  not (_02173_, _42152_);
  and (_02174_, _01724_, _02173_);
  or (_02175_, _02174_, _02172_);
  or (_02176_, _02175_, _02169_);
  or (_02177_, _02176_, _02166_);
  not (_02178_, _41906_);
  and (_02179_, _01714_, _02178_);
  not (_02180_, _41865_);
  and (_02181_, _01737_, _02180_);
  or (_02182_, _02181_, _02179_);
  or (_02183_, _02182_, _02177_);
  or (_02184_, _02183_, _02164_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _02184_, _02153_);
  not (_02185_, _41691_);
  and (_02186_, _01670_, _02185_);
  not (_02187_, _41780_);
  and (_02188_, _01665_, _02187_);
  or (_02189_, _02188_, _02186_);
  not (_02190_, _41732_);
  and (_02191_, _01661_, _02190_);
  not (_02193_, _42116_);
  and (_02194_, _01680_, _02193_);
  not (_02196_, _42075_);
  and (_02197_, _01676_, _02196_);
  or (_02198_, _02197_, _02194_);
  not (_02200_, _42034_);
  and (_02201_, _01685_, _02200_);
  not (_02202_, _41829_);
  and (_02204_, _01689_, _02202_);
  or (_02205_, _02204_, _02201_);
  or (_02206_, _02205_, _02198_);
  or (_02208_, _02206_, _02191_);
  or (_02209_, _02208_, _02189_);
  not (_02210_, _41952_);
  and (_02212_, _01701_, _02210_);
  not (_02213_, _41911_);
  and (_02214_, _01714_, _02213_);
  or (_02216_, _02214_, _02212_);
  not (_02217_, _41870_);
  and (_02218_, _01737_, _02217_);
  or (_02220_, _02218_, _02216_);
  not (_02221_, _42280_);
  and (_02222_, _01733_, _02221_);
  not (_02224_, _41993_);
  and (_02225_, _01717_, _02224_);
  not (_02226_, _42321_);
  and (_02227_, _01721_, _02226_);
  not (_02228_, _42157_);
  and (_02229_, _01724_, _02228_);
  or (_02230_, _02229_, _02227_);
  or (_02231_, _02230_, _02225_);
  or (_02232_, _02231_, _02222_);
  not (_02233_, _42239_);
  and (_02234_, _01706_, _02233_);
  not (_02235_, _42198_);
  and (_02236_, _01709_, _02235_);
  or (_02237_, _02236_, _02234_);
  or (_02238_, _02237_, _02232_);
  or (_02239_, _02238_, _02220_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _02239_, _02209_);
  and (_02240_, _01665_, _01871_);
  and (_02241_, _01680_, _01862_);
  and (_02242_, _01685_, _01888_);
  or (_02243_, _02242_, _02241_);
  and (_02244_, _01689_, _01853_);
  and (_02245_, _01676_, _01864_);
  or (_02246_, _02245_, _02244_);
  or (_02247_, _02246_, _02243_);
  or (_02248_, _02247_, _02240_);
  and (_02249_, _01670_, _01890_);
  and (_02250_, _01661_, _01869_);
  or (_02251_, _02250_, _02249_);
  or (_02252_, _02251_, _02248_);
  and (_02253_, _01709_, _01893_);
  and (_02254_, _01714_, _01900_);
  and (_02255_, _01706_, _01875_);
  or (_02256_, _02255_, _02254_);
  or (_02257_, _02256_, _02253_);
  and (_02258_, _01737_, _01856_);
  and (_02259_, _01717_, _01877_);
  and (_02260_, _01724_, _01859_);
  and (_02261_, _01721_, _01902_);
  or (_02262_, _02261_, _02260_);
  or (_02263_, _02262_, _02259_);
  or (_02264_, _02263_, _02258_);
  and (_02265_, _01701_, _01885_);
  and (_02266_, _01733_, _01879_);
  or (_02267_, _02266_, _02265_);
  or (_02268_, _02267_, _02264_);
  or (_02269_, _02268_, _02257_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _02269_, _02252_);
  and (_02270_, _01665_, _01926_);
  and (_02271_, _01689_, _01909_);
  and (_02272_, _01680_, _01912_);
  or (_02273_, _02272_, _02271_);
  and (_02274_, _01717_, _01933_);
  and (_02275_, _01676_, _01919_);
  or (_02276_, _02275_, _02274_);
  or (_02277_, _02276_, _02273_);
  or (_02278_, _02277_, _02270_);
  and (_02279_, _01670_, _01946_);
  and (_02280_, _01661_, _01924_);
  or (_02281_, _02280_, _02279_);
  or (_02282_, _02281_, _02278_);
  and (_02283_, _01706_, _01941_);
  and (_02284_, _01714_, _01956_);
  and (_02285_, _01733_, _01937_);
  or (_02286_, _02285_, _02284_);
  or (_02287_, _02286_, _02283_);
  and (_02288_, _01737_, _01944_);
  and (_02289_, _01685_, _01917_);
  and (_02290_, _01724_, _01914_);
  and (_02291_, _01721_, _01958_);
  or (_02292_, _02291_, _02290_);
  or (_02293_, _02292_, _02289_);
  or (_02294_, _02293_, _02288_);
  and (_02295_, _01701_, _01930_);
  and (_02296_, _01709_, _01949_);
  or (_02297_, _02296_, _02295_);
  or (_02298_, _02297_, _02294_);
  or (_02299_, _02298_, _02287_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _02299_, _02282_);
  and (_02300_, _01661_, _01965_);
  and (_02301_, _01689_, _01967_);
  and (_02302_, _01685_, _01977_);
  or (_02303_, _02302_, _02301_);
  and (_02304_, _01680_, _01974_);
  and (_02305_, _01676_, _02000_);
  or (_02306_, _02305_, _02304_);
  or (_02307_, _02306_, _02303_);
  or (_02308_, _02307_, _02300_);
  and (_02309_, _01670_, _02002_);
  and (_02310_, _01665_, _01970_);
  or (_02311_, _02310_, _02309_);
  or (_02312_, _02311_, _02308_);
  and (_02313_, _01714_, _02014_);
  and (_02314_, _01737_, _01979_);
  or (_02315_, _02314_, _02313_);
  and (_02316_, _01701_, _01986_);
  or (_02317_, _02316_, _02315_);
  and (_02318_, _01709_, _02005_);
  and (_02319_, _01717_, _01992_);
  and (_02320_, _01724_, _01972_);
  and (_02321_, _01721_, _01989_);
  or (_02322_, _02321_, _02320_);
  or (_02323_, _02322_, _02319_);
  or (_02324_, _02323_, _02318_);
  and (_02325_, _01733_, _01997_);
  and (_02326_, _01706_, _02012_);
  or (_02327_, _02326_, _02325_);
  or (_02328_, _02327_, _02324_);
  or (_02329_, _02328_, _02317_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _02329_, _02312_);
  and (_02330_, _01665_, _02037_);
  and (_02331_, _01685_, _02025_);
  and (_02332_, _01717_, _02042_);
  or (_02333_, _02332_, _02331_);
  and (_02334_, _01680_, _02032_);
  and (_02335_, _01676_, _02027_);
  or (_02336_, _02335_, _02334_);
  or (_02337_, _02336_, _02333_);
  or (_02338_, _02337_, _02330_);
  and (_02339_, _01670_, _02058_);
  and (_02340_, _01661_, _02020_);
  or (_02341_, _02340_, _02339_);
  or (_02342_, _02341_, _02338_);
  and (_02343_, _01733_, _02045_);
  and (_02344_, _01706_, _02070_);
  and (_02345_, _01701_, _02048_);
  or (_02346_, _02345_, _02344_);
  or (_02347_, _02346_, _02343_);
  and (_02348_, _01737_, _02056_);
  and (_02349_, _01714_, _02053_);
  or (_02350_, _02349_, _02348_);
  and (_02351_, _01709_, _02061_);
  and (_02352_, _01689_, _02022_);
  and (_02353_, _01721_, _02068_);
  and (_02354_, _01724_, _02030_);
  or (_02355_, _02354_, _02353_);
  or (_02356_, _02355_, _02352_);
  or (_02357_, _02356_, _02351_);
  or (_02358_, _02357_, _02350_);
  or (_02359_, _02358_, _02347_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02359_, _02342_);
  and (_02360_, _01661_, _02075_);
  and (_02361_, _01680_, _02082_);
  and (_02362_, _01689_, _02077_);
  or (_02363_, _02362_, _02361_);
  and (_02364_, _01676_, _02090_);
  and (_02365_, _01717_, _02123_);
  or (_02366_, _02365_, _02364_);
  or (_02367_, _02366_, _02363_);
  or (_02368_, _02367_, _02360_);
  and (_02369_, _01670_, _02114_);
  and (_02370_, _01665_, _02080_);
  or (_02371_, _02370_, _02369_);
  or (_02372_, _02371_, _02368_);
  and (_02373_, _01733_, _02104_);
  and (_02374_, _01701_, _02101_);
  and (_02375_, _01737_, _02112_);
  or (_02376_, _02375_, _02374_);
  or (_02377_, _02376_, _02373_);
  and (_02378_, _01709_, _02117_);
  and (_02379_, _01706_, _02109_);
  or (_02380_, _02379_, _02378_);
  and (_02381_, _01714_, _02125_);
  and (_02382_, _01685_, _02087_);
  and (_02383_, _01721_, _02098_);
  and (_02384_, _01724_, _02084_);
  or (_02385_, _02384_, _02383_);
  or (_02386_, _02385_, _02382_);
  or (_02387_, _02386_, _02381_);
  or (_02388_, _02387_, _02380_);
  or (_02389_, _02388_, _02377_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _02389_, _02372_);
  and (_02390_, _01665_, _02130_);
  and (_02391_, _01676_, _02168_);
  and (_02392_, _01689_, _02132_);
  or (_02393_, _02392_, _02391_);
  and (_02394_, _01685_, _02146_);
  and (_02395_, _01717_, _02160_);
  or (_02396_, _02395_, _02394_);
  or (_02397_, _02396_, _02393_);
  or (_02398_, _02397_, _02390_);
  and (_02399_, _01670_, _02170_);
  and (_02400_, _01661_, _02135_);
  or (_02401_, _02400_, _02399_);
  or (_02402_, _02401_, _02398_);
  and (_02403_, _01733_, _02165_);
  and (_02404_, _01701_, _02178_);
  and (_02405_, _01714_, _02180_);
  or (_02406_, _02405_, _02404_);
  or (_02407_, _02406_, _02403_);
  and (_02408_, _01709_, _02173_);
  and (_02409_, _01706_, _02157_);
  or (_02410_, _02409_, _02408_);
  and (_02411_, _01737_, _02139_);
  and (_02412_, _01680_, _02144_);
  and (_02413_, _01721_, _02154_);
  and (_02414_, _01724_, _02137_);
  or (_02415_, _02414_, _02413_);
  or (_02416_, _02415_, _02412_);
  or (_02417_, _02416_, _02411_);
  or (_02418_, _02417_, _02410_);
  or (_02419_, _02418_, _02407_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _02419_, _02402_);
  and (_02420_, _01670_, _02226_);
  and (_02421_, _01680_, _02196_);
  and (_02422_, _01685_, _02224_);
  or (_02423_, _02422_, _02421_);
  and (_02424_, _01676_, _02200_);
  and (_02425_, _01689_, _02187_);
  or (_02426_, _02425_, _02424_);
  or (_02427_, _02426_, _02423_);
  or (_02428_, _02427_, _02420_);
  and (_02429_, _01661_, _02185_);
  and (_02430_, _01665_, _02190_);
  or (_02431_, _02430_, _02429_);
  or (_02432_, _02431_, _02428_);
  and (_02433_, _01706_, _02235_);
  and (_02434_, _01733_, _02233_);
  and (_02435_, _01701_, _02213_);
  or (_02436_, _02435_, _02434_);
  or (_02437_, _02436_, _02433_);
  and (_02438_, _01714_, _02217_);
  and (_02439_, _01717_, _02210_);
  and (_02440_, _01721_, _02221_);
  and (_02441_, _01724_, _02193_);
  or (_02442_, _02441_, _02440_);
  or (_02443_, _02442_, _02439_);
  or (_02444_, _02443_, _02438_);
  and (_02445_, _01709_, _02228_);
  and (_02446_, _01737_, _02202_);
  or (_02447_, _02446_, _02445_);
  or (_02448_, _02447_, _02444_);
  or (_02449_, _02448_, _02437_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02449_, _02432_);
  and (_02450_, _01661_, _01890_);
  and (_02451_, _01670_, _01902_);
  or (_02452_, _02451_, _02450_);
  and (_02453_, _01665_, _01869_);
  and (_02454_, _01685_, _01877_);
  and (_02455_, _01676_, _01888_);
  or (_02456_, _02455_, _02454_);
  and (_02457_, _01717_, _01885_);
  and (_02458_, _01680_, _01864_);
  or (_02459_, _02458_, _02457_);
  or (_02460_, _02459_, _02456_);
  or (_02461_, _02460_, _02453_);
  or (_02462_, _02461_, _02452_);
  and (_02463_, _01706_, _01893_);
  and (_02464_, _01701_, _01900_);
  and (_02466_, _01733_, _01875_);
  or (_02467_, _02466_, _02464_);
  or (_02468_, _02467_, _02463_);
  and (_02469_, _01737_, _01853_);
  and (_02470_, _01689_, _01871_);
  and (_02471_, _01724_, _01862_);
  and (_02472_, _01721_, _01879_);
  or (_02473_, _02472_, _02471_);
  or (_02474_, _02473_, _02470_);
  or (_02475_, _02474_, _02469_);
  and (_02476_, _01714_, _01856_);
  and (_02477_, _01709_, _01859_);
  or (_02478_, _02477_, _02476_);
  or (_02479_, _02478_, _02475_);
  or (_02480_, _02479_, _02468_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _02480_, _02462_);
  and (_02481_, _01661_, _01946_);
  and (_02482_, _01676_, _01917_);
  and (_02483_, _01685_, _01933_);
  or (_02484_, _02483_, _02482_);
  and (_02485_, _01717_, _01930_);
  and (_02486_, _01689_, _01926_);
  or (_02487_, _02486_, _02485_);
  or (_02488_, _02487_, _02484_);
  or (_02489_, _02488_, _02481_);
  and (_02490_, _01670_, _01958_);
  and (_02491_, _01665_, _01924_);
  or (_02492_, _02491_, _02490_);
  or (_02493_, _02492_, _02489_);
  and (_02494_, _01706_, _01949_);
  and (_02495_, _01709_, _01914_);
  and (_02496_, _01737_, _01909_);
  or (_02497_, _02496_, _02495_);
  or (_02498_, _02497_, _02494_);
  and (_02499_, _01701_, _01956_);
  and (_02500_, _01714_, _01944_);
  or (_02501_, _02500_, _02499_);
  and (_02502_, _01733_, _01941_);
  and (_02503_, _01680_, _01919_);
  and (_02504_, _01721_, _01937_);
  and (_02505_, _01724_, _01912_);
  or (_02506_, _02505_, _02504_);
  or (_02507_, _02506_, _02503_);
  or (_02508_, _02507_, _02502_);
  or (_02509_, _02508_, _02501_);
  or (_02510_, _02509_, _02498_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _02510_, _02493_);
  and (_02511_, _01661_, _02002_);
  and (_02512_, _01670_, _01989_);
  or (_02513_, _02512_, _02511_);
  and (_02514_, _01665_, _01965_);
  and (_02515_, _01676_, _01977_);
  and (_02516_, _01685_, _01992_);
  or (_02517_, _02516_, _02515_);
  and (_02518_, _01717_, _01986_);
  and (_02519_, _01689_, _01970_);
  or (_02520_, _02519_, _02518_);
  or (_02521_, _02520_, _02517_);
  or (_02522_, _02521_, _02514_);
  or (_02523_, _02522_, _02513_);
  and (_02524_, _01737_, _01967_);
  and (_02525_, _01709_, _01972_);
  and (_02526_, _01706_, _02005_);
  or (_02527_, _02526_, _02525_);
  or (_02528_, _02527_, _02524_);
  and (_02529_, _01701_, _02014_);
  and (_02530_, _01714_, _01979_);
  or (_02531_, _02530_, _02529_);
  and (_02532_, _01733_, _02012_);
  and (_02533_, _01680_, _02000_);
  and (_02534_, _01724_, _01974_);
  and (_02535_, _01721_, _01997_);
  or (_02536_, _02535_, _02534_);
  or (_02537_, _02536_, _02533_);
  or (_02538_, _02537_, _02532_);
  or (_02539_, _02538_, _02531_);
  or (_02540_, _02539_, _02528_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _02540_, _02523_);
  and (_02541_, _01661_, _02058_);
  and (_02542_, _01676_, _02025_);
  and (_02543_, _01685_, _02042_);
  or (_02544_, _02543_, _02542_);
  and (_02545_, _01689_, _02037_);
  and (_02546_, _01717_, _02048_);
  or (_02547_, _02546_, _02545_);
  or (_02548_, _02547_, _02544_);
  or (_02549_, _02548_, _02541_);
  and (_02550_, _01670_, _02068_);
  and (_02551_, _01665_, _02020_);
  or (_02552_, _02551_, _02550_);
  or (_02553_, _02552_, _02549_);
  and (_02554_, _01706_, _02061_);
  and (_02555_, _01709_, _02030_);
  and (_02556_, _01737_, _02022_);
  or (_02557_, _02556_, _02555_);
  or (_02558_, _02557_, _02554_);
  and (_02559_, _01701_, _02053_);
  and (_02560_, _01714_, _02056_);
  or (_02561_, _02560_, _02559_);
  and (_02562_, _01733_, _02070_);
  and (_02563_, _01680_, _02027_);
  and (_02564_, _01721_, _02045_);
  and (_02565_, _01724_, _02032_);
  or (_02566_, _02565_, _02564_);
  or (_02567_, _02566_, _02563_);
  or (_02568_, _02567_, _02562_);
  or (_02569_, _02568_, _02561_);
  or (_02570_, _02569_, _02558_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _02570_, _02553_);
  and (_02571_, _01661_, _02114_);
  and (_02572_, _01680_, _02090_);
  and (_02573_, _01676_, _02087_);
  or (_02574_, _02573_, _02572_);
  and (_02575_, _01717_, _02101_);
  and (_02576_, _01689_, _02080_);
  or (_02577_, _02576_, _02575_);
  or (_02578_, _02577_, _02574_);
  or (_02579_, _02578_, _02571_);
  and (_02580_, _01665_, _02075_);
  and (_02581_, _01670_, _02098_);
  or (_02582_, _02581_, _02580_);
  or (_02583_, _02582_, _02579_);
  and (_02584_, _01737_, _02077_);
  and (_02585_, _01701_, _02125_);
  and (_02586_, _01706_, _02117_);
  or (_02587_, _02586_, _02585_);
  or (_02588_, _02587_, _02584_);
  and (_02589_, _01709_, _02084_);
  and (_02590_, _01685_, _02123_);
  and (_02591_, _01724_, _02082_);
  and (_02592_, _01721_, _02104_);
  or (_02593_, _02592_, _02591_);
  or (_02594_, _02593_, _02590_);
  or (_02595_, _02594_, _02589_);
  and (_02596_, _01714_, _02112_);
  and (_02597_, _01733_, _02109_);
  or (_02598_, _02597_, _02596_);
  or (_02599_, _02598_, _02595_);
  or (_02600_, _02599_, _02588_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _02600_, _02583_);
  and (_02601_, _01661_, _02170_);
  and (_02602_, _01670_, _02154_);
  or (_02603_, _02602_, _02601_);
  and (_02604_, _01665_, _02135_);
  and (_02605_, _01685_, _02160_);
  and (_02606_, _01676_, _02146_);
  or (_02607_, _02606_, _02605_);
  and (_02608_, _01717_, _02178_);
  and (_02609_, _01680_, _02168_);
  or (_02610_, _02609_, _02608_);
  or (_02611_, _02610_, _02607_);
  or (_02612_, _02611_, _02604_);
  or (_02613_, _02612_, _02603_);
  and (_02614_, _01709_, _02137_);
  and (_02615_, _01714_, _02139_);
  and (_02616_, _01706_, _02173_);
  or (_02617_, _02616_, _02615_);
  or (_02618_, _02617_, _02614_);
  and (_02619_, _01733_, _02157_);
  and (_02620_, _01689_, _02130_);
  and (_02621_, _01724_, _02144_);
  and (_02622_, _01721_, _02165_);
  or (_02623_, _02622_, _02621_);
  or (_02624_, _02623_, _02620_);
  or (_02625_, _02624_, _02619_);
  and (_02626_, _01701_, _02180_);
  and (_02627_, _01737_, _02132_);
  or (_02628_, _02627_, _02626_);
  or (_02629_, _02628_, _02625_);
  or (_02630_, _02629_, _02618_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _02630_, _02613_);
  and (_02631_, _01670_, _02221_);
  and (_02632_, _01676_, _02224_);
  and (_02633_, _01717_, _02213_);
  or (_02634_, _02633_, _02632_);
  and (_02635_, _01680_, _02200_);
  and (_02636_, _01689_, _02190_);
  or (_02637_, _02636_, _02635_);
  or (_02638_, _02637_, _02634_);
  or (_02639_, _02638_, _02631_);
  and (_02640_, _01661_, _02226_);
  and (_02641_, _01665_, _02185_);
  or (_02642_, _02641_, _02640_);
  or (_02643_, _02642_, _02639_);
  and (_02644_, _01709_, _02193_);
  and (_02645_, _01733_, _02235_);
  and (_02646_, _01714_, _02202_);
  or (_02647_, _02646_, _02645_);
  or (_02648_, _02647_, _02644_);
  and (_02649_, _01737_, _02187_);
  and (_02650_, _01685_, _02210_);
  and (_02651_, _01721_, _02233_);
  and (_02652_, _01724_, _02196_);
  or (_02653_, _02652_, _02651_);
  or (_02654_, _02653_, _02650_);
  or (_02655_, _02654_, _02649_);
  and (_02656_, _01706_, _02228_);
  and (_02657_, _01701_, _02217_);
  or (_02658_, _02657_, _02656_);
  or (_02659_, _02658_, _02655_);
  or (_02661_, _02659_, _02648_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _02661_, _02643_);
  and (_02662_, _01661_, _01902_);
  and (_02663_, _01670_, _01879_);
  or (_02664_, _02663_, _02662_);
  and (_02665_, _01665_, _01890_);
  and (_02666_, _01685_, _01885_);
  and (_02667_, _01717_, _01900_);
  or (_02668_, _02667_, _02666_);
  and (_02669_, _01680_, _01888_);
  and (_02670_, _01676_, _01877_);
  or (_02671_, _02670_, _02669_);
  or (_02672_, _02671_, _02668_);
  or (_02673_, _02672_, _02665_);
  or (_02674_, _02673_, _02664_);
  and (_02675_, _01706_, _01859_);
  and (_02676_, _01733_, _01893_);
  and (_02677_, _01701_, _01856_);
  or (_02678_, _02677_, _02676_);
  or (_02679_, _02678_, _02675_);
  and (_02680_, _01714_, _01853_);
  and (_02681_, _01689_, _01869_);
  and (_02682_, _01724_, _01864_);
  and (_02683_, _01721_, _01875_);
  or (_02684_, _02683_, _02682_);
  or (_02685_, _02684_, _02681_);
  or (_02686_, _02685_, _02680_);
  and (_02687_, _01709_, _01862_);
  and (_02688_, _01737_, _01871_);
  or (_02689_, _02688_, _02687_);
  or (_02690_, _02689_, _02686_);
  or (_02691_, _02690_, _02679_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02691_, _02674_);
  and (_02692_, _01670_, _01937_);
  and (_02693_, _01661_, _01958_);
  or (_02694_, _02693_, _02692_);
  and (_02695_, _01665_, _01946_);
  and (_02696_, _01717_, _01956_);
  and (_02697_, _01689_, _01924_);
  or (_02698_, _02697_, _02696_);
  and (_02699_, _01680_, _01917_);
  and (_02700_, _01676_, _01933_);
  or (_02701_, _02700_, _02699_);
  or (_02702_, _02701_, _02698_);
  or (_02703_, _02702_, _02695_);
  or (_02704_, _02703_, _02694_);
  and (_02705_, _01709_, _01912_);
  and (_02706_, _01706_, _01914_);
  and (_02707_, _01737_, _01926_);
  or (_02708_, _02707_, _02706_);
  or (_02709_, _02708_, _02705_);
  and (_02710_, _01714_, _01909_);
  and (_02711_, _01685_, _01930_);
  and (_02712_, _01721_, _01941_);
  and (_02713_, _01724_, _01919_);
  or (_02714_, _02713_, _02712_);
  or (_02715_, _02714_, _02711_);
  or (_02716_, _02715_, _02710_);
  and (_02717_, _01733_, _01949_);
  and (_02718_, _01701_, _01944_);
  or (_02719_, _02718_, _02717_);
  or (_02720_, _02719_, _02716_);
  or (_02721_, _02720_, _02709_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02721_, _02704_);
  and (_02722_, _01661_, _01989_);
  and (_02723_, _01680_, _01977_);
  and (_02724_, _01685_, _01986_);
  or (_02725_, _02724_, _02723_);
  and (_02726_, _01676_, _01992_);
  and (_02727_, _01717_, _02014_);
  or (_02728_, _02727_, _02726_);
  or (_02729_, _02728_, _02725_);
  or (_02730_, _02729_, _02722_);
  and (_02731_, _01665_, _02002_);
  and (_02732_, _01670_, _01997_);
  or (_02733_, _02732_, _02731_);
  or (_02734_, _02733_, _02730_);
  and (_02735_, _01709_, _01974_);
  and (_02736_, _01701_, _01979_);
  and (_02737_, _01714_, _01967_);
  or (_02738_, _02737_, _02736_);
  or (_02739_, _02738_, _02735_);
  and (_02740_, _01733_, _02005_);
  and (_02741_, _01689_, _01965_);
  and (_02742_, _01721_, _02012_);
  and (_02743_, _01724_, _02000_);
  or (_02744_, _02743_, _02742_);
  or (_02745_, _02744_, _02741_);
  or (_02746_, _02745_, _02740_);
  and (_02747_, _01706_, _01972_);
  and (_02748_, _01737_, _01970_);
  or (_02749_, _02748_, _02747_);
  or (_02750_, _02749_, _02746_);
  or (_02751_, _02750_, _02739_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02751_, _02734_);
  and (_02752_, _01661_, _02068_);
  and (_02753_, _01717_, _02053_);
  and (_02754_, _01680_, _02025_);
  or (_02755_, _02754_, _02753_);
  and (_02756_, _01676_, _02042_);
  and (_02757_, _01689_, _02020_);
  or (_02758_, _02757_, _02756_);
  or (_02759_, _02758_, _02755_);
  or (_02760_, _02759_, _02752_);
  and (_02761_, _01665_, _02058_);
  and (_02762_, _01670_, _02045_);
  or (_02763_, _02762_, _02761_);
  or (_02764_, _02763_, _02760_);
  and (_02765_, _01709_, _02032_);
  and (_02766_, _01737_, _02037_);
  and (_02767_, _01706_, _02030_);
  or (_02768_, _02767_, _02766_);
  or (_02769_, _02768_, _02765_);
  and (_02770_, _01701_, _02056_);
  and (_02771_, _01685_, _02048_);
  and (_02772_, _01724_, _02027_);
  and (_02773_, _01721_, _02070_);
  or (_02774_, _02773_, _02772_);
  or (_02775_, _02774_, _02771_);
  or (_02776_, _02775_, _02770_);
  and (_02777_, _01714_, _02022_);
  and (_02778_, _01733_, _02061_);
  or (_02779_, _02778_, _02777_);
  or (_02780_, _02779_, _02776_);
  or (_02781_, _02780_, _02769_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02781_, _02764_);
  and (_02782_, _01661_, _02098_);
  and (_02783_, _01689_, _02075_);
  and (_02784_, _01676_, _02123_);
  or (_02785_, _02784_, _02783_);
  and (_02786_, _01680_, _02087_);
  and (_02787_, _01685_, _02101_);
  or (_02788_, _02787_, _02786_);
  or (_02789_, _02788_, _02785_);
  or (_02790_, _02789_, _02782_);
  and (_02791_, _01665_, _02114_);
  and (_02792_, _01670_, _02104_);
  or (_02793_, _02792_, _02791_);
  or (_02794_, _02793_, _02790_);
  and (_02795_, _01714_, _02077_);
  and (_02796_, _01733_, _02117_);
  and (_02797_, _01709_, _02082_);
  or (_02798_, _02797_, _02796_);
  or (_02799_, _02798_, _02795_);
  and (_02800_, _01737_, _02080_);
  and (_02801_, _01717_, _02125_);
  and (_02802_, _01721_, _02109_);
  and (_02803_, _01724_, _02090_);
  or (_02804_, _02803_, _02802_);
  or (_02805_, _02804_, _02801_);
  or (_02806_, _02805_, _02800_);
  and (_02807_, _01706_, _02084_);
  and (_02808_, _01701_, _02112_);
  or (_02809_, _02808_, _02807_);
  or (_02810_, _02809_, _02806_);
  or (_02811_, _02810_, _02799_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02811_, _02794_);
  and (_02812_, _01661_, _02154_);
  and (_02813_, _01689_, _02135_);
  and (_02814_, _01676_, _02160_);
  or (_02815_, _02814_, _02813_);
  and (_02816_, _01685_, _02178_);
  and (_02817_, _01717_, _02180_);
  or (_02818_, _02817_, _02816_);
  or (_02819_, _02818_, _02815_);
  or (_02820_, _02819_, _02812_);
  and (_02821_, _01665_, _02170_);
  and (_02822_, _01670_, _02165_);
  or (_02823_, _02822_, _02821_);
  or (_02824_, _02823_, _02820_);
  and (_02825_, _01714_, _02132_);
  and (_02826_, _01733_, _02173_);
  and (_02827_, _01706_, _02137_);
  or (_02828_, _02827_, _02826_);
  or (_02829_, _02828_, _02825_);
  and (_02830_, _01701_, _02139_);
  and (_02831_, _01680_, _02146_);
  and (_02832_, _01721_, _02157_);
  and (_02833_, _01724_, _02168_);
  or (_02834_, _02833_, _02832_);
  or (_02835_, _02834_, _02831_);
  or (_02836_, _02835_, _02830_);
  and (_02837_, _01709_, _02144_);
  and (_02838_, _01737_, _02130_);
  or (_02839_, _02838_, _02837_);
  or (_02840_, _02839_, _02836_);
  or (_02841_, _02840_, _02829_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02841_, _02824_);
  and (_02842_, _01661_, _02221_);
  and (_02843_, _01676_, _02210_);
  and (_02844_, _01685_, _02213_);
  or (_02845_, _02844_, _02843_);
  and (_02846_, _01680_, _02224_);
  and (_02847_, _01689_, _02185_);
  or (_02848_, _02847_, _02846_);
  or (_02849_, _02848_, _02845_);
  or (_02850_, _02849_, _02842_);
  and (_02851_, _01665_, _02226_);
  and (_02852_, _01670_, _02233_);
  or (_02853_, _02852_, _02851_);
  or (_02855_, _02853_, _02850_);
  and (_02856_, _01733_, _02228_);
  and (_02857_, _01709_, _02196_);
  and (_02858_, _01737_, _02190_);
  or (_02859_, _02858_, _02857_);
  or (_02860_, _02859_, _02856_);
  and (_02861_, _01706_, _02193_);
  and (_02862_, _01717_, _02217_);
  and (_02863_, _01721_, _02235_);
  and (_02864_, _01724_, _02200_);
  or (_02865_, _02864_, _02863_);
  or (_02866_, _02865_, _02862_);
  or (_02867_, _02866_, _02861_);
  and (_02868_, _01701_, _02202_);
  and (_02869_, _01714_, _02187_);
  or (_02870_, _02869_, _02868_);
  or (_02871_, _02870_, _02867_);
  or (_02872_, _02871_, _02860_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02872_, _02855_);
  nand (_02873_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_02874_, \oc8051_golden_model_1.PC [3]);
  or (_02875_, \oc8051_golden_model_1.PC [2], _02874_);
  or (_02876_, _02875_, _02873_);
  or (_02877_, _02876_, _42137_);
  not (_02878_, \oc8051_golden_model_1.PC [1]);
  or (_02879_, _02878_, \oc8051_golden_model_1.PC [0]);
  or (_02880_, _02879_, _02875_);
  or (_02881_, _02880_, _42096_);
  and (_02882_, _02881_, _02877_);
  not (_02883_, \oc8051_golden_model_1.PC [2]);
  or (_02884_, _02883_, \oc8051_golden_model_1.PC [3]);
  or (_02885_, _02884_, _02873_);
  or (_02886_, _02885_, _41973_);
  or (_02887_, _02884_, _02879_);
  or (_02888_, _02887_, _41932_);
  and (_02889_, _02888_, _02886_);
  and (_02890_, _02889_, _02882_);
  nand (_02891_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02892_, _02891_, _02873_);
  or (_02893_, _02892_, _42301_);
  or (_02894_, _02891_, _02879_);
  or (_02895_, _02894_, _42260_);
  and (_02896_, _02895_, _02893_);
  or (_02897_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02898_, _02897_, _02873_);
  or (_02899_, _02898_, _41809_);
  or (_02900_, _02897_, _02879_);
  or (_02901_, _02900_, _41758_);
  and (_02902_, _02901_, _02899_);
  and (_02903_, _02902_, _02896_);
  and (_02904_, _02903_, _02890_);
  not (_02905_, \oc8051_golden_model_1.PC [0]);
  or (_02906_, \oc8051_golden_model_1.PC [1], _02905_);
  or (_02907_, _02906_, _02891_);
  or (_02908_, _02907_, _42219_);
  or (_02909_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_02910_, _02909_, _02891_);
  or (_02911_, _02910_, _42178_);
  and (_02912_, _02911_, _02908_);
  or (_02913_, _02897_, _02909_);
  or (_02914_, _02913_, _41671_);
  or (_02915_, _02897_, _02906_);
  or (_02916_, _02915_, _41712_);
  and (_02917_, _02916_, _02914_);
  and (_02918_, _02917_, _02912_);
  or (_02919_, _02906_, _02875_);
  or (_02920_, _02919_, _42055_);
  or (_02921_, _02909_, _02875_);
  or (_02922_, _02921_, _42014_);
  and (_02923_, _02922_, _02920_);
  or (_02924_, _02906_, _02884_);
  or (_02925_, _02924_, _41891_);
  or (_02926_, _02909_, _02884_);
  or (_02927_, _02926_, _41850_);
  and (_02928_, _02927_, _02925_);
  and (_02929_, _02928_, _02923_);
  and (_02930_, _02929_, _02918_);
  nand (_02931_, _02930_, _02904_);
  or (_02932_, _02876_, _42142_);
  or (_02933_, _02880_, _42101_);
  and (_02934_, _02933_, _02932_);
  or (_02935_, _02885_, _41978_);
  or (_02936_, _02887_, _41937_);
  and (_02937_, _02936_, _02935_);
  and (_02938_, _02937_, _02934_);
  or (_02939_, _02892_, _42306_);
  or (_02940_, _02894_, _42265_);
  and (_02941_, _02940_, _02939_);
  or (_02942_, _02898_, _41814_);
  or (_02943_, _02900_, _41765_);
  and (_02944_, _02943_, _02942_);
  and (_02945_, _02944_, _02941_);
  and (_02946_, _02945_, _02938_);
  or (_02947_, _02907_, _42224_);
  or (_02948_, _02910_, _42183_);
  and (_02949_, _02948_, _02947_);
  or (_02950_, _02913_, _41676_);
  or (_02951_, _02915_, _41717_);
  and (_02952_, _02951_, _02950_);
  and (_02953_, _02952_, _02949_);
  or (_02954_, _02919_, _42060_);
  or (_02955_, _02921_, _42019_);
  and (_02956_, _02955_, _02954_);
  or (_02957_, _02924_, _41896_);
  or (_02958_, _02926_, _41855_);
  and (_02959_, _02958_, _02957_);
  and (_02960_, _02959_, _02956_);
  and (_02961_, _02960_, _02953_);
  nand (_02962_, _02961_, _02946_);
  or (_02963_, _02962_, _02931_);
  or (_02964_, _02876_, _42127_);
  or (_02965_, _02880_, _42086_);
  and (_02966_, _02965_, _02964_);
  or (_02967_, _02885_, _41963_);
  or (_02968_, _02887_, _41922_);
  and (_02969_, _02968_, _02967_);
  and (_02970_, _02969_, _02966_);
  or (_02971_, _02892_, _42291_);
  or (_02972_, _02894_, _42250_);
  and (_02973_, _02972_, _02971_);
  or (_02974_, _02898_, _41791_);
  or (_02975_, _02900_, _41743_);
  and (_02976_, _02975_, _02974_);
  and (_02977_, _02976_, _02973_);
  and (_02978_, _02977_, _02970_);
  or (_02979_, _02907_, _42209_);
  or (_02980_, _02910_, _42168_);
  and (_02981_, _02980_, _02979_);
  or (_02982_, _02913_, _41661_);
  or (_02983_, _02915_, _41702_);
  and (_02984_, _02983_, _02982_);
  and (_02985_, _02984_, _02981_);
  or (_02986_, _02919_, _42045_);
  or (_02987_, _02921_, _42004_);
  and (_02988_, _02987_, _02986_);
  or (_02989_, _02924_, _41881_);
  or (_02990_, _02926_, _41840_);
  and (_02991_, _02990_, _02989_);
  and (_02992_, _02991_, _02988_);
  and (_02993_, _02992_, _02985_);
  and (_02994_, _02993_, _02978_);
  or (_02995_, _02876_, _42132_);
  or (_02996_, _02880_, _42091_);
  and (_02997_, _02996_, _02995_);
  or (_02998_, _02885_, _41968_);
  or (_02999_, _02887_, _41927_);
  and (_03000_, _02999_, _02998_);
  and (_03001_, _03000_, _02997_);
  or (_03002_, _02892_, _42296_);
  or (_03003_, _02894_, _42255_);
  and (_03004_, _03003_, _03002_);
  or (_03005_, _02898_, _41801_);
  or (_03006_, _02900_, _41749_);
  and (_03007_, _03006_, _03005_);
  and (_03008_, _03007_, _03004_);
  and (_03009_, _03008_, _03001_);
  or (_03010_, _02907_, _42214_);
  or (_03011_, _02910_, _42173_);
  and (_03012_, _03011_, _03010_);
  or (_03013_, _02913_, _41666_);
  or (_03015_, _02915_, _41707_);
  and (_03016_, _03015_, _03013_);
  and (_03017_, _03016_, _03012_);
  or (_03018_, _02919_, _42050_);
  or (_03019_, _02921_, _42009_);
  and (_03020_, _03019_, _03018_);
  or (_03021_, _02924_, _41886_);
  or (_03022_, _02926_, _41845_);
  and (_03023_, _03022_, _03021_);
  and (_03024_, _03023_, _03020_);
  and (_03026_, _03024_, _03017_);
  nand (_03027_, _03026_, _03009_);
  or (_03028_, _03027_, _02994_);
  or (_03029_, _03028_, _02963_);
  not (_03030_, _03029_);
  or (_03031_, _02876_, _42147_);
  or (_03032_, _02880_, _42106_);
  and (_03033_, _03032_, _03031_);
  or (_03034_, _02885_, _41983_);
  or (_03035_, _02887_, _41942_);
  and (_03036_, _03035_, _03034_);
  and (_03037_, _03036_, _03033_);
  or (_03038_, _02892_, _42311_);
  or (_03039_, _02894_, _42270_);
  and (_03040_, _03039_, _03038_);
  or (_03041_, _02898_, _41819_);
  or (_03042_, _02900_, _41770_);
  and (_03043_, _03042_, _03041_);
  and (_03044_, _03043_, _03040_);
  and (_03045_, _03044_, _03037_);
  or (_03047_, _02907_, _42229_);
  or (_03048_, _02910_, _42188_);
  and (_03049_, _03048_, _03047_);
  or (_03050_, _02913_, _41681_);
  or (_03051_, _02915_, _41722_);
  and (_03052_, _03051_, _03050_);
  and (_03053_, _03052_, _03049_);
  or (_03054_, _02919_, _42065_);
  or (_03055_, _02921_, _42024_);
  and (_03056_, _03055_, _03054_);
  or (_03058_, _02924_, _41901_);
  or (_03059_, _02926_, _41860_);
  and (_03060_, _03059_, _03058_);
  and (_03061_, _03060_, _03056_);
  and (_03062_, _03061_, _03053_);
  nand (_03063_, _03062_, _03045_);
  or (_03064_, _02876_, _42152_);
  or (_03065_, _02880_, _42111_);
  and (_03066_, _03065_, _03064_);
  or (_03067_, _02885_, _41988_);
  or (_03069_, _02887_, _41947_);
  and (_03070_, _03069_, _03067_);
  and (_03071_, _03070_, _03066_);
  or (_03072_, _02892_, _42316_);
  or (_03073_, _02894_, _42275_);
  and (_03074_, _03073_, _03072_);
  or (_03075_, _02898_, _41824_);
  or (_03076_, _02900_, _41775_);
  and (_03077_, _03076_, _03075_);
  and (_03078_, _03077_, _03074_);
  and (_03079_, _03078_, _03071_);
  or (_03080_, _02907_, _42234_);
  or (_03081_, _02910_, _42193_);
  and (_03082_, _03081_, _03080_);
  or (_03083_, _02913_, _41686_);
  or (_03084_, _02915_, _41727_);
  and (_03085_, _03084_, _03083_);
  and (_03086_, _03085_, _03082_);
  or (_03087_, _02919_, _42070_);
  or (_03088_, _02921_, _42029_);
  and (_03090_, _03088_, _03087_);
  or (_03091_, _02924_, _41906_);
  or (_03092_, _02926_, _41865_);
  and (_03093_, _03092_, _03091_);
  and (_03094_, _03093_, _03090_);
  and (_03095_, _03094_, _03086_);
  nand (_03096_, _03095_, _03079_);
  or (_03097_, _03096_, _03063_);
  or (_03098_, _02876_, _42157_);
  or (_03099_, _02880_, _42116_);
  and (_03101_, _03099_, _03098_);
  or (_03102_, _02885_, _41993_);
  or (_03103_, _02887_, _41952_);
  and (_03104_, _03103_, _03102_);
  and (_03105_, _03104_, _03101_);
  or (_03106_, _02892_, _42321_);
  or (_03107_, _02894_, _42280_);
  and (_03108_, _03107_, _03106_);
  or (_03109_, _02898_, _41829_);
  or (_03110_, _02900_, _41780_);
  and (_03112_, _03110_, _03109_);
  and (_03113_, _03112_, _03108_);
  and (_03114_, _03113_, _03105_);
  or (_03115_, _02907_, _42239_);
  or (_03116_, _02910_, _42198_);
  and (_03117_, _03116_, _03115_);
  or (_03118_, _02913_, _41691_);
  or (_03119_, _02915_, _41732_);
  and (_03120_, _03119_, _03118_);
  and (_03121_, _03120_, _03117_);
  or (_03123_, _02919_, _42075_);
  or (_03124_, _02921_, _42034_);
  and (_03125_, _03124_, _03123_);
  or (_03126_, _02924_, _41911_);
  or (_03127_, _02926_, _41870_);
  and (_03128_, _03127_, _03126_);
  and (_03129_, _03128_, _03125_);
  and (_03130_, _03129_, _03121_);
  nand (_03131_, _03130_, _03114_);
  or (_03132_, _02876_, _42122_);
  or (_03134_, _02880_, _42081_);
  and (_03135_, _03134_, _03132_);
  or (_03136_, _02885_, _41958_);
  or (_03137_, _02887_, _41917_);
  and (_03138_, _03137_, _03136_);
  and (_03139_, _03138_, _03135_);
  or (_03140_, _02892_, _42286_);
  or (_03141_, _02894_, _42245_);
  and (_03142_, _03141_, _03140_);
  or (_03143_, _02898_, _41786_);
  or (_03145_, _02900_, _41738_);
  and (_03146_, _03145_, _03143_);
  and (_03147_, _03146_, _03142_);
  and (_03148_, _03147_, _03139_);
  or (_03149_, _02907_, _42204_);
  or (_03150_, _02910_, _42163_);
  and (_03151_, _03150_, _03149_);
  or (_03152_, _02913_, _41656_);
  or (_03153_, _02915_, _41697_);
  and (_03154_, _03153_, _03152_);
  and (_03156_, _03154_, _03151_);
  or (_03157_, _02919_, _42040_);
  or (_03158_, _02921_, _41999_);
  and (_03159_, _03158_, _03157_);
  or (_03160_, _02924_, _41876_);
  or (_03161_, _02926_, _41835_);
  and (_03162_, _03161_, _03160_);
  and (_03163_, _03162_, _03159_);
  and (_03164_, _03163_, _03156_);
  and (_03165_, _03164_, _03148_);
  or (_03167_, _03165_, _03131_);
  nor (_03168_, _03167_, _03097_);
  and (_03169_, _03168_, _03030_);
  not (_03170_, _03169_);
  and (_03171_, _03165_, _03131_);
  and (_03172_, _03062_, _03045_);
  and (_03173_, _03095_, _03079_);
  or (_03174_, _03173_, _03172_);
  not (_03175_, _03174_);
  and (_03176_, _03175_, _03171_);
  and (_03178_, _03176_, _03030_);
  or (_03179_, _03173_, _03063_);
  not (_03180_, _03179_);
  and (_03181_, _03180_, _03171_);
  and (_03182_, _03181_, _03030_);
  nor (_03183_, _03182_, _03178_);
  and (_03184_, _03183_, _03170_);
  and (_03185_, _03130_, _03114_);
  and (_03186_, _03165_, _03185_);
  and (_03187_, _03175_, _03186_);
  and (_03188_, _03187_, _03030_);
  or (_03189_, _03096_, _03172_);
  not (_03190_, _03189_);
  and (_03191_, _03171_, _03190_);
  and (_03192_, _03191_, _03030_);
  nor (_03193_, _03192_, _03188_);
  not (_03194_, _03097_);
  and (_03195_, _03194_, _03186_);
  and (_03196_, _03195_, _03030_);
  and (_03197_, _03190_, _03186_);
  and (_03198_, _03030_, _03197_);
  nor (_03199_, _03198_, _03196_);
  and (_03200_, _03171_, _03194_);
  and (_03201_, _03200_, _03030_);
  and (_03202_, _03180_, _03186_);
  and (_03203_, _03202_, _03030_);
  nor (_03204_, _03203_, _03201_);
  and (_03205_, _03204_, _03199_);
  and (_03206_, _03205_, _03193_);
  and (_03207_, _03206_, _03184_);
  and (_03208_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03209_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03210_, _03209_, _03208_);
  or (_03211_, _03210_, _03207_);
  not (_03212_, _03168_);
  not (_03213_, _03027_);
  or (_03214_, _03213_, _02994_);
  or (_03215_, _03214_, _02963_);
  nor (_03216_, _03215_, _03212_);
  not (_03217_, _03216_);
  not (_03218_, _03028_);
  not (_03219_, _02962_);
  and (_03220_, _03219_, _02931_);
  and (_03221_, _03220_, _03218_);
  and (_03222_, _03221_, _03168_);
  nor (_03223_, _03167_, _03189_);
  and (_03224_, _03223_, _03030_);
  nor (_03225_, _03224_, _03222_);
  or (_03226_, _03167_, _03174_);
  or (_03227_, _03226_, _03029_);
  or (_03228_, _03165_, _03185_);
  or (_03229_, _03228_, _03189_);
  or (_03230_, _03229_, _03029_);
  and (_03231_, _03230_, _03227_);
  or (_03232_, _03228_, _03097_);
  or (_03233_, _03232_, _03029_);
  or (_03234_, _03228_, _03179_);
  or (_03235_, _03234_, _03029_);
  and (_03236_, _03235_, _03233_);
  or (_03237_, _03167_, _03179_);
  or (_03238_, _03237_, _03029_);
  or (_03239_, _03228_, _03174_);
  or (_03240_, _03239_, _03029_);
  and (_03241_, _03240_, _03238_);
  and (_03242_, _03241_, _03236_);
  and (_03243_, _03242_, _03231_);
  and (_03244_, _03243_, _03225_);
  not (_03245_, _03210_);
  or (_03246_, _03245_, _03244_);
  not (_03247_, _03223_);
  or (_03248_, _03247_, _03215_);
  and (_03249_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_03250_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03251_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_03252_, _03251_, _03249_);
  and (_03253_, _03252_, _03250_);
  nor (_03254_, _03253_, _03249_);
  and (_03255_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_03256_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_03257_, _03256_, _03255_);
  not (_03258_, _03257_);
  nor (_03259_, _03258_, _03254_);
  and (_03260_, _03258_, _03254_);
  nor (_03261_, _03260_, _03259_);
  not (_03262_, _03261_);
  or (_03263_, _03262_, _03248_);
  nor (_03264_, _02873_, _02883_);
  and (_03265_, _02873_, _02883_);
  nor (_03266_, _03265_, _03264_);
  and (_03267_, _03266_, _03248_);
  nand (_03269_, _03267_, _03243_);
  nand (_03270_, _03269_, _03263_);
  nand (_03271_, _03270_, _03225_);
  nand (_03272_, _03271_, _03246_);
  nand (_03273_, _03272_, _03217_);
  not (_03274_, \oc8051_golden_model_1.ACC [1]);
  and (_03275_, _02906_, _02879_);
  nor (_03276_, _03275_, _03274_);
  and (_03277_, \oc8051_golden_model_1.ACC [0], _02905_);
  and (_03278_, _03275_, _03274_);
  nor (_03279_, _03278_, _03276_);
  and (_03280_, _03279_, _03277_);
  nor (_03281_, _03280_, _03276_);
  and (_03282_, _03266_, \oc8051_golden_model_1.ACC [2]);
  nor (_03283_, _03266_, \oc8051_golden_model_1.ACC [2]);
  nor (_03284_, _03283_, _03282_);
  not (_03285_, _03284_);
  nor (_03286_, _03285_, _03281_);
  and (_03287_, _03285_, _03281_);
  nor (_03288_, _03287_, _03286_);
  and (_03289_, _03288_, _03216_);
  not (_03290_, _03289_);
  and (_03291_, _03290_, _03207_);
  nand (_03292_, _03291_, _03273_);
  nand (_03293_, _03292_, _03211_);
  and (_03294_, _03244_, _03207_);
  nor (_03295_, _02891_, _02878_);
  nor (_03296_, _03208_, \oc8051_golden_model_1.PC [3]);
  nor (_03297_, _03296_, _03295_);
  or (_03298_, _03297_, _03294_);
  and (_03299_, _03225_, _03217_);
  nor (_03300_, _03259_, _03255_);
  and (_03301_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03302_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03303_, _03302_, _03301_);
  not (_03304_, _03303_);
  nor (_03305_, _03304_, _03300_);
  and (_03306_, _03304_, _03300_);
  nor (_03307_, _03306_, _03305_);
  or (_03308_, _03307_, _03248_);
  not (_03309_, _02885_);
  nor (_03310_, _03264_, _02874_);
  nor (_03311_, _03310_, _03309_);
  and (_03312_, _03248_, _03311_);
  nand (_03313_, _03312_, _03243_);
  nand (_03314_, _03313_, _03308_);
  and (_03315_, _03314_, _03299_);
  nor (_03316_, _03286_, _03282_);
  nor (_03317_, _03311_, \oc8051_golden_model_1.ACC [3]);
  and (_03318_, _03311_, \oc8051_golden_model_1.ACC [3]);
  nor (_03319_, _03318_, _03317_);
  and (_03320_, _03319_, _03316_);
  nor (_03321_, _03319_, _03316_);
  nor (_03322_, _03321_, _03320_);
  nor (_03323_, _03322_, _03217_);
  or (_03324_, _03323_, _03315_);
  nand (_03325_, _03324_, _03207_);
  and (_03326_, _03325_, _03298_);
  or (_03327_, _03326_, _03293_);
  nor (_03328_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03329_, _03328_, _03250_);
  or (_03330_, _03329_, _03248_);
  and (_03331_, _03248_, \oc8051_golden_model_1.PC [0]);
  nand (_03332_, _03331_, _03243_);
  nand (_03333_, _03332_, _03330_);
  and (_03334_, _03333_, _03299_);
  not (_03335_, \oc8051_golden_model_1.ACC [0]);
  and (_03336_, _03335_, \oc8051_golden_model_1.PC [0]);
  nor (_03337_, _03336_, _03277_);
  nor (_03338_, _03337_, _03217_);
  or (_03339_, _03338_, _03334_);
  nand (_03340_, _03339_, _03207_);
  or (_03341_, _03294_, \oc8051_golden_model_1.PC [0]);
  and (_03342_, _03341_, _03340_);
  or (_03343_, _03294_, _02878_);
  nor (_03344_, _03252_, _03250_);
  nor (_03345_, _03344_, _03253_);
  or (_03346_, _03345_, _03248_);
  and (_03347_, _03275_, _03248_);
  nand (_03348_, _03347_, _03243_);
  nand (_03349_, _03348_, _03346_);
  and (_03350_, _03349_, _03299_);
  nor (_03351_, _03279_, _03277_);
  nor (_03352_, _03351_, _03280_);
  nor (_03353_, _03352_, _03217_);
  or (_03354_, _03353_, _03350_);
  nand (_03355_, _03354_, _03207_);
  nand (_03356_, _03355_, _03343_);
  or (_03357_, _03356_, _03342_);
  or (_03358_, _03357_, _03327_);
  nor (_03359_, _03358_, _41927_);
  nand (_03360_, _03341_, _03340_);
  and (_03361_, _03355_, _03343_);
  or (_03362_, _03361_, _03360_);
  or (_03363_, _03362_, _03327_);
  nor (_03364_, _03363_, _41886_);
  nor (_03365_, _03364_, _03359_);
  or (_03366_, _03356_, _03360_);
  and (_03367_, _03292_, _03211_);
  nand (_03368_, _03325_, _03298_);
  or (_03369_, _03368_, _03367_);
  or (_03370_, _03369_, _03366_);
  nor (_03371_, _03370_, _42132_);
  or (_03372_, _03326_, _03367_);
  or (_03373_, _03361_, _03342_);
  or (_03374_, _03373_, _03372_);
  nor (_03375_, _03374_, _41666_);
  nor (_03376_, _03375_, _03371_);
  and (_03377_, _03376_, _03365_);
  or (_03378_, _03369_, _03357_);
  nor (_03379_, _03378_, _42091_);
  or (_03380_, _03369_, _03362_);
  nor (_03381_, _03380_, _42050_);
  nor (_03382_, _03381_, _03379_);
  or (_03383_, _03368_, _03293_);
  or (_03384_, _03383_, _03357_);
  nor (_03385_, _03384_, _42255_);
  or (_03386_, _03372_, _03366_);
  nor (_03387_, _03386_, _41801_);
  nor (_03388_, _03387_, _03385_);
  and (_03389_, _03388_, _03382_);
  and (_03390_, _03389_, _03377_);
  or (_03391_, _03383_, _03366_);
  nor (_03392_, _03391_, _42296_);
  or (_03393_, _03373_, _03383_);
  nor (_03394_, _03393_, _42173_);
  nor (_03395_, _03394_, _03392_);
  or (_03396_, _03327_, _03366_);
  nor (_03397_, _03396_, _41968_);
  or (_03398_, _03373_, _03327_);
  nor (_03399_, _03398_, _41845_);
  nor (_03400_, _03399_, _03397_);
  and (_03401_, _03400_, _03395_);
  or (_03402_, _03369_, _03373_);
  nor (_03403_, _03402_, _42009_);
  or (_03404_, _03357_, _03372_);
  nor (_03405_, _03404_, _41749_);
  nor (_03406_, _03405_, _03403_);
  or (_03407_, _03362_, _03383_);
  nor (_03408_, _03407_, _42214_);
  or (_03409_, _03362_, _03372_);
  nor (_03410_, _03409_, _41707_);
  nor (_03411_, _03410_, _03408_);
  and (_03412_, _03411_, _03406_);
  and (_03413_, _03412_, _03401_);
  and (_03414_, _03413_, _03390_);
  not (_03415_, _03414_);
  or (_03416_, _03396_, _41958_);
  or (_03417_, _03386_, _41786_);
  and (_03418_, _03417_, _03416_);
  or (_03419_, _03384_, _42245_);
  or (_03420_, _03393_, _42163_);
  and (_03421_, _03420_, _03419_);
  and (_03422_, _03421_, _03418_);
  or (_03423_, _03358_, _41917_);
  or (_03424_, _03363_, _41876_);
  and (_03425_, _03424_, _03423_);
  or (_03426_, _03374_, _41656_);
  or (_03427_, _03404_, _41738_);
  and (_03428_, _03427_, _03426_);
  and (_03429_, _03428_, _03425_);
  and (_03430_, _03429_, _03422_);
  or (_03431_, _03378_, _42081_);
  or (_03432_, _03402_, _41999_);
  and (_03433_, _03432_, _03431_);
  or (_03434_, _03391_, _42286_);
  or (_03435_, _03407_, _42204_);
  and (_03436_, _03435_, _03434_);
  and (_03437_, _03436_, _03433_);
  or (_03438_, _03398_, _41835_);
  or (_03439_, _03409_, _41697_);
  and (_03440_, _03439_, _03438_);
  or (_03441_, _03370_, _42122_);
  or (_03442_, _03380_, _42040_);
  and (_03443_, _03442_, _03441_);
  and (_03444_, _03443_, _03440_);
  and (_03445_, _03444_, _03437_);
  and (_03446_, _03445_, _03430_);
  and (_03447_, _03221_, _03195_);
  and (_03448_, _03447_, _03446_);
  and (_03449_, _03448_, _03415_);
  not (_03450_, _02963_);
  and (_03451_, _03213_, _02994_);
  and (_03452_, _03451_, _03450_);
  and (_03453_, _03452_, _03197_);
  not (_03454_, _03446_);
  nor (_03455_, _03358_, _41942_);
  nor (_03456_, _03363_, _41901_);
  nor (_03457_, _03456_, _03455_);
  nor (_03458_, _03391_, _42311_);
  nor (_03459_, _03370_, _42147_);
  nor (_03460_, _03459_, _03458_);
  and (_03461_, _03460_, _03457_);
  nor (_03462_, _03384_, _42270_);
  nor (_03463_, _03407_, _42229_);
  nor (_03464_, _03463_, _03462_);
  nor (_03465_, _03378_, _42106_);
  nor (_03466_, _03402_, _42024_);
  nor (_03467_, _03466_, _03465_);
  and (_03468_, _03467_, _03464_);
  and (_03470_, _03468_, _03461_);
  nor (_03471_, _03374_, _41681_);
  nor (_03472_, _03404_, _41770_);
  nor (_03473_, _03472_, _03471_);
  nor (_03474_, _03396_, _41983_);
  nor (_03475_, _03398_, _41860_);
  nor (_03476_, _03475_, _03474_);
  and (_03477_, _03476_, _03473_);
  nor (_03478_, _03393_, _42188_);
  nor (_03479_, _03380_, _42065_);
  nor (_03480_, _03479_, _03478_);
  nor (_03481_, _03386_, _41819_);
  nor (_03482_, _03409_, _41722_);
  nor (_03483_, _03482_, _03481_);
  and (_03484_, _03483_, _03480_);
  and (_03485_, _03484_, _03477_);
  and (_03486_, _03485_, _03470_);
  nor (_03487_, _03486_, _03454_);
  and (_03488_, _03487_, _03453_);
  and (_03489_, _02962_, _02931_);
  and (_03490_, _03489_, _03213_);
  and (_03491_, _03490_, _03197_);
  not (_03492_, _03491_);
  nor (_03493_, _03219_, _02931_);
  and (_03494_, _03493_, _03213_);
  and (_03495_, _03494_, _03197_);
  not (_03496_, \oc8051_golden_model_1.SP [1]);
  and (_03497_, _03496_, \oc8051_golden_model_1.SP [0]);
  not (_03498_, \oc8051_golden_model_1.SP [0]);
  and (_03499_, \oc8051_golden_model_1.SP [1], _03498_);
  nor (_03500_, _03499_, _03497_);
  not (_03501_, _03500_);
  and (_03502_, _03501_, _03188_);
  and (_03503_, _03027_, _02994_);
  and (_03504_, _03503_, _03450_);
  and (_03505_, _03504_, _03223_);
  and (_03506_, _03487_, _03505_);
  not (_03507_, _03232_);
  and (_03508_, _03507_, _03452_);
  and (_03509_, _03501_, _03508_);
  not (_03510_, _03508_);
  nand (_03511_, _03220_, _03027_);
  nor (_03512_, _03511_, _03239_);
  not (_03513_, _03240_);
  not (_03514_, _03447_);
  and (_03515_, _03504_, _03202_);
  not (_03516_, _03515_);
  and (_03517_, _03221_, _03202_);
  not (_03518_, _03517_);
  nor (_03519_, _03396_, _41993_);
  nor (_03520_, _03409_, _41732_);
  nor (_03521_, _03520_, _03519_);
  nor (_03522_, _03402_, _42034_);
  nor (_03523_, _03386_, _41829_);
  nor (_03524_, _03523_, _03522_);
  and (_03525_, _03524_, _03521_);
  nor (_03526_, _03370_, _42157_);
  nor (_03527_, _03374_, _41691_);
  nor (_03528_, _03527_, _03526_);
  nor (_03529_, _03407_, _42239_);
  nor (_03530_, _03393_, _42198_);
  nor (_03531_, _03530_, _03529_);
  and (_03532_, _03531_, _03528_);
  and (_03533_, _03532_, _03525_);
  nor (_03534_, _03384_, _42280_);
  nor (_03535_, _03404_, _41780_);
  nor (_03536_, _03535_, _03534_);
  nor (_03537_, _03380_, _42075_);
  nor (_03538_, _03358_, _41952_);
  nor (_03539_, _03538_, _03537_);
  and (_03540_, _03539_, _03536_);
  nor (_03541_, _03378_, _42116_);
  nor (_03542_, _03398_, _41870_);
  nor (_03543_, _03542_, _03541_);
  nor (_03544_, _03391_, _42321_);
  nor (_03545_, _03363_, _41911_);
  nor (_03546_, _03545_, _03544_);
  and (_03547_, _03546_, _03543_);
  and (_03548_, _03547_, _03540_);
  and (_03549_, _03548_, _03533_);
  nor (_03550_, _03549_, _03454_);
  or (_03551_, _03391_, _42306_);
  or (_03552_, _03402_, _42019_);
  and (_03553_, _03552_, _03551_);
  or (_03554_, _03378_, _42101_);
  or (_03555_, _03386_, _41814_);
  and (_03556_, _03555_, _03554_);
  and (_03557_, _03556_, _03553_);
  or (_03558_, _03384_, _42265_);
  or (_03559_, _03407_, _42224_);
  and (_03560_, _03559_, _03558_);
  or (_03561_, _03396_, _41978_);
  or (_03562_, _03398_, _41855_);
  and (_03563_, _03562_, _03561_);
  and (_03564_, _03563_, _03560_);
  and (_03565_, _03564_, _03557_);
  or (_03566_, _03363_, _41896_);
  or (_03567_, _03404_, _41765_);
  and (_03568_, _03567_, _03566_);
  or (_03569_, _03374_, _41676_);
  or (_03570_, _03409_, _41717_);
  and (_03571_, _03570_, _03569_);
  and (_03572_, _03571_, _03568_);
  or (_03573_, _03393_, _42183_);
  or (_03574_, _03358_, _41937_);
  and (_03575_, _03574_, _03573_);
  or (_03576_, _03370_, _42142_);
  or (_03577_, _03380_, _42060_);
  and (_03578_, _03577_, _03576_);
  and (_03579_, _03578_, _03575_);
  and (_03580_, _03579_, _03572_);
  and (_03581_, _03580_, _03565_);
  nor (_03582_, _03581_, _03446_);
  nor (_03583_, _03582_, _03550_);
  and (_03584_, _03504_, _03176_);
  and (_03585_, _03504_, _03168_);
  nor (_03586_, _03585_, _03584_);
  not (_03587_, _03586_);
  and (_03588_, _03587_, _03583_);
  not (_03589_, _03222_);
  not (_03590_, _03226_);
  and (_03591_, _03489_, _03503_);
  and (_03592_, _03489_, _03218_);
  or (_03593_, _03592_, _03591_);
  and (_03594_, _03593_, _03590_);
  and (_03595_, _03489_, _03451_);
  nor (_03596_, _03493_, _03595_);
  nor (_03597_, _03596_, _03226_);
  nor (_03598_, _03597_, _03594_);
  not (_03599_, _03215_);
  and (_03600_, _03599_, _03181_);
  and (_03601_, _03221_, _03176_);
  nor (_03602_, _03601_, _03600_);
  and (_03603_, _03220_, _03451_);
  and (_03604_, _03603_, _03590_);
  and (_03605_, _03503_, _03220_);
  and (_03606_, _03605_, _03590_);
  nor (_03607_, _03606_, _03604_);
  and (_03608_, _03607_, _03602_);
  not (_03609_, _03229_);
  and (_03610_, _03609_, _03221_);
  not (_03611_, _03214_);
  and (_03612_, _03489_, _03611_);
  and (_03613_, _03612_, _03590_);
  nor (_03614_, _03613_, _03610_);
  and (_03615_, _03590_, _03221_);
  and (_03616_, _03220_, _03611_);
  and (_03617_, _03616_, _03590_);
  nor (_03618_, _03617_, _03615_);
  and (_03619_, _03618_, _03614_);
  and (_03620_, _03619_, _03608_);
  and (_03621_, _03187_, _03452_);
  and (_03622_, _03599_, _03191_);
  nor (_03623_, _03622_, _03621_);
  and (_03624_, _03599_, _03200_);
  and (_03625_, _03223_, _03452_);
  nor (_03626_, _03625_, _03624_);
  and (_03627_, _03626_, _03623_);
  and (_03628_, _03202_, _03452_);
  and (_03629_, _03504_, _03197_);
  nor (_03630_, _03629_, _03628_);
  and (_03631_, _03504_, _03195_);
  nor (_03632_, _03631_, _03453_);
  and (_03633_, _03632_, _03630_);
  and (_03634_, _03633_, _03627_);
  and (_03635_, _03634_, _03620_);
  and (_03636_, _03635_, _03598_);
  and (_03637_, _03636_, _02905_);
  nor (_03638_, _03637_, \oc8051_golden_model_1.PC [1]);
  and (_03639_, _03637_, \oc8051_golden_model_1.PC [1]);
  nor (_03640_, _03639_, _03638_);
  nor (_03641_, _03636_, _02905_);
  nor (_03642_, _03641_, _03637_);
  nor (_03643_, _03642_, _03640_);
  nor (_03644_, _03636_, _03245_);
  and (_03645_, _03636_, _03266_);
  nor (_03646_, _03645_, _03644_);
  not (_03647_, _03646_);
  not (_03648_, _03297_);
  nor (_03649_, _03636_, _03648_);
  not (_03650_, _03311_);
  and (_03651_, _03636_, _03650_);
  nor (_03652_, _03651_, _03649_);
  and (_03653_, _03652_, _03647_);
  and (_03654_, _03653_, _03643_);
  and (_03655_, _03654_, _02025_);
  and (_03656_, _03652_, _03646_);
  and (_03657_, _03656_, _03643_);
  and (_03658_, _03657_, _02056_);
  nor (_03659_, _03658_, _03655_);
  nor (_03660_, _03652_, _03646_);
  and (_03661_, _03642_, _03640_);
  and (_03662_, _03661_, _03660_);
  and (_03663_, _03662_, _02070_);
  nor (_03664_, _03652_, _03647_);
  and (_03665_, _03664_, _03661_);
  and (_03666_, _03665_, _02027_);
  nor (_03667_, _03666_, _03663_);
  and (_03668_, _03667_, _03659_);
  not (_03669_, _03642_);
  nor (_03671_, _03669_, _03640_);
  and (_03672_, _03671_, _03653_);
  and (_03673_, _03672_, _02042_);
  and (_03674_, _03669_, _03640_);
  and (_03675_, _03674_, _03653_);
  and (_03676_, _03675_, _02048_);
  nor (_03677_, _03676_, _03673_);
  and (_03678_, _03661_, _03653_);
  and (_03679_, _03678_, _02053_);
  and (_03680_, _03661_, _03656_);
  and (_03681_, _03680_, _02020_);
  nor (_03682_, _03681_, _03679_);
  and (_03683_, _03682_, _03677_);
  and (_03684_, _03683_, _03668_);
  and (_03685_, _03660_, _03643_);
  and (_03686_, _03685_, _02058_);
  and (_03687_, _03671_, _03660_);
  and (_03688_, _03687_, _02068_);
  nor (_03689_, _03688_, _03686_);
  and (_03690_, _03674_, _03660_);
  and (_03691_, _03690_, _02045_);
  and (_03692_, _03664_, _03643_);
  and (_03693_, _03692_, _02061_);
  nor (_03694_, _03693_, _03691_);
  and (_03695_, _03694_, _03689_);
  and (_03696_, _03671_, _03664_);
  and (_03697_, _03696_, _02030_);
  and (_03698_, _03674_, _03664_);
  and (_03699_, _03698_, _02032_);
  nor (_03700_, _03699_, _03697_);
  and (_03701_, _03671_, _03656_);
  and (_03702_, _03701_, _02022_);
  and (_03703_, _03674_, _03656_);
  and (_03704_, _03703_, _02037_);
  nor (_03705_, _03704_, _03702_);
  and (_03706_, _03705_, _03700_);
  and (_03707_, _03706_, _03695_);
  and (_03708_, _03707_, _03684_);
  nor (_03709_, _03708_, _03589_);
  not (_03710_, _03505_);
  nor (_03711_, _03615_, _03508_);
  nor (_03712_, _03711_, _03581_);
  not (_03713_, _03712_);
  and (_03714_, _03504_, _03507_);
  and (_03715_, _03504_, _03609_);
  or (_03716_, _03715_, _03714_);
  and (_03717_, _03716_, _03583_);
  and (_03718_, _03590_, _03452_);
  and (_03719_, _03504_, _03590_);
  nor (_03720_, _03719_, _03718_);
  not (_03721_, _03711_);
  not (_03722_, \oc8051_golden_model_1.SP [3]);
  and (_03723_, _03609_, _03452_);
  and (_03724_, _03723_, _03722_);
  not (_03725_, _03234_);
  and (_03726_, _03725_, _03221_);
  nor (_03727_, _03726_, _03610_);
  or (_03728_, _03727_, _03581_);
  and (_03729_, _03507_, _03221_);
  nor (_03730_, _03723_, _03715_);
  nand (_03731_, _03727_, \oc8051_golden_model_1.PSW [3]);
  and (_03732_, _03731_, _03730_);
  or (_03733_, _03732_, _03729_);
  and (_03734_, _03733_, _03728_);
  or (_03735_, _03734_, _03724_);
  not (_03736_, _03714_);
  not (_03737_, _03729_);
  or (_03738_, _03737_, _03581_);
  and (_03739_, _03738_, _03736_);
  and (_03740_, _03739_, _03735_);
  or (_03741_, _03740_, _03721_);
  and (_03742_, _03741_, _03720_);
  or (_03743_, _03742_, _03717_);
  and (_03744_, _03743_, _03713_);
  nor (_03745_, _03237_, _03219_);
  not (_03746_, _03720_);
  and (_03747_, _03746_, _03583_);
  nor (_03748_, _03747_, _03745_);
  not (_03749_, _03748_);
  nor (_03750_, _03749_, _03744_);
  not (_03751_, _03237_);
  and (_03752_, _03751_, _03452_);
  and (_03753_, _03504_, _03751_);
  nor (_03754_, _03753_, _03752_);
  not (_03755_, _03754_);
  not (_03756_, _03581_);
  and (_03757_, _03745_, _03756_);
  nor (_03758_, _03757_, _03755_);
  not (_03759_, _03758_);
  nor (_03760_, _03759_, _03750_);
  and (_03761_, _03223_, _03221_);
  and (_03762_, _03755_, _03583_);
  nor (_03763_, _03762_, _03761_);
  not (_03764_, _03763_);
  nor (_03765_, _03764_, _03760_);
  not (_03766_, _03761_);
  nor (_03767_, _03766_, _03581_);
  or (_03768_, _03767_, _03765_);
  and (_03769_, _03768_, _03710_);
  nor (_03770_, _03583_, _03710_);
  or (_03771_, _03770_, _03769_);
  and (_03772_, _03771_, _03589_);
  or (_03773_, _03772_, _03587_);
  nor (_03774_, _03773_, _03709_);
  nor (_03775_, _03774_, _03588_);
  and (_03776_, _03221_, _03187_);
  not (_03777_, _03776_);
  and (_03778_, _03221_, _03181_);
  not (_03779_, _03778_);
  and (_03780_, _03504_, _03181_);
  nor (_03781_, _03780_, _03600_);
  and (_03782_, _03781_, _03779_);
  and (_03783_, _03221_, _03200_);
  not (_03784_, _03783_);
  and (_03785_, _03504_, _03200_);
  nor (_03786_, _03785_, _03624_);
  and (_03787_, _03786_, _03784_);
  and (_03788_, _03221_, _03191_);
  not (_03789_, _03788_);
  and (_03790_, _03504_, _03191_);
  nor (_03791_, _03790_, _03622_);
  and (_03792_, _03791_, _03789_);
  and (_03793_, _03792_, _03787_);
  and (_03794_, _03793_, _03782_);
  and (_03795_, _03794_, _03777_);
  not (_03796_, _03795_);
  nor (_03797_, _03796_, _03775_);
  and (_03798_, _03504_, _03187_);
  and (_03799_, _03796_, _03581_);
  nor (_03800_, _03799_, _03798_);
  not (_03801_, _03800_);
  nor (_03802_, _03801_, _03797_);
  and (_03803_, _03798_, \oc8051_golden_model_1.SP [3]);
  or (_03804_, _03803_, _03621_);
  nor (_03805_, _03804_, _03802_);
  and (_03806_, _03583_, _03621_);
  or (_03807_, _03806_, _03805_);
  and (_03808_, _03807_, _03518_);
  and (_03809_, _03517_, _03581_);
  or (_03810_, _03809_, _03808_);
  nand (_03811_, _03810_, _03516_);
  and (_03812_, _03515_, _03722_);
  nor (_03813_, _03812_, _03628_);
  nand (_03814_, _03813_, _03811_);
  and (_03815_, _03221_, _03197_);
  not (_03816_, _03628_);
  nor (_03817_, _03816_, _03583_);
  nor (_03818_, _03817_, _03815_);
  nand (_03819_, _03818_, _03814_);
  and (_03820_, _03815_, _03581_);
  nor (_03821_, _03820_, _03453_);
  and (_03822_, _03821_, _03819_);
  not (_03823_, _03453_);
  nor (_03824_, _03583_, _03823_);
  or (_03825_, _03824_, _03822_);
  nand (_03826_, _03825_, _03514_);
  nor (_03827_, _03514_, _03581_);
  not (_03828_, _03827_);
  and (_03829_, _03828_, _03826_);
  nor (_03830_, _03391_, _42316_);
  nor (_03831_, _03370_, _42152_);
  nor (_03832_, _03831_, _03830_);
  nor (_03833_, _03363_, _41906_);
  nor (_03834_, _03374_, _41686_);
  nor (_03835_, _03834_, _03833_);
  and (_03836_, _03835_, _03832_);
  nor (_03837_, _03378_, _42111_);
  nor (_03838_, _03380_, _42070_);
  nor (_03839_, _03838_, _03837_);
  nor (_03840_, _03384_, _42275_);
  nor (_03841_, _03393_, _42193_);
  nor (_03842_, _03841_, _03840_);
  and (_03843_, _03842_, _03839_);
  and (_03844_, _03843_, _03836_);
  nor (_03845_, _03386_, _41824_);
  nor (_03846_, _03404_, _41775_);
  nor (_03847_, _03846_, _03845_);
  nor (_03848_, _03396_, _41988_);
  nor (_03849_, _03409_, _41727_);
  nor (_03850_, _03849_, _03848_);
  and (_03851_, _03850_, _03847_);
  nor (_03852_, _03407_, _42234_);
  nor (_03853_, _03402_, _42029_);
  nor (_03854_, _03853_, _03852_);
  nor (_03855_, _03358_, _41947_);
  nor (_03856_, _03398_, _41865_);
  nor (_03857_, _03856_, _03855_);
  and (_03858_, _03857_, _03854_);
  and (_03859_, _03858_, _03851_);
  and (_03860_, _03859_, _03844_);
  nor (_03861_, _03860_, _03454_);
  and (_03862_, _03861_, _03715_);
  not (_03863_, _03862_);
  not (_03864_, _03861_);
  nor (_03865_, _03621_, _03453_);
  and (_03866_, _03865_, _03754_);
  and (_03867_, _03866_, _03720_);
  nor (_03868_, _03628_, _03714_);
  and (_03869_, _03586_, _03710_);
  and (_03870_, _03869_, _03868_);
  and (_03872_, _03870_, _03867_);
  nor (_03873_, _03872_, _03864_);
  nor (_03874_, _03396_, _41973_);
  nor (_03875_, _03386_, _41809_);
  nor (_03876_, _03875_, _03874_);
  nor (_03877_, _03393_, _42178_);
  nor (_03878_, _03380_, _42055_);
  nor (_03879_, _03878_, _03877_);
  and (_03880_, _03879_, _03876_);
  nor (_03881_, _03358_, _41932_);
  nor (_03882_, _03363_, _41891_);
  nor (_03883_, _03882_, _03881_);
  nor (_03884_, _03404_, _41758_);
  nor (_03885_, _03409_, _41712_);
  nor (_03886_, _03885_, _03884_);
  and (_03887_, _03886_, _03883_);
  and (_03888_, _03887_, _03880_);
  nor (_03889_, _03370_, _42137_);
  nor (_03890_, _03378_, _42096_);
  nor (_03891_, _03890_, _03889_);
  nor (_03892_, _03391_, _42301_);
  nor (_03893_, _03402_, _42014_);
  nor (_03894_, _03893_, _03892_);
  and (_03895_, _03894_, _03891_);
  nor (_03896_, _03384_, _42260_);
  nor (_03897_, _03407_, _42219_);
  nor (_03898_, _03897_, _03896_);
  nor (_03899_, _03398_, _41850_);
  nor (_03900_, _03374_, _41671_);
  nor (_03901_, _03900_, _03899_);
  and (_03902_, _03901_, _03898_);
  and (_03903_, _03902_, _03895_);
  and (_03904_, _03903_, _03888_);
  nor (_03905_, _03761_, _03745_);
  and (_03906_, _03905_, _03737_);
  and (_03907_, _03727_, _03711_);
  and (_03908_, _03907_, _03906_);
  nor (_03909_, _03815_, _03447_);
  and (_03910_, _03909_, _03777_);
  and (_03911_, _03910_, _03518_);
  and (_03912_, _03911_, _03908_);
  and (_03913_, _03912_, _03794_);
  nor (_03914_, _03913_, _03904_);
  not (_03915_, _03914_);
  and (_03916_, _03690_, _01997_);
  and (_03917_, _03654_, _01977_);
  nor (_03918_, _03917_, _03916_);
  and (_03919_, _03672_, _01992_);
  and (_03920_, _03680_, _01965_);
  nor (_03921_, _03920_, _03919_);
  and (_03922_, _03921_, _03918_);
  and (_03923_, _03692_, _02005_);
  and (_03924_, _03657_, _01979_);
  nor (_03925_, _03924_, _03923_);
  and (_03926_, _03696_, _01972_);
  and (_03927_, _03665_, _02000_);
  nor (_03928_, _03927_, _03926_);
  and (_03929_, _03928_, _03925_);
  and (_03930_, _03929_, _03922_);
  and (_03931_, _03675_, _01986_);
  and (_03932_, _03678_, _02014_);
  nor (_03933_, _03932_, _03931_);
  and (_03934_, _03687_, _01989_);
  and (_03935_, _03703_, _01970_);
  nor (_03936_, _03935_, _03934_);
  and (_03937_, _03936_, _03933_);
  and (_03938_, _03685_, _02002_);
  and (_03939_, _03701_, _01967_);
  nor (_03940_, _03939_, _03938_);
  and (_03941_, _03662_, _02012_);
  and (_03942_, _03698_, _01974_);
  nor (_03943_, _03942_, _03941_);
  and (_03944_, _03943_, _03940_);
  and (_03945_, _03944_, _03937_);
  and (_03946_, _03945_, _03930_);
  nor (_03947_, _03946_, _03589_);
  not (_03948_, _03490_);
  not (_03949_, _03202_);
  nor (_03950_, _03590_, _03191_);
  and (_03951_, _03950_, _03949_);
  nor (_03952_, _03951_, _03948_);
  not (_03953_, _03952_);
  and (_03954_, _03489_, _03027_);
  not (_03955_, _03954_);
  nor (_03956_, _03590_, _03187_);
  and (_03957_, _03956_, _03212_);
  nor (_03958_, _03957_, _03955_);
  not (_03959_, _03958_);
  and (_03960_, _03489_, _03195_);
  not (_03961_, _03960_);
  and (_03962_, _03489_, _03609_);
  and (_03963_, _03490_, _03181_);
  nor (_03964_, _03963_, _03962_);
  and (_03965_, _03964_, _03961_);
  and (_03966_, _03965_, _03959_);
  and (_03967_, _03966_, _03953_);
  and (_03968_, _03592_, _03187_);
  and (_03969_, _03595_, _03168_);
  nor (_03970_, _03969_, _03968_);
  and (_03971_, _03954_, _03200_);
  and (_03972_, _03954_, _03197_);
  nor (_03973_, _03972_, _03971_);
  nor (_03974_, _03223_, _03181_);
  nor (_03975_, _03974_, _03955_);
  not (_03976_, _03975_);
  and (_03977_, _03976_, _03973_);
  and (_03978_, _03977_, _03970_);
  and (_03979_, _03954_, _03725_);
  and (_03980_, _03592_, _03725_);
  or (_03981_, _03980_, _03979_);
  and (_03982_, _03954_, _03191_);
  nor (_03983_, _03982_, _03981_);
  and (_03984_, _03490_, _03200_);
  and (_03985_, _03489_, _03507_);
  nor (_03986_, _03985_, _03984_);
  and (_03987_, _03986_, _03983_);
  and (_03988_, _03595_, _03223_);
  not (_03989_, _03988_);
  and (_03990_, _03954_, _03202_);
  nor (_03991_, _03491_, _03990_);
  and (_03992_, _03991_, _03989_);
  and (_03993_, _03992_, _03987_);
  and (_03994_, _03993_, _03978_);
  not (_03995_, \oc8051_golden_model_1.SP [2]);
  not (_03996_, _03723_);
  nor (_03997_, _03798_, _03515_);
  and (_03998_, _03997_, _03996_);
  nor (_03999_, _03998_, _03995_);
  or (_04000_, _03223_, _03168_);
  and (_04001_, _04000_, _03592_);
  not (_04002_, _04001_);
  and (_04003_, _03595_, _03187_);
  and (_04004_, _03595_, _03725_);
  nor (_04005_, _04004_, _04003_);
  and (_04006_, _04005_, _04002_);
  not (_04007_, _04006_);
  nor (_04008_, _04007_, _03999_);
  and (_04009_, _04008_, _03994_);
  and (_04010_, _04009_, _03967_);
  not (_04011_, _04010_);
  nor (_04012_, _04011_, _03947_);
  and (_04013_, _04012_, _03915_);
  not (_04014_, _04013_);
  nor (_04015_, _04014_, _03873_);
  and (_04016_, _04015_, _03863_);
  not (_04017_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_04018_, _03384_, _42250_);
  or (_04019_, _03407_, _42209_);
  and (_04020_, _04019_, _04018_);
  or (_04021_, _03370_, _42127_);
  or (_04022_, _03378_, _42086_);
  and (_04023_, _04022_, _04021_);
  and (_04024_, _04023_, _04020_);
  or (_04025_, _03374_, _41661_);
  or (_04026_, _03409_, _41702_);
  and (_04027_, _04026_, _04025_);
  or (_04028_, _03363_, _41881_);
  or (_04029_, _03398_, _41840_);
  and (_04030_, _04029_, _04028_);
  and (_04031_, _04030_, _04027_);
  and (_04032_, _04031_, _04024_);
  or (_04033_, _03380_, _42045_);
  or (_04034_, _03402_, _42004_);
  and (_04035_, _04034_, _04033_);
  or (_04036_, _03391_, _42291_);
  or (_04037_, _03393_, _42168_);
  and (_04038_, _04037_, _04036_);
  and (_04039_, _04038_, _04035_);
  or (_04040_, _03396_, _41963_);
  or (_04041_, _03358_, _41922_);
  and (_04042_, _04041_, _04040_);
  or (_04043_, _03386_, _41791_);
  or (_04044_, _03404_, _41743_);
  and (_04045_, _04044_, _04043_);
  and (_04046_, _04045_, _04042_);
  and (_04047_, _04046_, _04039_);
  and (_04048_, _04047_, _04032_);
  nor (_04049_, _04048_, _03514_);
  not (_04050_, _04049_);
  and (_04051_, _03756_, _03446_);
  and (_04052_, _04051_, _03453_);
  and (_04053_, _03505_, _04051_);
  nor (_04054_, _04048_, _03766_);
  not (_04055_, _03715_);
  not (_04056_, _03726_);
  nor (_04057_, _04048_, _04056_);
  and (_04058_, _03493_, _03451_);
  nor (_04059_, _03605_, _04058_);
  nor (_04060_, _04059_, _03234_);
  not (_04061_, _04060_);
  not (_04062_, _03239_);
  and (_04063_, _03605_, _04062_);
  and (_04064_, _03591_, _03725_);
  nor (_04065_, _04064_, _04063_);
  and (_04066_, _03493_, _03503_);
  and (_04067_, _04066_, _03725_);
  not (_04068_, _04067_);
  nor (_04069_, _04004_, _03726_);
  and (_04070_, _04069_, _04068_);
  and (_04071_, _04070_, _04065_);
  and (_04073_, _04071_, _04061_);
  or (_04074_, _04073_, _04057_);
  and (_04075_, _03489_, _02994_);
  nor (_04076_, _04066_, _04075_);
  and (_04077_, _04076_, _04059_);
  nor (_04078_, _04077_, _03229_);
  nor (_04079_, _04078_, _03610_);
  nand (_04080_, _04079_, _04074_);
  not (_04081_, _03610_);
  or (_04082_, _04048_, _04081_);
  nand (_04083_, _04082_, _04080_);
  nand (_04084_, _04083_, _04055_);
  nand (_04085_, _03715_, _04051_);
  nand (_04086_, _04085_, _04084_);
  and (_04087_, _03723_, _03498_);
  nor (_04088_, _04087_, _03729_);
  not (_04089_, _04088_);
  nor (_04090_, _04077_, _03232_);
  nor (_04091_, _04090_, _04089_);
  and (_04092_, _04091_, _04086_);
  nor (_04093_, _04048_, _03737_);
  or (_04094_, _04093_, _04092_);
  and (_04095_, _04094_, _03736_);
  and (_04096_, _03714_, _04051_);
  or (_04097_, _04096_, _04095_);
  and (_04098_, _04048_, _03508_);
  nor (_04099_, _03606_, _03615_);
  and (_04100_, _02994_, _02962_);
  and (_04101_, _04100_, _03590_);
  not (_04102_, _04101_);
  and (_04103_, _04102_, _04099_);
  not (_04104_, _04103_);
  nor (_04105_, _04104_, _04098_);
  and (_04106_, _04105_, _04097_);
  not (_04107_, _03615_);
  nor (_04108_, _04048_, _04107_);
  or (_04109_, _04108_, _04106_);
  nand (_04110_, _04109_, _03720_);
  and (_04111_, _03746_, _04051_);
  nor (_04112_, _04111_, _03745_);
  nand (_04113_, _04112_, _04110_);
  and (_04114_, _04048_, _03745_);
  and (_04115_, _03605_, _03751_);
  nor (_04116_, _04115_, _03755_);
  not (_04117_, _04116_);
  nor (_04118_, _04117_, _04114_);
  and (_04119_, _04118_, _04113_);
  and (_04120_, _03755_, _04051_);
  nor (_04121_, _04120_, _04119_);
  nor (_04122_, _04066_, _03591_);
  nor (_04123_, _03595_, _03221_);
  and (_04124_, _04123_, _04059_);
  and (_04125_, _04124_, _04122_);
  nor (_04126_, _04125_, _03247_);
  nor (_04127_, _04126_, _04121_);
  or (_04128_, _04127_, _04054_);
  and (_04129_, _04128_, _03710_);
  nor (_04130_, _04129_, _04053_);
  nor (_04131_, _04077_, _03212_);
  nor (_04132_, _04131_, _04130_);
  and (_04133_, _03665_, _01864_);
  and (_04134_, _03678_, _01900_);
  nor (_04135_, _04134_, _04133_);
  and (_04136_, _03685_, _01890_);
  and (_04137_, _03654_, _01888_);
  nor (_04138_, _04137_, _04136_);
  and (_04139_, _04138_, _04135_);
  and (_04140_, _03698_, _01862_);
  and (_04141_, _03675_, _01885_);
  nor (_04142_, _04141_, _04140_);
  and (_04143_, _03680_, _01869_);
  and (_04144_, _03703_, _01871_);
  nor (_04145_, _04144_, _04143_);
  and (_04146_, _04145_, _04142_);
  and (_04147_, _04146_, _04139_);
  and (_04148_, _03662_, _01875_);
  and (_04149_, _03692_, _01893_);
  nor (_04150_, _04149_, _04148_);
  and (_04151_, _03672_, _01877_);
  and (_04152_, _03701_, _01853_);
  nor (_04153_, _04152_, _04151_);
  and (_04154_, _04153_, _04150_);
  and (_04155_, _03690_, _01879_);
  and (_04156_, _03696_, _01859_);
  nor (_04157_, _04156_, _04155_);
  and (_04158_, _03687_, _01902_);
  and (_04159_, _03657_, _01856_);
  nor (_04160_, _04159_, _04158_);
  and (_04161_, _04160_, _04157_);
  and (_04162_, _04161_, _04154_);
  and (_04163_, _04162_, _04147_);
  and (_04164_, _04163_, _03222_);
  nor (_04165_, _04164_, _03585_);
  and (_04166_, _04165_, _04132_);
  and (_04167_, _03585_, _04051_);
  or (_04168_, _04167_, _04166_);
  and (_04169_, _03605_, _03176_);
  nor (_04170_, _04169_, _03584_);
  and (_04171_, _04170_, _04168_);
  and (_04172_, _03584_, _04051_);
  or (_04174_, _04172_, _04171_);
  not (_04175_, _03181_);
  nor (_04176_, _04058_, _03591_);
  nor (_04177_, _04176_, _04175_);
  not (_04178_, _04177_);
  and (_04179_, _03963_, _02994_);
  not (_04180_, _04179_);
  and (_04181_, _04066_, _03181_);
  and (_04182_, _03605_, _03181_);
  nor (_04183_, _04182_, _04181_);
  and (_04184_, _04183_, _04180_);
  and (_04185_, _04184_, _04178_);
  and (_04186_, _04185_, _04174_);
  and (_04187_, _03792_, _03782_);
  not (_04188_, _04048_);
  nor (_04189_, _04188_, _04187_);
  not (_04190_, _03200_);
  nor (_04191_, _04077_, _04190_);
  not (_04192_, _04191_);
  not (_04193_, _03191_);
  nor (_04194_, _03605_, _04075_);
  nor (_04195_, _04194_, _04193_);
  not (_04196_, _04195_);
  and (_04197_, _04066_, _03191_);
  and (_04198_, _03494_, _03191_);
  and (_04199_, _04198_, _02994_);
  nor (_04200_, _04199_, _04197_);
  and (_04201_, _04200_, _04196_);
  and (_04202_, _04201_, _04192_);
  not (_04203_, _04202_);
  nor (_04204_, _04203_, _04189_);
  and (_04205_, _04204_, _04186_);
  nor (_04206_, _04188_, _03787_);
  not (_04207_, _03187_);
  nor (_04208_, _03605_, _03221_);
  and (_04209_, _04208_, _04122_);
  nor (_04210_, _04209_, _04207_);
  and (_04211_, _04058_, _03187_);
  nor (_04212_, _04211_, _04003_);
  not (_04213_, _04212_);
  nor (_04214_, _04213_, _04210_);
  not (_04215_, _04214_);
  nor (_04216_, _04215_, _04206_);
  and (_04217_, _04216_, _04205_);
  nor (_04218_, _04048_, _03777_);
  or (_04219_, _04218_, _04217_);
  and (_04220_, _03798_, _03498_);
  nor (_04221_, _04220_, _03621_);
  and (_04222_, _04221_, _04219_);
  and (_04223_, _03621_, _04051_);
  or (_04224_, _04223_, _04222_);
  and (_04225_, _03591_, _03202_);
  and (_04226_, _04066_, _03202_);
  nor (_04227_, _04226_, _04225_);
  not (_04228_, _04227_);
  nor (_04229_, _04124_, _03949_);
  nor (_04230_, _04229_, _04228_);
  and (_04231_, _04230_, _04224_);
  nor (_04232_, _04048_, _03518_);
  or (_04233_, _04232_, _04231_);
  and (_04234_, _03515_, _03498_);
  nor (_04235_, _04234_, _03628_);
  and (_04236_, _04235_, _04233_);
  and (_04237_, _03628_, _04051_);
  or (_04238_, _04237_, _04236_);
  and (_04239_, _02994_, _03197_);
  and (_04240_, _04239_, _02962_);
  not (_04241_, _04240_);
  and (_04242_, _03605_, _03197_);
  nor (_04243_, _04242_, _03815_);
  and (_04244_, _04243_, _04241_);
  and (_04245_, _04244_, _04238_);
  not (_04246_, _03815_);
  nor (_04247_, _04048_, _04246_);
  or (_04248_, _04247_, _04245_);
  and (_04249_, _04248_, _03823_);
  or (_04250_, _04249_, _04052_);
  and (_04251_, _03960_, _02994_);
  not (_04252_, _04251_);
  and (_04253_, _03493_, _03195_);
  and (_04254_, _04253_, _02994_);
  not (_04255_, _04254_);
  and (_04256_, _03605_, _03195_);
  nor (_04257_, _04256_, _03447_);
  and (_04258_, _04257_, _04255_);
  and (_04259_, _04258_, _04252_);
  nand (_04260_, _04259_, _04250_);
  nand (_04261_, _04260_, _04050_);
  or (_04262_, _04261_, _04017_);
  nor (_04263_, _03715_, _03505_);
  and (_04264_, _03868_, _03586_);
  and (_04265_, _04264_, _04263_);
  and (_04266_, _04265_, _03867_);
  not (_04267_, _04266_);
  and (_04268_, _04267_, _03487_);
  not (_04269_, _04268_);
  nor (_04270_, _03414_, _03913_);
  not (_04271_, _04270_);
  and (_04272_, _03692_, _01949_);
  and (_04273_, _03654_, _01917_);
  nor (_04275_, _04273_, _04272_);
  and (_04276_, _03672_, _01933_);
  and (_04277_, _03680_, _01924_);
  nor (_04278_, _04277_, _04276_);
  and (_04279_, _04278_, _04275_);
  and (_04280_, _03685_, _01946_);
  and (_04281_, _03657_, _01944_);
  nor (_04282_, _04281_, _04280_);
  and (_04283_, _03687_, _01958_);
  and (_04284_, _03665_, _01919_);
  nor (_04285_, _04284_, _04283_);
  and (_04286_, _04285_, _04282_);
  and (_04287_, _04286_, _04279_);
  and (_04288_, _03675_, _01930_);
  and (_04289_, _03678_, _01956_);
  nor (_04290_, _04289_, _04288_);
  and (_04291_, _03696_, _01914_);
  and (_04292_, _03703_, _01926_);
  nor (_04293_, _04292_, _04291_);
  and (_04294_, _04293_, _04290_);
  and (_04295_, _03662_, _01941_);
  and (_04296_, _03701_, _01909_);
  nor (_04297_, _04296_, _04295_);
  and (_04298_, _03690_, _01937_);
  and (_04299_, _03698_, _01912_);
  nor (_04300_, _04299_, _04298_);
  and (_04301_, _04300_, _04297_);
  and (_04302_, _04301_, _04294_);
  and (_04303_, _04302_, _04287_);
  nor (_04304_, _04303_, _03589_);
  and (_04305_, _03493_, _03027_);
  and (_04306_, _04305_, _03200_);
  and (_04307_, _04305_, _03609_);
  nor (_04308_, _04307_, _04306_);
  and (_04309_, _04305_, _03168_);
  and (_04310_, _04305_, _03202_);
  nor (_04311_, _04310_, _04309_);
  and (_04312_, _04311_, _04308_);
  and (_04313_, _03954_, _03609_);
  nor (_04314_, _03982_, _04313_);
  and (_04315_, _04305_, _03191_);
  nor (_04316_, _04315_, _03979_);
  and (_04317_, _04316_, _04314_);
  and (_04318_, _04317_, _04312_);
  and (_04319_, _04318_, _03959_);
  and (_04320_, _04305_, _03195_);
  not (_04321_, _04320_);
  and (_04322_, _04305_, _03197_);
  and (_04323_, _03985_, _03027_);
  nor (_04324_, _04323_, _04322_);
  and (_04325_, _04324_, _04321_);
  and (_04326_, _04305_, _03590_);
  nor (_04327_, _03990_, _04326_);
  and (_04328_, _04327_, _03973_);
  and (_04329_, _03954_, _03195_);
  nor (_04330_, _04329_, _03975_);
  and (_04331_, _04330_, _04328_);
  and (_04332_, _04331_, _04325_);
  not (_04333_, _04305_);
  and (_04334_, _03234_, _03247_);
  nor (_04335_, _03181_, _03187_);
  and (_04336_, _04335_, _03232_);
  and (_04337_, _04336_, _04334_);
  nor (_04338_, _04337_, _04333_);
  nor (_04339_, _03998_, _03496_);
  nor (_04340_, _04339_, _04338_);
  and (_04341_, _04340_, _04332_);
  and (_04342_, _04341_, _04319_);
  not (_04343_, _04342_);
  nor (_04344_, _04343_, _04304_);
  and (_04345_, _04344_, _04271_);
  and (_04346_, _04345_, _04269_);
  not (_04347_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_04348_, _04260_, _04050_);
  or (_04349_, _04348_, _04347_);
  and (_04350_, _04349_, _04346_);
  nand (_04351_, _04350_, _04262_);
  not (_04352_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_04353_, _04348_, _04352_);
  not (_04354_, _04346_);
  not (_04355_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_04356_, _04261_, _04355_);
  and (_04357_, _04356_, _04354_);
  nand (_04358_, _04357_, _04353_);
  nand (_04359_, _04358_, _04351_);
  nand (_04360_, _04359_, _04016_);
  not (_04361_, _04016_);
  not (_04362_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_04363_, _04348_, _04362_);
  not (_04364_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_04365_, _04261_, _04364_);
  and (_04366_, _04365_, _04354_);
  nand (_04367_, _04366_, _04363_);
  not (_04368_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_04369_, _04261_, _04368_);
  not (_04370_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_04371_, _04348_, _04370_);
  and (_04372_, _04371_, _04346_);
  nand (_04373_, _04372_, _04369_);
  nand (_04374_, _04373_, _04367_);
  nand (_04376_, _04374_, _04361_);
  nand (_04377_, _04376_, _04360_);
  nand (_04378_, _04377_, _03829_);
  not (_04379_, _03829_);
  not (_04380_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_04381_, _04348_, _04380_);
  nand (_04382_, _04348_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_04383_, _04382_, _04354_);
  nand (_04384_, _04383_, _04381_);
  not (_04385_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_04386_, _04261_, _04385_);
  nand (_04387_, _04261_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_04388_, _04387_, _04346_);
  nand (_04389_, _04388_, _04386_);
  nand (_04390_, _04389_, _04384_);
  nand (_04391_, _04390_, _04016_);
  not (_04392_, \oc8051_golden_model_1.IRAM[15] [1]);
  or (_04393_, _04348_, _04392_);
  nand (_04394_, _04348_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_04395_, _04394_, _04354_);
  nand (_04396_, _04395_, _04393_);
  not (_04397_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_04398_, _04261_, _04397_);
  nand (_04399_, _04261_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_04400_, _04399_, _04346_);
  nand (_04401_, _04400_, _04398_);
  nand (_04402_, _04401_, _04396_);
  nand (_04403_, _04402_, _04361_);
  nand (_04404_, _04403_, _04391_);
  nand (_04405_, _04404_, _04379_);
  nand (_04406_, _04405_, _04378_);
  and (_04407_, _04406_, _03513_);
  or (_04408_, _04407_, _03512_);
  and (_04409_, _03612_, _03725_);
  and (_04410_, _04409_, _03446_);
  and (_04411_, _03414_, _04410_);
  or (_04412_, _04411_, _04408_);
  and (_04413_, _03500_, _03980_);
  not (_04414_, _04413_);
  and (_04415_, _03490_, _03609_);
  and (_04416_, _03494_, _03609_);
  nor (_04417_, _04416_, _04415_);
  and (_04418_, _04417_, _04414_);
  not (_04419_, _04418_);
  nor (_04420_, _04419_, _04412_);
  and (_04421_, _03610_, _03446_);
  nor (_04422_, _03511_, _03229_);
  and (_04423_, _04406_, _04422_);
  nor (_04424_, _04423_, _04421_);
  and (_04425_, _04424_, _04420_);
  and (_04426_, _04421_, _03415_);
  nor (_04427_, _04426_, _04425_);
  and (_04428_, _03715_, _03446_);
  and (_04429_, _03486_, _04428_);
  nor (_04430_, _04429_, _04427_);
  and (_04431_, _03723_, _03446_);
  nor (_04432_, _03501_, _03230_);
  nor (_04433_, _04432_, _04431_);
  and (_04434_, _04433_, _04430_);
  and (_04435_, _04431_, _03415_);
  nor (_04436_, _04435_, _04434_);
  and (_04437_, _03490_, _03507_);
  and (_04438_, _03494_, _03507_);
  nor (_04439_, _04438_, _04437_);
  not (_04440_, _04439_);
  nor (_04441_, _04440_, _04436_);
  and (_04442_, _03729_, _03446_);
  nor (_04443_, _03511_, _03232_);
  and (_04444_, _04406_, _04443_);
  nor (_04445_, _04444_, _04442_);
  and (_04446_, _04445_, _04441_);
  and (_04447_, _04442_, _03415_);
  nor (_04448_, _04447_, _04446_);
  and (_04449_, _03714_, _03446_);
  and (_04450_, _03486_, _04449_);
  nor (_04451_, _04450_, _04448_);
  and (_04452_, _04451_, _03510_);
  nor (_04453_, _04452_, _03509_);
  and (_04454_, _03719_, _03446_);
  and (_04455_, _04454_, _03486_);
  or (_04456_, _04455_, _04453_);
  nor (_04457_, _03501_, _03227_);
  and (_04458_, _03745_, _03213_);
  nor (_04459_, _04458_, _04457_);
  not (_04460_, _04459_);
  nor (_04461_, _04460_, _04456_);
  and (_04462_, _03505_, _03446_);
  nor (_04463_, _03511_, _03237_);
  and (_04464_, _04406_, _04463_);
  nor (_04465_, _04464_, _04462_);
  and (_04466_, _04465_, _04461_);
  nor (_04467_, _04466_, _03506_);
  nor (_04468_, _04467_, _03224_);
  and (_04469_, _03501_, _03224_);
  nor (_04470_, _04469_, _04468_);
  and (_04471_, _03446_, _03168_);
  and (_04472_, _04471_, _03494_);
  not (_04473_, _04309_);
  or (_04474_, _03592_, _03954_);
  and (_04475_, _04474_, _03168_);
  nor (_04477_, _04475_, _03969_);
  and (_04478_, _04477_, _04473_);
  nor (_04479_, _04478_, _03454_);
  nor (_04480_, _04479_, _04472_);
  nor (_04481_, _03511_, _03212_);
  and (_04482_, _04481_, _03446_);
  and (_04483_, _04471_, _03221_);
  nor (_04484_, _04483_, _04482_);
  and (_04485_, _04484_, _04480_);
  nor (_04486_, _04485_, _03415_);
  and (_04487_, _03592_, _03176_);
  and (_04488_, _03493_, _03218_);
  and (_04489_, _04488_, _03176_);
  or (_04490_, _04489_, _04487_);
  not (_04491_, _04490_);
  and (_04492_, _04058_, _03176_);
  and (_04493_, _03595_, _03176_);
  nor (_04494_, _04493_, _04492_);
  and (_04495_, _04494_, _04491_);
  not (_04496_, _04495_);
  nor (_04497_, _04496_, _04486_);
  not (_04498_, _04497_);
  nor (_04499_, _04498_, _04470_);
  and (_04500_, _03601_, _03446_);
  not (_04501_, _03176_);
  nor (_04502_, _03511_, _04501_);
  and (_04503_, _04406_, _04502_);
  nor (_04504_, _04503_, _04500_);
  and (_04505_, _04504_, _04499_);
  and (_04506_, _04500_, _03415_);
  nor (_04507_, _04506_, _04505_);
  nor (_04508_, _04507_, _03178_);
  and (_04509_, _03501_, _03178_);
  nor (_04510_, _04509_, _04508_);
  and (_04511_, _03780_, _03446_);
  and (_04512_, _03600_, _03446_);
  nor (_04513_, _04512_, _04511_);
  and (_04514_, _03790_, _03446_);
  and (_04515_, _03622_, _03446_);
  nor (_04516_, _04515_, _04514_);
  and (_04517_, _04516_, _04513_);
  nor (_04518_, _04517_, _03415_);
  nor (_04519_, _04518_, _03192_);
  not (_04520_, _04519_);
  nor (_04521_, _04520_, _04510_);
  and (_04522_, _03501_, _03192_);
  nor (_04523_, _04522_, _04521_);
  nor (_04524_, _03786_, _03454_);
  and (_04525_, _04524_, _03414_);
  or (_04526_, _04525_, _03188_);
  nor (_04527_, _04526_, _04523_);
  nor (_04528_, _04527_, _03502_);
  nor (_04529_, _04528_, _03495_);
  and (_04530_, _04529_, _03492_);
  and (_04531_, _03815_, _03446_);
  not (_04532_, _03197_);
  nor (_04533_, _03511_, _04532_);
  and (_04534_, _04406_, _04533_);
  nor (_04535_, _04534_, _04531_);
  and (_04536_, _04535_, _04530_);
  and (_04537_, _04531_, _03415_);
  nor (_04538_, _04537_, _04536_);
  and (_04539_, _03446_, _03453_);
  nor (_04540_, _03629_, _03198_);
  nor (_04541_, _03501_, _04540_);
  nor (_04542_, _04541_, _04539_);
  not (_04543_, _04542_);
  nor (_04544_, _04543_, _04538_);
  nor (_04545_, _04544_, _03488_);
  and (_04546_, _03490_, _03195_);
  and (_04547_, _03494_, _03195_);
  nor (_04548_, _04547_, _04546_);
  not (_04549_, _04548_);
  nor (_04550_, _04549_, _04545_);
  not (_04551_, _03195_);
  nor (_04552_, _03511_, _04551_);
  and (_04553_, _04406_, _04552_);
  nor (_04554_, _04553_, _03448_);
  and (_04555_, _04554_, _04550_);
  nor (_04556_, _04555_, _03449_);
  not (_04557_, _04556_);
  not (_04558_, _04539_);
  and (_04559_, _03188_, _03498_);
  nor (_04560_, _04485_, _04188_);
  and (_04561_, _03719_, _04051_);
  not (_04562_, _04454_);
  not (_04563_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_04564_, _04261_, _04563_);
  not (_04565_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_04566_, _04348_, _04565_);
  and (_04567_, _04566_, _04346_);
  nand (_04568_, _04567_, _04564_);
  not (_04569_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_04570_, _04348_, _04569_);
  not (_04571_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_04572_, _04261_, _04571_);
  and (_04573_, _04572_, _04354_);
  nand (_04574_, _04573_, _04570_);
  nand (_04575_, _04574_, _04568_);
  nand (_04576_, _04575_, _04016_);
  not (_04578_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_04579_, _04348_, _04578_);
  not (_04580_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_04581_, _04261_, _04580_);
  and (_04582_, _04581_, _04354_);
  nand (_04583_, _04582_, _04579_);
  not (_04584_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_04585_, _04261_, _04584_);
  not (_04586_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_04587_, _04348_, _04586_);
  and (_04588_, _04587_, _04346_);
  nand (_04589_, _04588_, _04585_);
  nand (_04590_, _04589_, _04583_);
  nand (_04591_, _04590_, _04361_);
  nand (_04592_, _04591_, _04576_);
  nand (_04593_, _04592_, _03829_);
  not (_04594_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_04595_, _04348_, _04594_);
  nand (_04596_, _04348_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_04597_, _04596_, _04354_);
  nand (_04598_, _04597_, _04595_);
  not (_04599_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_04600_, _04261_, _04599_);
  nand (_04601_, _04261_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_04602_, _04601_, _04346_);
  nand (_04603_, _04602_, _04600_);
  nand (_04604_, _04603_, _04598_);
  nand (_04605_, _04604_, _04016_);
  not (_04606_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_04607_, _04348_, _04606_);
  nand (_04608_, _04348_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_04609_, _04608_, _04354_);
  nand (_04610_, _04609_, _04607_);
  not (_04611_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_04612_, _04261_, _04611_);
  nand (_04613_, _04261_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_04614_, _04613_, _04346_);
  nand (_04615_, _04614_, _04612_);
  nand (_04616_, _04615_, _04610_);
  nand (_04617_, _04616_, _04361_);
  nand (_04618_, _04617_, _04605_);
  nand (_04619_, _04618_, _04379_);
  and (_04620_, _04619_, _04593_);
  and (_04621_, _04620_, _03513_);
  nor (_04622_, _03603_, _03030_);
  and (_04623_, _04622_, _04059_);
  nor (_04624_, _04623_, _03239_);
  not (_04625_, _04624_);
  nor (_04626_, _04625_, _04621_);
  and (_04627_, _04048_, _04410_);
  or (_04628_, _04627_, _04626_);
  and (_04629_, _03980_, \oc8051_golden_model_1.SP [0]);
  and (_04630_, _04100_, _03609_);
  nor (_04631_, _04630_, _04629_);
  not (_04632_, _04631_);
  nor (_04633_, _04632_, _04628_);
  nand (_04634_, _04619_, _04593_);
  and (_04635_, _04422_, _04634_);
  nor (_04636_, _04635_, _04421_);
  and (_04637_, _04636_, _04633_);
  and (_04638_, _04421_, _04188_);
  nor (_04639_, _04638_, _04637_);
  nor (_04640_, _04639_, _04428_);
  not (_04641_, _04640_);
  and (_04642_, _04641_, _04085_);
  nor (_04643_, _03230_, _03498_);
  nor (_04644_, _04643_, _04642_);
  and (_04645_, _04431_, _04048_);
  and (_04646_, _04100_, _03507_);
  nor (_04647_, _04646_, _04645_);
  and (_04648_, _04647_, _04644_);
  and (_04649_, _04443_, _04634_);
  not (_04650_, _04649_);
  and (_04651_, _04650_, _04648_);
  and (_04652_, _04442_, _04048_);
  nor (_04653_, _04652_, _04449_);
  and (_04654_, _04653_, _04651_);
  nor (_04655_, _04654_, _04096_);
  nor (_04656_, _04655_, _03508_);
  and (_04657_, _03508_, _03498_);
  or (_04658_, _04657_, _04656_);
  and (_04659_, _04658_, _04562_);
  nor (_04660_, _04659_, _04561_);
  nor (_04661_, _03227_, _03498_);
  and (_04662_, _04100_, _03751_);
  nor (_04663_, _04662_, _04661_);
  not (_04664_, _04663_);
  nor (_04665_, _04664_, _04660_);
  and (_04666_, _04463_, _04634_);
  nor (_04667_, _04666_, _04462_);
  and (_04668_, _04667_, _04665_);
  nor (_04669_, _04668_, _04053_);
  nor (_04670_, _04669_, _03224_);
  and (_04671_, _03224_, _03498_);
  nor (_04672_, _04671_, _04670_);
  and (_04673_, _04100_, _03176_);
  or (_04674_, _04673_, _04672_);
  nor (_04675_, _04674_, _04560_);
  and (_04676_, _04502_, _04634_);
  not (_04677_, _04676_);
  and (_04679_, _04677_, _04675_);
  and (_04680_, _04500_, _04048_);
  nor (_04681_, _04680_, _03178_);
  and (_04682_, _04681_, _04679_);
  and (_04683_, _03178_, _03498_);
  nor (_04684_, _04683_, _04682_);
  nor (_04685_, _04517_, _04188_);
  nor (_04686_, _04685_, _03192_);
  not (_04687_, _04686_);
  nor (_04688_, _04687_, _04684_);
  and (_04689_, _03192_, _03498_);
  nor (_04690_, _04689_, _04688_);
  and (_04691_, _04524_, _04048_);
  or (_04692_, _04691_, _03188_);
  nor (_04693_, _04692_, _04690_);
  nor (_04694_, _04693_, _04559_);
  nor (_04695_, _04694_, _04240_);
  and (_04696_, _04533_, _04634_);
  nor (_04697_, _04696_, _04531_);
  and (_04698_, _04697_, _04695_);
  and (_04699_, _04531_, _04188_);
  nor (_04700_, _04699_, _04698_);
  nor (_04701_, _04540_, _03498_);
  nor (_04702_, _04701_, _04700_);
  and (_04703_, _04702_, _04558_);
  nor (_04704_, _04703_, _04052_);
  and (_04705_, _04100_, _03195_);
  nor (_04706_, _04705_, _04704_);
  and (_04707_, _04552_, _04634_);
  nor (_04708_, _04707_, _03448_);
  and (_04709_, _04708_, _04706_);
  and (_04710_, _03448_, _04188_);
  nor (_04711_, _04710_, _04709_);
  nor (_04712_, _04483_, _04472_);
  not (_04713_, _03448_);
  and (_04714_, _03593_, _03176_);
  not (_04715_, _04714_);
  and (_04716_, _03493_, _03176_);
  and (_04717_, _04716_, _03027_);
  nor (_04718_, _04717_, _04546_);
  and (_04719_, _04718_, _04715_);
  and (_04720_, _04719_, _04325_);
  or (_04721_, _03593_, _03595_);
  and (_04722_, _04721_, _03751_);
  not (_04723_, _03221_);
  and (_04724_, _04622_, _04723_);
  nor (_04725_, _04724_, _03239_);
  not (_04726_, _03494_);
  and (_04727_, _03511_, _04726_);
  nor (_04728_, _04727_, _03239_);
  or (_04729_, _04728_, _04725_);
  nor (_04730_, _04729_, _04722_);
  and (_04731_, _04730_, _04720_);
  and (_04732_, _04716_, _03218_);
  nor (_04733_, _04732_, _04493_);
  nor (_04734_, _04502_, _04492_);
  and (_04735_, _04540_, _03193_);
  and (_04736_, _04735_, _04734_);
  and (_04737_, _04736_, _04733_);
  nor (_04738_, _04463_, _04443_);
  nor (_04739_, _04552_, _04422_);
  and (_04740_, _04739_, _04738_);
  nor (_04741_, _03491_, _03972_);
  nor (_04742_, _04307_, _03962_);
  and (_04743_, _04742_, _04741_);
  and (_04744_, _04743_, _04740_);
  not (_04745_, _03495_);
  and (_04746_, _03612_, _03751_);
  nor (_04747_, _04416_, _04746_);
  and (_04748_, _04747_, _04745_);
  and (_04749_, _04305_, _03751_);
  or (_04750_, _04488_, _04305_);
  and (_04751_, _04750_, _03507_);
  nor (_04752_, _04751_, _04749_);
  and (_04753_, _03494_, _03751_);
  and (_04754_, _03612_, _03176_);
  nor (_04755_, _04754_, _04753_);
  and (_04756_, _04755_, _04752_);
  and (_04757_, _04756_, _04748_);
  and (_04758_, _04757_, _04744_);
  and (_04759_, _04058_, _03507_);
  nor (_04760_, _04329_, _04759_);
  nor (_04761_, _04547_, _04437_);
  and (_04762_, _04761_, _04760_);
  not (_04763_, _03980_);
  nor (_04764_, _04533_, _03508_);
  and (_04765_, _04764_, _04763_);
  not (_04766_, _03227_);
  nor (_04767_, _04766_, _03224_);
  not (_04768_, _03230_);
  nor (_04769_, _04768_, _03178_);
  and (_04770_, _04769_, _04767_);
  and (_04771_, _04770_, _04765_);
  and (_04772_, _04771_, _04762_);
  and (_04773_, _04772_, _04758_);
  and (_04774_, _04773_, _04737_);
  and (_04775_, _04774_, _04731_);
  and (_04776_, _04775_, _04713_);
  nor (_04777_, _04500_, _04442_);
  and (_04778_, _04777_, _04776_);
  and (_04780_, _04778_, _04712_);
  nor (_04781_, _04482_, _04479_);
  nor (_04782_, _03714_, _03453_);
  and (_04783_, _04782_, _04246_);
  and (_04784_, _04783_, _04263_);
  nor (_04785_, _04784_, _03454_);
  nor (_04786_, _04785_, _04524_);
  and (_04787_, _04786_, _04781_);
  nor (_04788_, _04431_, _04410_);
  nor (_04789_, _04454_, _04421_);
  and (_04790_, _04789_, _04788_);
  and (_04791_, _04790_, _04787_);
  and (_04792_, _04791_, _04517_);
  and (_04793_, _04792_, _04780_);
  and (_04794_, _43868_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_04795_, _04794_);
  nor (_04796_, _04795_, _04793_);
  not (_04797_, _04796_);
  nor (_04798_, _04797_, _04711_);
  and (_04799_, _04798_, _04557_);
  not (_04800_, _03904_);
  and (_04801_, _03448_, _04800_);
  and (_04802_, _03861_, _03453_);
  and (_04803_, _03493_, _03197_);
  and (_04804_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04805_, _04804_, \oc8051_golden_model_1.SP [2]);
  nor (_04806_, _04804_, \oc8051_golden_model_1.SP [2]);
  nor (_04807_, _04806_, _04805_);
  and (_04808_, _04807_, _03188_);
  and (_04809_, _04500_, _04800_);
  and (_04810_, _03861_, _03505_);
  and (_04811_, _04807_, _03508_);
  and (_04812_, _04421_, _04800_);
  not (_04813_, _04807_);
  and (_04814_, _04813_, _03980_);
  and (_04815_, _03493_, _03609_);
  nor (_04816_, _04815_, _04814_);
  and (_04817_, _03904_, _04410_);
  not (_04818_, _04725_);
  not (_04819_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_04820_, _04261_, _04819_);
  not (_04821_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_04822_, _04348_, _04821_);
  and (_04823_, _04822_, _04346_);
  nand (_04824_, _04823_, _04820_);
  not (_04825_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_04826_, _04348_, _04825_);
  not (_04827_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_04828_, _04261_, _04827_);
  and (_04829_, _04828_, _04354_);
  nand (_04830_, _04829_, _04826_);
  nand (_04831_, _04830_, _04824_);
  nand (_04832_, _04831_, _04016_);
  not (_04833_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_04834_, _04348_, _04833_);
  not (_04835_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_04836_, _04261_, _04835_);
  and (_04837_, _04836_, _04354_);
  nand (_04838_, _04837_, _04834_);
  not (_04839_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_04840_, _04261_, _04839_);
  not (_04841_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_04842_, _04348_, _04841_);
  and (_04843_, _04842_, _04346_);
  nand (_04844_, _04843_, _04840_);
  nand (_04845_, _04844_, _04838_);
  nand (_04846_, _04845_, _04361_);
  nand (_04847_, _04846_, _04832_);
  nand (_04848_, _04847_, _03829_);
  not (_04849_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_04850_, _04348_, _04849_);
  not (_04851_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_04852_, _04261_, _04851_);
  and (_04853_, _04852_, _04354_);
  nand (_04854_, _04853_, _04850_);
  nand (_04855_, _04348_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_04856_, _04261_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_04857_, _04856_, _04346_);
  nand (_04858_, _04857_, _04855_);
  nand (_04859_, _04858_, _04854_);
  nand (_04860_, _04859_, _04016_);
  not (_04861_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_04862_, _04348_, _04861_);
  not (_04863_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_04864_, _04261_, _04863_);
  and (_04865_, _04864_, _04354_);
  nand (_04866_, _04865_, _04862_);
  nand (_04867_, _04348_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_04868_, _04261_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_04869_, _04868_, _04346_);
  nand (_04870_, _04869_, _04867_);
  nand (_04871_, _04870_, _04866_);
  nand (_04872_, _04871_, _04361_);
  nand (_04873_, _04872_, _04860_);
  nand (_04874_, _04873_, _04379_);
  nand (_04875_, _04874_, _04848_);
  nor (_04876_, _04875_, _03029_);
  nor (_04877_, _04876_, _04818_);
  nor (_04878_, _04877_, _04817_);
  and (_04879_, _04878_, _04816_);
  and (_04880_, _04875_, _04422_);
  nor (_04881_, _04880_, _04421_);
  and (_04882_, _04881_, _04879_);
  nor (_04883_, _04882_, _04812_);
  nor (_04884_, _04883_, _04428_);
  nor (_04885_, _04884_, _03862_);
  nor (_04886_, _04807_, _03230_);
  nor (_04887_, _04886_, _04885_);
  and (_04888_, _03493_, _03507_);
  and (_04889_, _04431_, _03904_);
  nor (_04890_, _04889_, _04888_);
  and (_04891_, _04890_, _04887_);
  and (_04892_, _04875_, _04443_);
  nor (_04893_, _04892_, _04442_);
  and (_04894_, _04893_, _04891_);
  and (_04895_, _04442_, _04800_);
  nor (_04896_, _04895_, _04894_);
  and (_04897_, _03860_, _04449_);
  nor (_04898_, _04897_, _04896_);
  and (_04899_, _04898_, _03510_);
  nor (_04900_, _04899_, _04811_);
  and (_04901_, _04454_, _03860_);
  or (_04902_, _04901_, _04900_);
  and (_04903_, _03493_, _03751_);
  nor (_04904_, _04807_, _03227_);
  nor (_04905_, _04904_, _04903_);
  not (_04906_, _04905_);
  nor (_04907_, _04906_, _04902_);
  and (_04908_, _04875_, _04463_);
  nor (_04909_, _04908_, _04462_);
  and (_04910_, _04909_, _04907_);
  nor (_04911_, _04910_, _04810_);
  nor (_04912_, _04911_, _03224_);
  and (_04913_, _04807_, _03224_);
  nor (_04914_, _04913_, _04912_);
  nor (_04915_, _04485_, _04800_);
  nor (_04916_, _04915_, _04716_);
  not (_04917_, _04916_);
  nor (_04918_, _04917_, _04914_);
  and (_04919_, _04875_, _04502_);
  nor (_04920_, _04919_, _04500_);
  and (_04921_, _04920_, _04918_);
  nor (_04922_, _04921_, _04809_);
  nor (_04923_, _04922_, _03178_);
  and (_04924_, _04807_, _03178_);
  nor (_04925_, _04924_, _04923_);
  nor (_04926_, _04517_, _04800_);
  nor (_04927_, _04926_, _03192_);
  not (_04928_, _04927_);
  nor (_04929_, _04928_, _04925_);
  and (_04930_, _04807_, _03192_);
  nor (_04931_, _04930_, _04929_);
  and (_04932_, _04524_, _03904_);
  or (_04933_, _04932_, _03188_);
  nor (_04934_, _04933_, _04931_);
  nor (_04935_, _04934_, _04808_);
  nor (_04936_, _04935_, _04803_);
  and (_04937_, _04875_, _04533_);
  nor (_04938_, _04937_, _04531_);
  and (_04939_, _04938_, _04936_);
  and (_04940_, _04531_, _04800_);
  nor (_04941_, _04940_, _04939_);
  nor (_04942_, _04807_, _04540_);
  nor (_04943_, _04942_, _04539_);
  not (_04944_, _04943_);
  nor (_04945_, _04944_, _04941_);
  nor (_04946_, _04945_, _04802_);
  nor (_04947_, _04946_, _04253_);
  and (_04948_, _04875_, _04552_);
  nor (_04949_, _04948_, _03448_);
  and (_04950_, _04949_, _04947_);
  nor (_04951_, _04950_, _04801_);
  not (_04952_, _04951_);
  not (_04953_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_04954_, _04261_, _04953_);
  not (_04955_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_04956_, _04348_, _04955_);
  and (_04957_, _04956_, _04346_);
  nand (_04958_, _04957_, _04954_);
  not (_04959_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_04960_, _04348_, _04959_);
  not (_04961_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_04962_, _04261_, _04961_);
  and (_04963_, _04962_, _04354_);
  nand (_04964_, _04963_, _04960_);
  nand (_04965_, _04964_, _04958_);
  nand (_04966_, _04965_, _04016_);
  not (_04967_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_04968_, _04348_, _04967_);
  not (_04969_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_04970_, _04261_, _04969_);
  and (_04971_, _04970_, _04354_);
  nand (_04972_, _04971_, _04968_);
  not (_04973_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_04974_, _04261_, _04973_);
  not (_04975_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_04976_, _04348_, _04975_);
  and (_04977_, _04976_, _04346_);
  nand (_04978_, _04977_, _04974_);
  nand (_04979_, _04978_, _04972_);
  nand (_04980_, _04979_, _04361_);
  nand (_04981_, _04980_, _04966_);
  nand (_04982_, _04981_, _03829_);
  nand (_04983_, _04261_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_04984_, _04348_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_04985_, _04984_, _04354_);
  nand (_04986_, _04985_, _04983_);
  nand (_04987_, _04348_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_04988_, _04261_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_04989_, _04988_, _04346_);
  nand (_04990_, _04989_, _04987_);
  nand (_04991_, _04990_, _04986_);
  nand (_04992_, _04991_, _04016_);
  nand (_04993_, _04261_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_04994_, _04348_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_04995_, _04994_, _04354_);
  nand (_04996_, _04995_, _04993_);
  nand (_04997_, _04348_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_04998_, _04261_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_04999_, _04998_, _04346_);
  nand (_05000_, _04999_, _04997_);
  nand (_05001_, _05000_, _04996_);
  nand (_05002_, _05001_, _04361_);
  nand (_05003_, _05002_, _04992_);
  nand (_05004_, _05003_, _04379_);
  nand (_05005_, _05004_, _04982_);
  and (_05006_, _05005_, _04502_);
  and (_05007_, _05005_, _04463_);
  nor (_05008_, _04805_, \oc8051_golden_model_1.SP [3]);
  and (_05009_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_05010_, _05009_, \oc8051_golden_model_1.SP [3]);
  and (_05011_, _05010_, \oc8051_golden_model_1.SP [0]);
  nor (_05012_, _05011_, _05008_);
  and (_05013_, _05012_, _04766_);
  and (_05014_, _03549_, _04428_);
  and (_05015_, _05005_, _04422_);
  and (_05016_, _05012_, _03980_);
  and (_05017_, _05005_, _03513_);
  not (_05018_, \oc8051_golden_model_1.PSW [3]);
  and (_05019_, _03240_, _05018_);
  nor (_05020_, _05019_, _04410_);
  not (_05021_, _05020_);
  nor (_05022_, _05021_, _05017_);
  and (_05023_, _04409_, _04051_);
  nor (_05024_, _05023_, _05022_);
  nor (_05025_, _05024_, _03980_);
  or (_05026_, _05025_, _04422_);
  nor (_05027_, _05026_, _05016_);
  or (_05028_, _05027_, _04421_);
  nor (_05029_, _05028_, _05015_);
  and (_05030_, _04421_, _03756_);
  or (_05031_, _05030_, _04428_);
  nor (_05032_, _05031_, _05029_);
  nor (_05033_, _05032_, _05014_);
  nor (_05034_, _05033_, _04768_);
  nor (_05035_, _05012_, _03230_);
  nor (_05036_, _05035_, _04431_);
  not (_05037_, _05036_);
  nor (_05038_, _05037_, _05034_);
  and (_05039_, _04431_, _03756_);
  nor (_05040_, _05039_, _04443_);
  not (_05041_, _05040_);
  nor (_05042_, _05041_, _05038_);
  and (_05043_, _05005_, _04443_);
  nor (_05044_, _05043_, _04442_);
  not (_05045_, _05044_);
  nor (_05046_, _05045_, _05042_);
  and (_05047_, _04442_, _03756_);
  or (_05048_, _05047_, _04449_);
  nor (_05049_, _05048_, _05046_);
  and (_05050_, _03549_, _04449_);
  nor (_05051_, _05050_, _05049_);
  and (_05052_, _05051_, _03510_);
  and (_05053_, _05012_, _03508_);
  nor (_05054_, _05053_, _05052_);
  nor (_05055_, _05054_, _04454_);
  nor (_05056_, _04562_, _03583_);
  or (_05057_, _05056_, _05055_);
  and (_05058_, _05057_, _03227_);
  or (_05059_, _05058_, _04463_);
  nor (_05060_, _05059_, _05013_);
  or (_05061_, _05060_, _04462_);
  nor (_05062_, _05061_, _05007_);
  not (_05063_, _04462_);
  nor (_05064_, _05063_, _03583_);
  nor (_05065_, _05064_, _05062_);
  nor (_05066_, _05065_, _03224_);
  and (_05067_, _05012_, _03224_);
  not (_05068_, _05067_);
  and (_05069_, _05068_, _04485_);
  not (_05070_, _05069_);
  nor (_05071_, _05070_, _05066_);
  nor (_05072_, _04485_, _03756_);
  nor (_05073_, _05072_, _05071_);
  nor (_05074_, _05073_, _04502_);
  or (_05075_, _05074_, _04500_);
  nor (_05076_, _05075_, _05006_);
  and (_05077_, _04500_, _03756_);
  nor (_05078_, _05077_, _05076_);
  nor (_05079_, _05078_, _03178_);
  and (_05080_, _05012_, _03178_);
  not (_05081_, _05080_);
  and (_05082_, _05081_, _04517_);
  not (_05083_, _05082_);
  nor (_05084_, _05083_, _05079_);
  nor (_05085_, _04517_, _03756_);
  nor (_05086_, _05085_, _03192_);
  not (_05087_, _05086_);
  nor (_05088_, _05087_, _05084_);
  and (_05089_, _05012_, _03192_);
  or (_05090_, _05089_, _04524_);
  nor (_05091_, _05090_, _05088_);
  and (_05092_, _04524_, _03581_);
  or (_05093_, _05092_, _03188_);
  nor (_05094_, _05093_, _05091_);
  and (_05095_, _05012_, _03188_);
  nor (_05096_, _05095_, _04533_);
  not (_05097_, _05096_);
  nor (_05098_, _05097_, _05094_);
  and (_05099_, _05005_, _04533_);
  nor (_05100_, _05099_, _04531_);
  not (_05101_, _05100_);
  nor (_05102_, _05101_, _05098_);
  not (_05103_, _04540_);
  and (_05104_, _04531_, _03756_);
  nor (_05105_, _05104_, _05103_);
  not (_05106_, _05105_);
  nor (_05107_, _05106_, _05102_);
  nor (_05108_, _05012_, _04540_);
  nor (_05109_, _05108_, _04539_);
  not (_05110_, _05109_);
  nor (_05111_, _05110_, _05107_);
  not (_05112_, _03549_);
  and (_05113_, _04539_, _05112_);
  nor (_05114_, _05113_, _04552_);
  not (_05115_, _05114_);
  nor (_05116_, _05115_, _05111_);
  and (_05117_, _05005_, _04552_);
  nor (_05118_, _05117_, _03448_);
  not (_05119_, _05118_);
  nor (_05120_, _05119_, _05116_);
  and (_05121_, _03827_, _03446_);
  nor (_05122_, _05121_, _05120_);
  nor (_05123_, _04797_, _05122_);
  and (_05124_, _05123_, _04952_);
  and (_05125_, _05124_, _04799_);
  or (_05126_, _05125_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_05127_, _05009_, _03498_);
  nor (_05128_, _04807_, _03499_);
  nor (_05129_, _05128_, _05127_);
  and (_05130_, _05127_, _03722_);
  nor (_05131_, _05010_, _05008_);
  nor (_05132_, _05131_, _05130_);
  not (_05133_, _05132_);
  and (_05134_, _04769_, _04763_);
  and (_05135_, _05134_, _04767_);
  and (_05136_, _05135_, _04735_);
  nor (_05137_, _05136_, _04795_);
  and (_05138_, _05137_, _05133_);
  and (_05139_, _05138_, _05129_);
  and (_05140_, _05139_, _03497_);
  not (_05141_, _05140_);
  and (_05142_, _05141_, _05126_);
  not (_05143_, _05125_);
  not (_05144_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_05145_, _04261_, _05144_);
  not (_05146_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_05147_, _04348_, _05146_);
  and (_05148_, _05147_, _04346_);
  nand (_05149_, _05148_, _05145_);
  not (_05150_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_05151_, _04348_, _05150_);
  not (_05152_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_05153_, _04261_, _05152_);
  and (_05154_, _05153_, _04354_);
  nand (_05155_, _05154_, _05151_);
  nand (_05156_, _05155_, _05149_);
  nand (_05157_, _05156_, _04016_);
  not (_05158_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_05159_, _04348_, _05158_);
  not (_05160_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_05161_, _04261_, _05160_);
  and (_05162_, _05161_, _04354_);
  nand (_05163_, _05162_, _05159_);
  not (_05164_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_05165_, _04261_, _05164_);
  not (_05166_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_05167_, _04348_, _05166_);
  and (_05168_, _05167_, _04346_);
  nand (_05169_, _05168_, _05165_);
  nand (_05170_, _05169_, _05163_);
  nand (_05171_, _05170_, _04361_);
  nand (_05172_, _05171_, _05157_);
  nand (_05173_, _05172_, _03829_);
  not (_05174_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_05175_, _04348_, _05174_);
  not (_05176_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_05177_, _04261_, _05176_);
  and (_05178_, _05177_, _04354_);
  nand (_05179_, _05178_, _05175_);
  not (_05180_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_05181_, _04261_, _05180_);
  not (_05182_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_05183_, _04348_, _05182_);
  and (_05184_, _05183_, _04346_);
  nand (_05185_, _05184_, _05181_);
  nand (_05186_, _05185_, _05179_);
  nand (_05187_, _05186_, _04016_);
  not (_05188_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_05189_, _04348_, _05188_);
  not (_05190_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_05191_, _04261_, _05190_);
  and (_05192_, _05191_, _04354_);
  nand (_05193_, _05192_, _05189_);
  not (_05194_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_05195_, _04261_, _05194_);
  not (_05196_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_05197_, _04348_, _05196_);
  and (_05198_, _05197_, _04346_);
  nand (_05199_, _05198_, _05195_);
  nand (_05200_, _05199_, _05193_);
  nand (_05201_, _05200_, _04361_);
  nand (_05202_, _05201_, _05187_);
  nand (_05203_, _05202_, _04379_);
  nand (_05204_, _05203_, _05173_);
  or (_05205_, _05204_, _03454_);
  and (_05206_, _03549_, _03454_);
  and (_05207_, _05206_, _03860_);
  and (_05208_, _05207_, _03486_);
  and (_05209_, _05208_, _03581_);
  nor (_05210_, _03414_, _04048_);
  and (_05211_, _05210_, _04800_);
  and (_05212_, _05211_, _05209_);
  and (_05213_, _05212_, \oc8051_golden_model_1.PCON [7]);
  not (_05214_, _05213_);
  and (_05215_, _03414_, _04188_);
  and (_05216_, _05215_, _03904_);
  and (_05217_, _05216_, _03756_);
  not (_05218_, _03486_);
  and (_05219_, _05218_, _03860_);
  and (_05220_, _05219_, _05206_);
  and (_05221_, _05220_, _05217_);
  and (_05222_, _05221_, \oc8051_golden_model_1.SBUF [7]);
  and (_05223_, _03414_, _04048_);
  and (_05224_, _05223_, _03904_);
  and (_05225_, _05224_, _03756_);
  not (_05226_, _03860_);
  and (_05227_, _03486_, _05226_);
  and (_05228_, _05227_, _05206_);
  and (_05229_, _05228_, _05225_);
  and (_05230_, _05229_, \oc8051_golden_model_1.IE [7]);
  nor (_05231_, _05230_, _05222_);
  and (_05232_, _05231_, _05214_);
  and (_05233_, _03904_, _03581_);
  and (_05234_, _05233_, _05223_);
  and (_05235_, _05234_, _05228_);
  and (_05236_, _05235_, \oc8051_golden_model_1.P2 [7]);
  nor (_05237_, _03486_, _03860_);
  and (_05238_, _05237_, _05206_);
  and (_05239_, _05238_, _05234_);
  and (_05240_, _05239_, \oc8051_golden_model_1.P3 [7]);
  nor (_05241_, _05240_, _05236_);
  and (_05242_, _05241_, _05232_);
  nor (_05243_, _03549_, _03446_);
  and (_05244_, _05243_, _05219_);
  and (_05245_, _05244_, _05234_);
  and (_05246_, _05245_, \oc8051_golden_model_1.PSW [7]);
  and (_05247_, _05243_, _05237_);
  and (_05248_, _05247_, _05234_);
  and (_05249_, _05248_, \oc8051_golden_model_1.B [7]);
  nor (_05250_, _05249_, _05246_);
  and (_05251_, _05238_, _05225_);
  and (_05252_, _05251_, \oc8051_golden_model_1.IP [7]);
  and (_05253_, _05243_, _05227_);
  and (_05254_, _05253_, _05234_);
  and (_05255_, _05254_, \oc8051_golden_model_1.ACC [7]);
  nor (_05256_, _05255_, _05252_);
  and (_05257_, _05256_, _05250_);
  and (_05258_, _05225_, _05208_);
  and (_05259_, _05258_, \oc8051_golden_model_1.TCON [7]);
  not (_05260_, _05208_);
  nor (_05261_, _03904_, _03581_);
  nand (_05262_, _05261_, _05223_);
  nor (_05263_, _05262_, _05260_);
  and (_05264_, _05263_, \oc8051_golden_model_1.TH0 [7]);
  nor (_05265_, _05264_, _05259_);
  and (_05266_, _05234_, _05220_);
  and (_05267_, _05266_, \oc8051_golden_model_1.P1 [7]);
  not (_05268_, _05210_);
  nand (_05269_, _03904_, _03756_);
  or (_05270_, _05269_, _05268_);
  nor (_05271_, _05270_, _05260_);
  and (_05272_, _05271_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05273_, _05272_, _05267_);
  and (_05274_, _05273_, _05265_);
  and (_05275_, _05225_, _05220_);
  and (_05276_, _05275_, \oc8051_golden_model_1.SCON [7]);
  nand (_05277_, _05261_, _05215_);
  nor (_05278_, _05277_, _05260_);
  and (_05279_, _05278_, \oc8051_golden_model_1.TH1 [7]);
  nor (_05280_, _05279_, _05276_);
  nor (_05281_, _03414_, _04188_);
  not (_05282_, _05281_);
  or (_05283_, _05282_, _05269_);
  nor (_05284_, _05283_, _05260_);
  and (_05285_, _05284_, \oc8051_golden_model_1.TL0 [7]);
  and (_05286_, _05217_, _05208_);
  and (_05287_, _05286_, \oc8051_golden_model_1.TMOD [7]);
  nor (_05288_, _05287_, _05285_);
  and (_05289_, _05288_, _05280_);
  and (_05290_, _05289_, _05274_);
  and (_05291_, _05290_, _05257_);
  and (_05292_, _05291_, _05242_);
  and (_05293_, _05234_, _05208_);
  and (_05294_, _05293_, \oc8051_golden_model_1.P0 [7]);
  not (_05295_, _05294_);
  and (_05296_, _05210_, _03904_);
  and (_05297_, _05296_, _05209_);
  and (_05298_, _05297_, \oc8051_golden_model_1.DPH [7]);
  not (_05299_, _05298_);
  and (_05300_, _05216_, _05209_);
  and (_05301_, _05300_, \oc8051_golden_model_1.SP [7]);
  and (_05302_, _05281_, _03904_);
  and (_05303_, _05302_, _05209_);
  and (_05304_, _05303_, \oc8051_golden_model_1.DPL [7]);
  nor (_05305_, _05304_, _05301_);
  and (_05306_, _05305_, _05299_);
  and (_05307_, _05306_, _05295_);
  and (_05308_, _05307_, _05292_);
  and (_05309_, _05308_, _05205_);
  not (_05310_, _05309_);
  not (_05311_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_05312_, _04261_, _05311_);
  not (_05313_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_05314_, _04348_, _05313_);
  and (_05315_, _05314_, _04346_);
  nand (_05316_, _05315_, _05312_);
  not (_05317_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_05318_, _04348_, _05317_);
  not (_05319_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_05320_, _04261_, _05319_);
  and (_05321_, _05320_, _04354_);
  nand (_05322_, _05321_, _05318_);
  nand (_05323_, _05322_, _05316_);
  nand (_05324_, _05323_, _04016_);
  not (_05325_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_05326_, _04348_, _05325_);
  not (_05327_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_05328_, _04261_, _05327_);
  and (_05329_, _05328_, _04354_);
  nand (_05330_, _05329_, _05326_);
  not (_05331_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_05332_, _04261_, _05331_);
  not (_05333_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_05334_, _04348_, _05333_);
  and (_05335_, _05334_, _04346_);
  nand (_05336_, _05335_, _05332_);
  nand (_05337_, _05336_, _05330_);
  nand (_05338_, _05337_, _04361_);
  nand (_05339_, _05338_, _05324_);
  nand (_05340_, _05339_, _03829_);
  nand (_05341_, _04261_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_05342_, _04348_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_05343_, _05342_, _04354_);
  nand (_05344_, _05343_, _05341_);
  nand (_05345_, _04348_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_05346_, _04261_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_05347_, _05346_, _04346_);
  nand (_05348_, _05347_, _05345_);
  nand (_05349_, _05348_, _05344_);
  nand (_05350_, _05349_, _04016_);
  nand (_05351_, _04261_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_05352_, _04348_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_05353_, _05352_, _04354_);
  nand (_05354_, _05353_, _05351_);
  nand (_05355_, _04348_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_05356_, _04261_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_05357_, _05356_, _04346_);
  nand (_05358_, _05357_, _05355_);
  nand (_05359_, _05358_, _05354_);
  nand (_05360_, _05359_, _04361_);
  nand (_05361_, _05360_, _05350_);
  nand (_05362_, _05361_, _04379_);
  nand (_05363_, _05362_, _05340_);
  or (_05364_, _05363_, _03454_);
  and (_05365_, _05297_, \oc8051_golden_model_1.DPH [6]);
  not (_05366_, _05365_);
  and (_05367_, _05263_, \oc8051_golden_model_1.TH0 [6]);
  and (_05368_, _05271_, \oc8051_golden_model_1.TL1 [6]);
  nor (_05369_, _05368_, _05367_);
  and (_05370_, _05369_, _05366_);
  and (_05371_, _05300_, \oc8051_golden_model_1.SP [6]);
  and (_05372_, _05303_, \oc8051_golden_model_1.DPL [6]);
  nor (_05373_, _05372_, _05371_);
  and (_05374_, _05212_, \oc8051_golden_model_1.PCON [6]);
  not (_05375_, _05374_);
  and (_05376_, _05221_, \oc8051_golden_model_1.SBUF [6]);
  and (_05377_, _05229_, \oc8051_golden_model_1.IE [6]);
  nor (_05378_, _05377_, _05376_);
  and (_05379_, _05378_, _05375_);
  and (_05380_, _05379_, _05373_);
  and (_05381_, _05380_, _05370_);
  and (_05382_, _05284_, \oc8051_golden_model_1.TL0 [6]);
  and (_05383_, _05275_, \oc8051_golden_model_1.SCON [6]);
  nor (_05384_, _05383_, _05382_);
  and (_05385_, _05278_, \oc8051_golden_model_1.TH1 [6]);
  not (_05386_, _05385_);
  and (_05387_, _05258_, \oc8051_golden_model_1.TCON [6]);
  and (_05388_, _05286_, \oc8051_golden_model_1.TMOD [6]);
  nor (_05389_, _05388_, _05387_);
  and (_05390_, _05389_, _05386_);
  and (_05391_, _05390_, _05384_);
  and (_05392_, _05251_, \oc8051_golden_model_1.IP [6]);
  and (_05393_, _05248_, \oc8051_golden_model_1.B [6]);
  nor (_05394_, _05393_, _05392_);
  and (_05395_, _05245_, \oc8051_golden_model_1.PSW [6]);
  and (_05396_, _05254_, \oc8051_golden_model_1.ACC [6]);
  nor (_05397_, _05396_, _05395_);
  and (_05398_, _05397_, _05394_);
  and (_05399_, _05293_, \oc8051_golden_model_1.P0 [6]);
  not (_05400_, _05399_);
  and (_05401_, _05266_, \oc8051_golden_model_1.P1 [6]);
  not (_05402_, _05401_);
  and (_05403_, _05235_, \oc8051_golden_model_1.P2 [6]);
  and (_05404_, _05239_, \oc8051_golden_model_1.P3 [6]);
  nor (_05405_, _05404_, _05403_);
  and (_05406_, _05405_, _05402_);
  and (_05407_, _05406_, _05400_);
  and (_05408_, _05407_, _05398_);
  and (_05409_, _05408_, _05391_);
  and (_05410_, _05409_, _05381_);
  and (_05411_, _05410_, _05364_);
  not (_05412_, _05411_);
  not (_05413_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_05414_, _04261_, _05413_);
  not (_05415_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_05416_, _04348_, _05415_);
  and (_05417_, _05416_, _04346_);
  nand (_05418_, _05417_, _05414_);
  not (_05419_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_05420_, _04348_, _05419_);
  not (_05421_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_05422_, _04261_, _05421_);
  and (_05423_, _05422_, _04354_);
  nand (_05424_, _05423_, _05420_);
  nand (_05425_, _05424_, _05418_);
  nand (_05426_, _05425_, _04016_);
  not (_05427_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_05428_, _04348_, _05427_);
  not (_05429_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_05430_, _04261_, _05429_);
  and (_05431_, _05430_, _04354_);
  nand (_05432_, _05431_, _05428_);
  not (_05433_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_05434_, _04261_, _05433_);
  not (_05435_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_05436_, _04348_, _05435_);
  and (_05437_, _05436_, _04346_);
  nand (_05438_, _05437_, _05434_);
  nand (_05439_, _05438_, _05432_);
  nand (_05440_, _05439_, _04361_);
  nand (_05441_, _05440_, _05426_);
  nand (_05442_, _05441_, _03829_);
  nand (_05443_, _04261_, \oc8051_golden_model_1.IRAM[11] [5]);
  not (_05444_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_05445_, _04261_, _05444_);
  and (_05446_, _05445_, _04354_);
  nand (_05447_, _05446_, _05443_);
  nand (_05448_, _04348_, \oc8051_golden_model_1.IRAM[8] [5]);
  not (_05449_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_05450_, _04348_, _05449_);
  and (_05451_, _05450_, _04346_);
  nand (_05452_, _05451_, _05448_);
  nand (_05453_, _05452_, _05447_);
  nand (_05454_, _05453_, _04016_);
  nand (_05455_, _04261_, \oc8051_golden_model_1.IRAM[15] [5]);
  not (_05456_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_05457_, _04261_, _05456_);
  and (_05458_, _05457_, _04354_);
  nand (_05459_, _05458_, _05455_);
  nand (_05460_, _04348_, \oc8051_golden_model_1.IRAM[12] [5]);
  not (_05461_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_05462_, _04348_, _05461_);
  and (_05463_, _05462_, _04346_);
  nand (_05464_, _05463_, _05460_);
  nand (_05465_, _05464_, _05459_);
  nand (_05466_, _05465_, _04361_);
  nand (_05467_, _05466_, _05454_);
  nand (_05468_, _05467_, _04379_);
  nand (_05469_, _05468_, _05442_);
  or (_05470_, _05469_, _03454_);
  and (_05471_, _05297_, \oc8051_golden_model_1.DPH [5]);
  not (_05472_, _05471_);
  and (_05473_, _05300_, \oc8051_golden_model_1.SP [5]);
  and (_05474_, _05303_, \oc8051_golden_model_1.DPL [5]);
  nor (_05475_, _05474_, _05473_);
  and (_05476_, _05475_, _05472_);
  and (_05477_, _05258_, \oc8051_golden_model_1.TCON [5]);
  not (_05478_, _05477_);
  and (_05479_, _05284_, \oc8051_golden_model_1.TL0 [5]);
  and (_05480_, _05275_, \oc8051_golden_model_1.SCON [5]);
  nor (_05481_, _05480_, _05479_);
  and (_05482_, _05481_, _05478_);
  and (_05483_, _05263_, \oc8051_golden_model_1.TH0 [5]);
  and (_05484_, _05278_, \oc8051_golden_model_1.TH1 [5]);
  nor (_05485_, _05484_, _05483_);
  and (_05486_, _05286_, \oc8051_golden_model_1.TMOD [5]);
  and (_05487_, _05271_, \oc8051_golden_model_1.TL1 [5]);
  nor (_05488_, _05487_, _05486_);
  and (_05489_, _05488_, _05485_);
  and (_05490_, _05489_, _05482_);
  and (_05491_, _05490_, _05476_);
  and (_05492_, _05212_, \oc8051_golden_model_1.PCON [5]);
  not (_05493_, _05492_);
  and (_05494_, _05221_, \oc8051_golden_model_1.SBUF [5]);
  and (_05495_, _05229_, \oc8051_golden_model_1.IE [5]);
  nor (_05496_, _05495_, _05494_);
  and (_05497_, _05496_, _05493_);
  and (_05498_, _05293_, \oc8051_golden_model_1.P0 [5]);
  not (_05499_, _05498_);
  and (_05500_, _05245_, \oc8051_golden_model_1.PSW [5]);
  and (_05501_, _05254_, \oc8051_golden_model_1.ACC [5]);
  nor (_05502_, _05501_, _05500_);
  and (_05503_, _05251_, \oc8051_golden_model_1.IP [5]);
  and (_05504_, _05248_, \oc8051_golden_model_1.B [5]);
  nor (_05505_, _05504_, _05503_);
  and (_05506_, _05505_, _05502_);
  and (_05507_, _05266_, \oc8051_golden_model_1.P1 [5]);
  not (_05508_, _05507_);
  and (_05509_, _05235_, \oc8051_golden_model_1.P2 [5]);
  and (_05510_, _05239_, \oc8051_golden_model_1.P3 [5]);
  nor (_05511_, _05510_, _05509_);
  and (_05512_, _05511_, _05508_);
  and (_05513_, _05512_, _05506_);
  and (_05514_, _05513_, _05499_);
  and (_05515_, _05514_, _05497_);
  and (_05516_, _05515_, _05491_);
  and (_05517_, _05516_, _05470_);
  not (_05518_, _05517_);
  or (_05519_, _05005_, _03454_);
  and (_05520_, _05297_, \oc8051_golden_model_1.DPH [3]);
  not (_05521_, _05520_);
  and (_05522_, _05300_, \oc8051_golden_model_1.SP [3]);
  and (_05523_, _05303_, \oc8051_golden_model_1.DPL [3]);
  nor (_05524_, _05523_, _05522_);
  and (_05525_, _05524_, _05521_);
  and (_05526_, _05258_, \oc8051_golden_model_1.TCON [3]);
  not (_05527_, _05526_);
  and (_05528_, _05284_, \oc8051_golden_model_1.TL0 [3]);
  and (_05529_, _05275_, \oc8051_golden_model_1.SCON [3]);
  nor (_05530_, _05529_, _05528_);
  and (_05531_, _05530_, _05527_);
  and (_05532_, _05263_, \oc8051_golden_model_1.TH0 [3]);
  and (_05533_, _05278_, \oc8051_golden_model_1.TH1 [3]);
  nor (_05534_, _05533_, _05532_);
  and (_05535_, _05286_, \oc8051_golden_model_1.TMOD [3]);
  and (_05536_, _05271_, \oc8051_golden_model_1.TL1 [3]);
  nor (_05537_, _05536_, _05535_);
  and (_05538_, _05537_, _05534_);
  and (_05539_, _05538_, _05531_);
  and (_05540_, _05539_, _05525_);
  and (_05541_, _05212_, \oc8051_golden_model_1.PCON [3]);
  not (_05542_, _05541_);
  and (_05543_, _05221_, \oc8051_golden_model_1.SBUF [3]);
  and (_05544_, _05229_, \oc8051_golden_model_1.IE [3]);
  nor (_05545_, _05544_, _05543_);
  and (_05546_, _05545_, _05542_);
  and (_05547_, _05293_, \oc8051_golden_model_1.P0 [3]);
  not (_05548_, _05547_);
  and (_05549_, _05245_, \oc8051_golden_model_1.PSW [3]);
  and (_05550_, _05248_, \oc8051_golden_model_1.B [3]);
  nor (_05551_, _05550_, _05549_);
  and (_05552_, _05251_, \oc8051_golden_model_1.IP [3]);
  and (_05553_, _05254_, \oc8051_golden_model_1.ACC [3]);
  nor (_05554_, _05553_, _05552_);
  and (_05555_, _05554_, _05551_);
  and (_05556_, _05266_, \oc8051_golden_model_1.P1 [3]);
  not (_05557_, _05556_);
  and (_05558_, _05235_, \oc8051_golden_model_1.P2 [3]);
  and (_05559_, _05239_, \oc8051_golden_model_1.P3 [3]);
  nor (_05560_, _05559_, _05558_);
  and (_05561_, _05560_, _05557_);
  and (_05562_, _05561_, _05555_);
  and (_05563_, _05562_, _05548_);
  and (_05564_, _05563_, _05546_);
  and (_05565_, _05564_, _05540_);
  and (_05566_, _05565_, _05519_);
  not (_05567_, _05566_);
  or (_05568_, _04406_, _03454_);
  and (_05569_, _05300_, \oc8051_golden_model_1.SP [1]);
  not (_05570_, _05569_);
  and (_05571_, _05303_, \oc8051_golden_model_1.DPL [1]);
  and (_05572_, _05258_, \oc8051_golden_model_1.TCON [1]);
  nor (_05573_, _05572_, _05571_);
  and (_05574_, _05573_, _05570_);
  and (_05575_, _05293_, \oc8051_golden_model_1.P0 [1]);
  not (_05576_, _05575_);
  and (_05577_, _05266_, \oc8051_golden_model_1.P1 [1]);
  not (_05578_, _05577_);
  and (_05579_, _05235_, \oc8051_golden_model_1.P2 [1]);
  and (_05580_, _05239_, \oc8051_golden_model_1.P3 [1]);
  nor (_05581_, _05580_, _05579_);
  and (_05582_, _05581_, _05578_);
  and (_05583_, _05582_, _05576_);
  and (_05584_, _05583_, _05574_);
  and (_05585_, _05271_, \oc8051_golden_model_1.TL1 [1]);
  and (_05586_, _05278_, \oc8051_golden_model_1.TH1 [1]);
  nor (_05587_, _05586_, _05585_);
  and (_05588_, _05286_, \oc8051_golden_model_1.TMOD [1]);
  and (_05589_, _05275_, \oc8051_golden_model_1.SCON [1]);
  nor (_05590_, _05589_, _05588_);
  and (_05591_, _05590_, _05587_);
  and (_05592_, _05297_, \oc8051_golden_model_1.DPH [1]);
  not (_05593_, _05592_);
  and (_05594_, _05284_, \oc8051_golden_model_1.TL0 [1]);
  and (_05595_, _05263_, \oc8051_golden_model_1.TH0 [1]);
  nor (_05596_, _05595_, _05594_);
  and (_05597_, _05596_, _05593_);
  and (_05598_, _05597_, _05591_);
  and (_05599_, _05212_, \oc8051_golden_model_1.PCON [1]);
  not (_05600_, _05599_);
  and (_05601_, _05251_, \oc8051_golden_model_1.IP [1]);
  not (_05602_, _05601_);
  and (_05603_, _05245_, \oc8051_golden_model_1.PSW [1]);
  and (_05604_, _05248_, \oc8051_golden_model_1.B [1]);
  nor (_05605_, _05604_, _05603_);
  and (_05606_, _05605_, _05602_);
  and (_05607_, _05221_, \oc8051_golden_model_1.SBUF [1]);
  not (_05608_, _05607_);
  and (_05609_, _05229_, \oc8051_golden_model_1.IE [1]);
  and (_05610_, _05254_, \oc8051_golden_model_1.ACC [1]);
  nor (_05611_, _05610_, _05609_);
  and (_05612_, _05611_, _05608_);
  and (_05613_, _05612_, _05606_);
  and (_05614_, _05613_, _05600_);
  and (_05615_, _05614_, _05598_);
  and (_05616_, _05615_, _05584_);
  and (_05617_, _05616_, _05568_);
  not (_05618_, _05617_);
  or (_05619_, _04634_, _03454_);
  and (_05620_, _05297_, \oc8051_golden_model_1.DPH [0]);
  not (_05621_, _05620_);
  and (_05622_, _05300_, \oc8051_golden_model_1.SP [0]);
  and (_05623_, _05303_, \oc8051_golden_model_1.DPL [0]);
  nor (_05624_, _05623_, _05622_);
  and (_05625_, _05624_, _05621_);
  and (_05626_, _05258_, \oc8051_golden_model_1.TCON [0]);
  not (_05627_, _05626_);
  and (_05628_, _05284_, \oc8051_golden_model_1.TL0 [0]);
  and (_05629_, _05275_, \oc8051_golden_model_1.SCON [0]);
  nor (_05630_, _05629_, _05628_);
  and (_05631_, _05630_, _05627_);
  and (_05632_, _05263_, \oc8051_golden_model_1.TH0 [0]);
  and (_05633_, _05278_, \oc8051_golden_model_1.TH1 [0]);
  nor (_05634_, _05633_, _05632_);
  and (_05635_, _05286_, \oc8051_golden_model_1.TMOD [0]);
  and (_05636_, _05271_, \oc8051_golden_model_1.TL1 [0]);
  nor (_05637_, _05636_, _05635_);
  and (_05638_, _05637_, _05634_);
  and (_05639_, _05638_, _05631_);
  and (_05640_, _05639_, _05625_);
  and (_05641_, _05212_, \oc8051_golden_model_1.PCON [0]);
  not (_05642_, _05641_);
  and (_05643_, _05221_, \oc8051_golden_model_1.SBUF [0]);
  and (_05644_, _05229_, \oc8051_golden_model_1.IE [0]);
  nor (_05645_, _05644_, _05643_);
  and (_05646_, _05645_, _05642_);
  and (_05647_, _05293_, \oc8051_golden_model_1.P0 [0]);
  not (_05648_, _05647_);
  and (_05649_, _05251_, \oc8051_golden_model_1.IP [0]);
  and (_05650_, _05248_, \oc8051_golden_model_1.B [0]);
  nor (_05651_, _05650_, _05649_);
  and (_05652_, _05245_, \oc8051_golden_model_1.PSW [0]);
  and (_05653_, _05254_, \oc8051_golden_model_1.ACC [0]);
  nor (_05654_, _05653_, _05652_);
  and (_05655_, _05654_, _05651_);
  and (_05656_, _05266_, \oc8051_golden_model_1.P1 [0]);
  not (_05657_, _05656_);
  and (_05658_, _05235_, \oc8051_golden_model_1.P2 [0]);
  and (_05659_, _05239_, \oc8051_golden_model_1.P3 [0]);
  nor (_05660_, _05659_, _05658_);
  and (_05661_, _05660_, _05657_);
  and (_05662_, _05661_, _05655_);
  and (_05663_, _05662_, _05648_);
  and (_05664_, _05663_, _05646_);
  and (_05665_, _05664_, _05640_);
  nand (_05666_, _05665_, _05619_);
  and (_05667_, _05666_, _05618_);
  or (_05668_, _04875_, _03454_);
  and (_05669_, _05300_, \oc8051_golden_model_1.SP [2]);
  not (_05670_, _05669_);
  and (_05671_, _05303_, \oc8051_golden_model_1.DPL [2]);
  and (_05672_, _05258_, \oc8051_golden_model_1.TCON [2]);
  nor (_05673_, _05672_, _05671_);
  and (_05674_, _05673_, _05670_);
  and (_05675_, _05293_, \oc8051_golden_model_1.P0 [2]);
  not (_05676_, _05675_);
  and (_05677_, _05266_, \oc8051_golden_model_1.P1 [2]);
  not (_05678_, _05677_);
  and (_05679_, _05235_, \oc8051_golden_model_1.P2 [2]);
  and (_05680_, _05239_, \oc8051_golden_model_1.P3 [2]);
  nor (_05681_, _05680_, _05679_);
  and (_05682_, _05681_, _05678_);
  and (_05683_, _05682_, _05676_);
  and (_05684_, _05683_, _05674_);
  and (_05685_, _05271_, \oc8051_golden_model_1.TL1 [2]);
  and (_05686_, _05278_, \oc8051_golden_model_1.TH1 [2]);
  nor (_05687_, _05686_, _05685_);
  and (_05688_, _05286_, \oc8051_golden_model_1.TMOD [2]);
  and (_05689_, _05275_, \oc8051_golden_model_1.SCON [2]);
  nor (_05690_, _05689_, _05688_);
  and (_05691_, _05690_, _05687_);
  and (_05692_, _05297_, \oc8051_golden_model_1.DPH [2]);
  not (_05693_, _05692_);
  and (_05694_, _05284_, \oc8051_golden_model_1.TL0 [2]);
  and (_05695_, _05263_, \oc8051_golden_model_1.TH0 [2]);
  nor (_05696_, _05695_, _05694_);
  and (_05697_, _05696_, _05693_);
  and (_05698_, _05697_, _05691_);
  and (_05699_, _05212_, \oc8051_golden_model_1.PCON [2]);
  not (_05700_, _05699_);
  and (_05701_, _05251_, \oc8051_golden_model_1.IP [2]);
  not (_05702_, _05701_);
  and (_05703_, _05245_, \oc8051_golden_model_1.PSW [2]);
  and (_05704_, _05254_, \oc8051_golden_model_1.ACC [2]);
  nor (_05705_, _05704_, _05703_);
  and (_05706_, _05705_, _05702_);
  and (_05707_, _05221_, \oc8051_golden_model_1.SBUF [2]);
  not (_05708_, _05707_);
  and (_05709_, _05229_, \oc8051_golden_model_1.IE [2]);
  and (_05710_, _05248_, \oc8051_golden_model_1.B [2]);
  nor (_05711_, _05710_, _05709_);
  and (_05712_, _05711_, _05708_);
  and (_05713_, _05712_, _05706_);
  and (_05714_, _05713_, _05700_);
  and (_05715_, _05714_, _05698_);
  and (_05716_, _05715_, _05684_);
  and (_05717_, _05716_, _05668_);
  not (_05718_, _05717_);
  and (_05719_, _05718_, _05667_);
  and (_05720_, _05719_, _05567_);
  not (_05721_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_05722_, _04261_, _05721_);
  not (_05723_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_05724_, _04348_, _05723_);
  and (_05725_, _05724_, _04346_);
  nand (_05726_, _05725_, _05722_);
  not (_05727_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_05728_, _04348_, _05727_);
  not (_05729_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05730_, _04261_, _05729_);
  and (_05731_, _05730_, _04354_);
  nand (_05732_, _05731_, _05728_);
  nand (_05733_, _05732_, _05726_);
  nand (_05734_, _05733_, _04016_);
  not (_05735_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_05736_, _04348_, _05735_);
  not (_05737_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05738_, _04261_, _05737_);
  and (_05739_, _05738_, _04354_);
  nand (_05740_, _05739_, _05736_);
  not (_05741_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_05742_, _04261_, _05741_);
  not (_05743_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_05744_, _04348_, _05743_);
  and (_05745_, _05744_, _04346_);
  nand (_05746_, _05745_, _05742_);
  nand (_05747_, _05746_, _05740_);
  nand (_05748_, _05747_, _04361_);
  nand (_05749_, _05748_, _05734_);
  nand (_05750_, _05749_, _03829_);
  nand (_05751_, _04261_, \oc8051_golden_model_1.IRAM[11] [4]);
  not (_05752_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_05753_, _04261_, _05752_);
  and (_05754_, _05753_, _04354_);
  nand (_05755_, _05754_, _05751_);
  nand (_05756_, _04348_, \oc8051_golden_model_1.IRAM[8] [4]);
  not (_05757_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_05758_, _04348_, _05757_);
  and (_05759_, _05758_, _04346_);
  nand (_05760_, _05759_, _05756_);
  nand (_05761_, _05760_, _05755_);
  nand (_05762_, _05761_, _04016_);
  nand (_05763_, _04261_, \oc8051_golden_model_1.IRAM[15] [4]);
  not (_05764_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_05765_, _04261_, _05764_);
  and (_05766_, _05765_, _04354_);
  nand (_05767_, _05766_, _05763_);
  nand (_05768_, _04348_, \oc8051_golden_model_1.IRAM[12] [4]);
  not (_05769_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_05770_, _04348_, _05769_);
  and (_05771_, _05770_, _04346_);
  nand (_05772_, _05771_, _05768_);
  nand (_05773_, _05772_, _05767_);
  nand (_05774_, _05773_, _04361_);
  nand (_05775_, _05774_, _05762_);
  nand (_05776_, _05775_, _04379_);
  nand (_05777_, _05776_, _05750_);
  or (_05778_, _05777_, _03454_);
  and (_05779_, _05278_, \oc8051_golden_model_1.TH1 [4]);
  and (_05780_, _05221_, \oc8051_golden_model_1.SBUF [4]);
  nor (_05781_, _05780_, _05779_);
  and (_05782_, _05286_, \oc8051_golden_model_1.TMOD [4]);
  and (_05783_, _05275_, \oc8051_golden_model_1.SCON [4]);
  nor (_05784_, _05783_, _05782_);
  and (_05785_, _05784_, _05781_);
  and (_05786_, _05303_, \oc8051_golden_model_1.DPL [4]);
  not (_05787_, _05786_);
  and (_05788_, _05284_, \oc8051_golden_model_1.TL0 [4]);
  and (_05789_, _05229_, \oc8051_golden_model_1.IE [4]);
  nor (_05790_, _05789_, _05788_);
  and (_05791_, _05790_, _05787_);
  and (_05792_, _05300_, \oc8051_golden_model_1.SP [4]);
  and (_05793_, _05297_, \oc8051_golden_model_1.DPH [4]);
  nor (_05794_, _05793_, _05792_);
  and (_05795_, _05794_, _05791_);
  and (_05796_, _05795_, _05785_);
  not (_05797_, _05796_);
  and (_05798_, _05266_, \oc8051_golden_model_1.P1 [4]);
  and (_05799_, _05258_, \oc8051_golden_model_1.TCON [4]);
  and (_05800_, _05235_, \oc8051_golden_model_1.P2 [4]);
  and (_05801_, _05239_, \oc8051_golden_model_1.P3 [4]);
  or (_05802_, _05801_, _05800_);
  or (_05803_, _05802_, _05799_);
  or (_05804_, _05803_, _05798_);
  and (_05805_, _05212_, \oc8051_golden_model_1.PCON [4]);
  not (_05806_, _05805_);
  and (_05807_, _05245_, \oc8051_golden_model_1.PSW [4]);
  and (_05808_, _05248_, \oc8051_golden_model_1.B [4]);
  nor (_05809_, _05808_, _05807_);
  and (_05810_, _05251_, \oc8051_golden_model_1.IP [4]);
  and (_05811_, _05254_, \oc8051_golden_model_1.ACC [4]);
  nor (_05812_, _05811_, _05810_);
  and (_05813_, _05812_, _05809_);
  and (_05814_, _05813_, _05806_);
  and (_05815_, _05293_, \oc8051_golden_model_1.P0 [4]);
  not (_05816_, _05815_);
  and (_05817_, _05263_, \oc8051_golden_model_1.TH0 [4]);
  and (_05818_, _05271_, \oc8051_golden_model_1.TL1 [4]);
  nor (_05819_, _05818_, _05817_);
  and (_05820_, _05819_, _05816_);
  nand (_05821_, _05820_, _05814_);
  or (_05822_, _05821_, _05804_);
  nor (_05823_, _05822_, _05797_);
  and (_05824_, _05823_, _05778_);
  not (_05825_, _05824_);
  and (_05826_, _05825_, _05720_);
  and (_05827_, _05826_, _05518_);
  and (_05828_, _05827_, _05412_);
  nor (_05829_, _05828_, _05310_);
  and (_05830_, _05828_, _05310_);
  nor (_05831_, _05830_, _05829_);
  and (_05832_, _05831_, _03448_);
  not (_05833_, _05204_);
  and (_05834_, _05777_, _05469_);
  and (_05835_, _04406_, _04634_);
  and (_05836_, _04875_, _05005_);
  and (_05837_, _05836_, _05835_);
  and (_05838_, _05837_, _05834_);
  and (_05839_, _05838_, _05363_);
  or (_05840_, _05839_, _05833_);
  nand (_05841_, _05839_, _05833_);
  and (_05842_, _05841_, _05840_);
  and (_05843_, _03595_, _03197_);
  nor (_05844_, _04322_, _05843_);
  and (_05845_, _04474_, _03197_);
  not (_05846_, _05845_);
  and (_05847_, _05846_, _05844_);
  and (_05848_, _05847_, _04745_);
  or (_05849_, _05848_, _05842_);
  not (_05850_, _04511_);
  and (_05851_, _03654_, _01716_);
  and (_05852_, _03657_, _01688_);
  nor (_05853_, _05852_, _05851_);
  and (_05854_, _03685_, _01719_);
  and (_05855_, _03698_, _01673_);
  nor (_05856_, _05855_, _05854_);
  and (_05857_, _05856_, _05853_);
  and (_05858_, _03701_, _01663_);
  and (_05859_, _03703_, _01632_);
  nor (_05860_, _05859_, _05858_);
  and (_05861_, _03672_, _01697_);
  and (_05862_, _03678_, _01735_);
  nor (_05863_, _05862_, _05861_);
  and (_05864_, _05863_, _05860_);
  and (_05865_, _05864_, _05857_);
  and (_05866_, _03662_, _01708_);
  and (_05867_, _03692_, _01723_);
  nor (_05868_, _05867_, _05866_);
  and (_05869_, _03687_, _01731_);
  and (_05870_, _03690_, _01704_);
  nor (_05871_, _05870_, _05869_);
  and (_05872_, _05871_, _05868_);
  and (_05873_, _03675_, _01713_);
  and (_05874_, _03680_, _01668_);
  nor (_05875_, _05874_, _05873_);
  and (_05876_, _03696_, _01678_);
  and (_05877_, _03665_, _01684_);
  nor (_05878_, _05877_, _05876_);
  and (_05879_, _05878_, _05875_);
  and (_05880_, _05879_, _05872_);
  and (_05881_, _05880_, _05865_);
  and (_05882_, _05881_, _05309_);
  nor (_05883_, _05881_, _05309_);
  nor (_05884_, _05883_, _05882_);
  and (_05885_, _05884_, _04512_);
  not (_05886_, _03601_);
  not (_05887_, _04754_);
  not (_05888_, _04502_);
  nor (_05889_, _04717_, _04714_);
  and (_05890_, _03494_, _03176_);
  nor (_05891_, _05890_, _04493_);
  and (_05892_, _05891_, _05889_);
  and (_05893_, _05892_, _05888_);
  and (_05894_, _05893_, _05887_);
  and (_05895_, _05894_, _05886_);
  or (_05896_, _05895_, _03454_);
  not (_05897_, _03224_);
  nor (_05898_, _03487_, _04051_);
  and (_05899_, _03864_, _03583_);
  and (_05900_, _05899_, _05898_);
  and (_05901_, _05244_, _05900_);
  and (_05902_, _05901_, \oc8051_golden_model_1.PSW [7]);
  and (_05903_, _05253_, _05900_);
  and (_05904_, _05903_, \oc8051_golden_model_1.ACC [7]);
  nor (_05905_, _05904_, _05902_);
  nor (_05906_, _03861_, _03583_);
  and (_05907_, _05906_, _05898_);
  and (_05908_, _05907_, _05238_);
  and (_05909_, _05908_, \oc8051_golden_model_1.IP [7]);
  and (_05910_, _05247_, _05900_);
  and (_05911_, _05910_, \oc8051_golden_model_1.B [7]);
  nor (_05912_, _05911_, _05909_);
  and (_05913_, _05912_, _05905_);
  and (_05914_, _05209_, \oc8051_golden_model_1.P0INREG [7]);
  not (_05915_, _05914_);
  and (_05916_, _05220_, _05900_);
  and (_05917_, _05916_, \oc8051_golden_model_1.P1INREG [7]);
  and (_05918_, _05228_, _05900_);
  and (_05919_, _05918_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_05920_, _05919_, _05917_);
  and (_05921_, _05920_, _05915_);
  and (_05922_, _05907_, _05220_);
  and (_05923_, _05922_, \oc8051_golden_model_1.SCON [7]);
  and (_05924_, _05907_, _05228_);
  and (_05925_, _05924_, \oc8051_golden_model_1.IE [7]);
  nor (_05926_, _05925_, _05923_);
  and (_05927_, _05907_, _05208_);
  and (_05928_, _05927_, \oc8051_golden_model_1.TCON [7]);
  and (_05929_, _05238_, _05900_);
  and (_05930_, _05929_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05931_, _05930_, _05928_);
  and (_05932_, _05931_, _05926_);
  and (_05933_, _05932_, _05921_);
  and (_05934_, _05933_, _05913_);
  and (_05935_, _05934_, _05205_);
  nor (_05936_, _05935_, _05211_);
  and (_05937_, _05211_, \oc8051_golden_model_1.PSW [7]);
  nor (_05938_, _05937_, _05936_);
  nor (_05939_, _05938_, _05063_);
  not (_05940_, _04449_);
  and (_05941_, _05918_, \oc8051_golden_model_1.P2 [7]);
  and (_05942_, _05929_, \oc8051_golden_model_1.P3 [7]);
  or (_05943_, _05942_, _05941_);
  nor (_05944_, _05943_, _05928_);
  and (_05945_, _05209_, \oc8051_golden_model_1.P0 [7]);
  and (_05946_, _05916_, \oc8051_golden_model_1.P1 [7]);
  nor (_05947_, _05946_, _05945_);
  and (_05948_, _05947_, _05926_);
  and (_05949_, _05948_, _05913_);
  and (_05950_, _05949_, _05944_);
  and (_05951_, _05950_, _05205_);
  nor (_05952_, _05951_, _05211_);
  or (_05953_, _05952_, _05940_);
  not (_05954_, _04428_);
  and (_05955_, _05824_, _05517_);
  not (_05956_, _05666_);
  and (_05957_, _05956_, _05617_);
  and (_05958_, _05717_, _05566_);
  and (_05959_, _05958_, _05957_);
  and (_05960_, _05959_, _05955_);
  and (_05961_, _05960_, _05411_);
  nor (_05962_, _05961_, _05310_);
  and (_05963_, _05961_, _05310_);
  nor (_05964_, _05963_, _05962_);
  and (_05965_, _05964_, _04421_);
  not (_05966_, _04422_);
  nor (_05967_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_05968_, _05967_, _03995_);
  nor (_05969_, _05968_, _03722_);
  nor (_05970_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_05971_, _05970_, _03722_);
  and (_05972_, _05971_, _03498_);
  nor (_05973_, _05972_, _05969_);
  nor (_05974_, _05973_, _03997_);
  not (_05975_, _05974_);
  not (_05976_, _04463_);
  nand (_05977_, _05005_, _05976_);
  and (_05978_, _04463_, _03581_);
  not (_05979_, _05978_);
  and (_05980_, _05979_, _03997_);
  nand (_05981_, _05980_, _05977_);
  and (_05982_, _05981_, _05975_);
  nor (_05983_, _05967_, _03995_);
  nor (_05984_, _05983_, _05968_);
  nor (_05985_, _05984_, _03997_);
  not (_05986_, _05985_);
  nand (_05987_, _04875_, _05976_);
  and (_05988_, _04463_, _03904_);
  not (_05989_, _05988_);
  and (_05990_, _05989_, _03997_);
  nand (_05991_, _05990_, _05987_);
  and (_05992_, _05991_, _05986_);
  or (_05993_, _04463_, _04620_);
  not (_05994_, _03997_);
  and (_05995_, _04463_, _04048_);
  nor (_05997_, _05995_, _05994_);
  nand (_05998_, _05997_, _05993_);
  nor (_06000_, _03997_, \oc8051_golden_model_1.SP [0]);
  not (_06001_, _06000_);
  nand (_06003_, _06001_, _05998_);
  or (_06004_, _06003_, _05144_);
  nor (_06006_, _03500_, _03997_);
  not (_06007_, _06006_);
  or (_06009_, _04406_, _04463_);
  or (_06010_, _05976_, _03414_);
  and (_06012_, _06010_, _03997_);
  nand (_06013_, _06012_, _06009_);
  and (_06015_, _06013_, _06007_);
  not (_06016_, _06015_);
  and (_06018_, _06001_, _05998_);
  or (_06019_, _06018_, _05146_);
  and (_06021_, _06019_, _06016_);
  nand (_06022_, _06021_, _06004_);
  or (_06024_, _06003_, _05152_);
  or (_06025_, _06018_, _05150_);
  and (_06027_, _06025_, _06015_);
  nand (_06028_, _06027_, _06024_);
  nand (_06030_, _06028_, _06022_);
  nand (_06031_, _06030_, _05992_);
  not (_06033_, _05992_);
  or (_06034_, _06003_, _05164_);
  or (_06035_, _06018_, _05166_);
  and (_06036_, _06035_, _06016_);
  nand (_06037_, _06036_, _06034_);
  or (_06038_, _06003_, _05160_);
  or (_06039_, _06018_, _05158_);
  and (_06040_, _06039_, _06015_);
  nand (_06041_, _06040_, _06038_);
  nand (_06042_, _06041_, _06037_);
  nand (_06043_, _06042_, _06033_);
  nand (_06044_, _06043_, _06031_);
  nand (_06045_, _06044_, _05982_);
  not (_06046_, _05982_);
  or (_06047_, _06003_, _05176_);
  or (_06048_, _06018_, _05174_);
  and (_06049_, _06048_, _06015_);
  nand (_06050_, _06049_, _06047_);
  or (_06051_, _06003_, _05180_);
  or (_06052_, _06018_, _05182_);
  and (_06053_, _06052_, _06016_);
  nand (_06054_, _06053_, _06051_);
  nand (_06055_, _06054_, _06050_);
  nand (_06056_, _06055_, _05992_);
  or (_06057_, _06003_, _05194_);
  or (_06058_, _06018_, _05196_);
  and (_06059_, _06058_, _06016_);
  nand (_06060_, _06059_, _06057_);
  or (_06061_, _06003_, _05190_);
  or (_06062_, _06018_, _05188_);
  and (_06063_, _06062_, _06015_);
  nand (_06064_, _06063_, _06061_);
  nand (_06065_, _06064_, _06060_);
  nand (_06066_, _06065_, _06033_);
  nand (_06067_, _06066_, _06056_);
  nand (_06068_, _06067_, _06046_);
  and (_06069_, _06068_, _06045_);
  or (_06070_, _06069_, _05966_);
  not (_06071_, _04421_);
  or (_06072_, _03229_, _03219_);
  not (_06073_, _06072_);
  and (_06074_, _06073_, _05842_);
  not (_06075_, \oc8051_golden_model_1.ACC [7]);
  nor (_06076_, _03980_, _06075_);
  and (_06077_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_06078_, _06077_, \oc8051_golden_model_1.PC [6]);
  and (_06079_, _06078_, _03295_);
  and (_06080_, _06079_, \oc8051_golden_model_1.PC [7]);
  nor (_06081_, _06079_, \oc8051_golden_model_1.PC [7]);
  nor (_06082_, _06081_, _06080_);
  and (_06083_, _06082_, _03980_);
  or (_06084_, _06083_, _06076_);
  and (_06085_, _06084_, _06072_);
  or (_06086_, _06085_, _04422_);
  or (_06087_, _06086_, _06074_);
  and (_06088_, _06087_, _06071_);
  and (_06089_, _06088_, _06070_);
  or (_06090_, _06089_, _05965_);
  and (_06092_, _06090_, _05954_);
  not (_06094_, _05211_);
  nand (_06095_, _05951_, _06094_);
  and (_06097_, _06095_, _04428_);
  or (_06098_, _06097_, _04768_);
  or (_06100_, _06098_, _06092_);
  nor (_06101_, _06082_, _03230_);
  nor (_06103_, _06101_, _04431_);
  and (_06104_, _06103_, _06100_);
  and (_06106_, _05833_, _04431_);
  or (_06107_, _06106_, _04449_);
  or (_06109_, _06107_, _06104_);
  and (_06110_, _06109_, _05953_);
  or (_06112_, _06110_, _03508_);
  not (_06113_, _05259_);
  nor (_06115_, _05272_, _05264_);
  and (_06116_, _06115_, _05288_);
  and (_06118_, _06116_, _06113_);
  and (_06119_, _06118_, _05306_);
  and (_06121_, _05280_, _05232_);
  and (_06122_, _05235_, \oc8051_golden_model_1.P2INREG [7]);
  and (_06124_, _05239_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06125_, _06124_, _06122_);
  and (_06126_, _05266_, \oc8051_golden_model_1.P1INREG [7]);
  and (_06127_, _05293_, \oc8051_golden_model_1.P0INREG [7]);
  nor (_06128_, _06127_, _06126_);
  and (_06129_, _06128_, _06125_);
  and (_06130_, _06129_, _05257_);
  and (_06131_, _06130_, _06121_);
  and (_06132_, _06131_, _06119_);
  and (_06133_, _06132_, _05205_);
  nand (_06134_, _06133_, _03508_);
  and (_06135_, _06134_, _04562_);
  and (_06136_, _06135_, _06112_);
  nor (_06137_, _05951_, _06094_);
  not (_06138_, _06137_);
  and (_06139_, _06138_, _06095_);
  and (_06140_, _06139_, _04454_);
  or (_06141_, _06140_, _06136_);
  and (_06142_, _06141_, _03227_);
  not (_06143_, _06082_);
  nor (_06144_, _06143_, _03227_);
  or (_06145_, _06144_, _03745_);
  or (_06146_, _06145_, _06142_);
  nand (_06147_, _06133_, _03745_);
  and (_06148_, _06147_, _06146_);
  or (_06149_, _06148_, _04463_);
  and (_06150_, _06069_, _03446_);
  nand (_06151_, _06132_, _04463_);
  or (_06152_, _06151_, _06150_);
  and (_06153_, _06152_, _05063_);
  and (_06154_, _06153_, _06149_);
  or (_06155_, _06154_, _05939_);
  and (_06156_, _06155_, _05897_);
  nand (_06157_, _06082_, _03224_);
  nand (_06158_, _06157_, _04480_);
  or (_06159_, _06158_, _06156_);
  or (_06160_, _05833_, _04480_);
  and (_06161_, _06160_, _06159_);
  or (_06162_, _06161_, _04482_);
  not (_06163_, _04483_);
  not (_06164_, _04482_);
  or (_06165_, _06069_, _06164_);
  and (_06166_, _06165_, _06163_);
  and (_06167_, _06166_, _06162_);
  not (_06168_, _05894_);
  and (_06169_, _03446_, _03222_);
  not (_06170_, _06169_);
  not (_06171_, _05881_);
  nor (_06172_, _06171_, _05204_);
  and (_06173_, _03946_, _03708_);
  and (_06174_, _03654_, _02224_);
  and (_06175_, _03657_, _02202_);
  nor (_06176_, _06175_, _06174_);
  and (_06177_, _03687_, _02221_);
  and (_06178_, _03698_, _02196_);
  nor (_06179_, _06178_, _06177_);
  and (_06180_, _06179_, _06176_);
  and (_06181_, _03701_, _02187_);
  and (_06182_, _03703_, _02190_);
  nor (_06183_, _06182_, _06181_);
  and (_06184_, _03675_, _02213_);
  and (_06185_, _03678_, _02217_);
  nor (_06186_, _06185_, _06184_);
  and (_06187_, _06186_, _06183_);
  and (_06188_, _06187_, _06180_);
  and (_06189_, _03690_, _02233_);
  and (_06190_, _03692_, _02228_);
  nor (_06191_, _06190_, _06189_);
  and (_06192_, _03685_, _02226_);
  and (_06193_, _03662_, _02235_);
  nor (_06194_, _06193_, _06192_);
  and (_06195_, _06194_, _06191_);
  and (_06196_, _03672_, _02210_);
  and (_06197_, _03680_, _02185_);
  nor (_06198_, _06197_, _06196_);
  and (_06199_, _03696_, _02193_);
  and (_06200_, _03665_, _02200_);
  nor (_06201_, _06200_, _06199_);
  and (_06202_, _06201_, _06198_);
  and (_06203_, _06202_, _06195_);
  and (_06204_, _06203_, _06188_);
  and (_06205_, _06204_, _06171_);
  and (_06206_, _03685_, _02114_);
  and (_06207_, _03703_, _02080_);
  nor (_06208_, _06207_, _06206_);
  and (_06209_, _03692_, _02117_);
  and (_06210_, _03680_, _02075_);
  nor (_06211_, _06210_, _06209_);
  and (_06212_, _06211_, _06208_);
  and (_06213_, _03665_, _02090_);
  and (_06214_, _03701_, _02077_);
  nor (_06215_, _06214_, _06213_);
  and (_06216_, _03654_, _02087_);
  and (_06217_, _03678_, _02125_);
  nor (_06218_, _06217_, _06216_);
  and (_06219_, _06218_, _06215_);
  and (_06220_, _06219_, _06212_);
  and (_06221_, _03675_, _02101_);
  and (_06222_, _03657_, _02112_);
  nor (_06223_, _06222_, _06221_);
  and (_06224_, _03687_, _02098_);
  and (_06225_, _03696_, _02084_);
  nor (_06226_, _06225_, _06224_);
  and (_06227_, _06226_, _06223_);
  and (_06228_, _03690_, _02104_);
  and (_06229_, _03698_, _02082_);
  nor (_06230_, _06229_, _06228_);
  and (_06231_, _03662_, _02109_);
  and (_06232_, _03672_, _02123_);
  nor (_06233_, _06232_, _06231_);
  and (_06234_, _06233_, _06230_);
  and (_06235_, _06234_, _06227_);
  and (_06236_, _06235_, _06220_);
  and (_06237_, _03685_, _02170_);
  and (_06238_, _03657_, _02139_);
  nor (_06239_, _06238_, _06237_);
  and (_06240_, _03687_, _02154_);
  and (_06241_, _03698_, _02144_);
  nor (_06242_, _06241_, _06240_);
  and (_06243_, _06242_, _06239_);
  and (_06244_, _03675_, _02178_);
  and (_06245_, _03672_, _02160_);
  nor (_06246_, _06245_, _06244_);
  and (_06247_, _03692_, _02173_);
  and (_06248_, _03654_, _02146_);
  nor (_06249_, _06248_, _06247_);
  and (_06250_, _06249_, _06246_);
  and (_06251_, _06250_, _06243_);
  and (_06252_, _03690_, _02165_);
  and (_06253_, _03662_, _02157_);
  nor (_06254_, _06253_, _06252_);
  and (_06255_, _03665_, _02168_);
  and (_06256_, _03701_, _02132_);
  nor (_06257_, _06256_, _06255_);
  and (_06258_, _06257_, _06254_);
  and (_06259_, _03696_, _02137_);
  and (_06260_, _03678_, _02180_);
  nor (_06261_, _06260_, _06259_);
  and (_06262_, _03680_, _02135_);
  and (_06263_, _03703_, _02130_);
  nor (_06264_, _06263_, _06262_);
  and (_06265_, _06264_, _06261_);
  and (_06266_, _06265_, _06258_);
  and (_06267_, _06266_, _06251_);
  and (_06268_, _06267_, _06236_);
  and (_06269_, _06268_, _06205_);
  nor (_06270_, _04303_, _04163_);
  and (_06271_, _06270_, _06269_);
  and (_06272_, _06271_, _06173_);
  and (_06273_, _06272_, \oc8051_golden_model_1.DPH [7]);
  not (_06274_, _04163_);
  and (_06275_, _04303_, _06274_);
  not (_06276_, _03708_);
  and (_06277_, _03946_, _06276_);
  and (_06278_, _06277_, _06269_);
  and (_06279_, _06278_, _06275_);
  and (_06280_, _06279_, \oc8051_golden_model_1.TMOD [7]);
  nor (_06281_, _06280_, _06273_);
  not (_06282_, _04303_);
  and (_06283_, _06282_, _04163_);
  and (_06284_, _06283_, _06278_);
  and (_06285_, _06284_, \oc8051_golden_model_1.TL0 [7]);
  nor (_06286_, _03946_, _03708_);
  and (_06287_, _06286_, _06269_);
  and (_06288_, _06287_, _06275_);
  and (_06289_, _06288_, \oc8051_golden_model_1.TH1 [7]);
  nor (_06290_, _06289_, _06285_);
  and (_06291_, _06290_, _06281_);
  and (_06292_, _04303_, _04163_);
  and (_06293_, _06292_, _06277_);
  nor (_06294_, _06267_, _06236_);
  and (_06295_, _06294_, _06205_);
  and (_06296_, _06295_, _06293_);
  and (_06297_, _06296_, \oc8051_golden_model_1.IP [7]);
  not (_06298_, _06236_);
  and (_06299_, _06267_, _06298_);
  and (_06300_, _06292_, _06173_);
  nor (_06301_, _06204_, _05881_);
  and (_06302_, _06301_, _06300_);
  and (_06303_, _06302_, _06299_);
  and (_06304_, _06303_, \oc8051_golden_model_1.PSW [7]);
  nor (_06305_, _06304_, _06297_);
  not (_06306_, _06267_);
  and (_06307_, _06306_, _06236_);
  and (_06308_, _06307_, _06302_);
  and (_06309_, _06308_, \oc8051_golden_model_1.ACC [7]);
  and (_06310_, _06302_, _06294_);
  and (_06311_, _06310_, \oc8051_golden_model_1.B [7]);
  nor (_06312_, _06311_, _06309_);
  and (_06313_, _06312_, _06305_);
  and (_06314_, _06307_, _06205_);
  and (_06315_, _06314_, _06293_);
  and (_06316_, _06315_, \oc8051_golden_model_1.IE [7]);
  and (_06317_, _06299_, _06205_);
  and (_06318_, _06277_, _06275_);
  and (_06319_, _06318_, _06317_);
  and (_06320_, _06319_, \oc8051_golden_model_1.SBUF [7]);
  and (_06321_, _06317_, _06293_);
  and (_06322_, _06321_, \oc8051_golden_model_1.SCON [7]);
  or (_06323_, _06322_, _06320_);
  nor (_06324_, _06323_, _06316_);
  and (_06325_, _06324_, _06313_);
  and (_06326_, _06325_, _06291_);
  and (_06327_, _06292_, _06287_);
  and (_06328_, _06327_, \oc8051_golden_model_1.TH0 [7]);
  and (_06329_, _06277_, _06271_);
  and (_06330_, _06329_, \oc8051_golden_model_1.TL1 [7]);
  nor (_06331_, _06330_, _06328_);
  not (_06332_, _03946_);
  and (_06333_, _06332_, _03708_);
  and (_06334_, _06333_, _06271_);
  and (_06335_, _06334_, \oc8051_golden_model_1.PCON [7]);
  and (_06336_, _06292_, _06278_);
  and (_06337_, _06336_, \oc8051_golden_model_1.TCON [7]);
  nor (_06338_, _06337_, _06335_);
  and (_06339_, _06338_, _06331_);
  and (_06340_, _06317_, _06300_);
  and (_06341_, _06340_, \oc8051_golden_model_1.P1INREG [7]);
  not (_06342_, _06341_);
  and (_06343_, _06300_, _06269_);
  and (_06344_, _06343_, \oc8051_golden_model_1.P0INREG [7]);
  not (_06345_, _06344_);
  and (_06346_, _06314_, _06300_);
  and (_06347_, _06346_, \oc8051_golden_model_1.P2INREG [7]);
  and (_06348_, _06300_, _06295_);
  and (_06349_, _06348_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06350_, _06349_, _06347_);
  and (_06351_, _06350_, _06345_);
  and (_06352_, _06351_, _06342_);
  and (_06353_, _06269_, _06173_);
  and (_06354_, _06353_, _06275_);
  and (_06355_, _06354_, \oc8051_golden_model_1.SP [7]);
  and (_06356_, _06353_, _06283_);
  and (_06357_, _06356_, \oc8051_golden_model_1.DPL [7]);
  nor (_06358_, _06357_, _06355_);
  and (_06359_, _06358_, _06352_);
  and (_06360_, _06359_, _06339_);
  and (_06361_, _06360_, _06326_);
  not (_06362_, _06361_);
  nor (_06363_, _06362_, _06172_);
  nor (_06364_, _06363_, _06170_);
  or (_06365_, _06364_, _06168_);
  or (_06366_, _06365_, _06167_);
  and (_06367_, _06366_, _05896_);
  and (_06368_, _06171_, _04500_);
  or (_06369_, _06368_, _03178_);
  or (_06370_, _06369_, _06367_);
  and (_06371_, _06143_, _03178_);
  nor (_06372_, _06371_, _04512_);
  and (_06373_, _06372_, _06370_);
  or (_06374_, _06373_, _05885_);
  and (_06375_, _06374_, _05850_);
  nor (_06376_, _05309_, _06075_);
  and (_06377_, _05309_, _06075_);
  nor (_06378_, _06377_, _06376_);
  and (_06379_, _06378_, _04511_);
  or (_06380_, _06379_, _04515_);
  or (_06381_, _06380_, _06375_);
  not (_06382_, _04514_);
  not (_06383_, _04515_);
  or (_06384_, _05883_, _06383_);
  and (_06385_, _06384_, _06382_);
  and (_06386_, _06385_, _06381_);
  and (_06387_, _06376_, _04514_);
  or (_06388_, _06387_, _03192_);
  or (_06389_, _06388_, _06386_);
  and (_06390_, _03624_, _03446_);
  and (_06391_, _06143_, _03192_);
  nor (_06392_, _06391_, _06390_);
  and (_06393_, _06392_, _06389_);
  and (_06394_, _03785_, _03446_);
  not (_06395_, _06390_);
  nor (_06396_, _05882_, _06395_);
  or (_06397_, _06396_, _06394_);
  or (_06398_, _06397_, _06393_);
  not (_06399_, _03188_);
  nand (_06400_, _06377_, _06394_);
  and (_06401_, _06400_, _06399_);
  and (_06402_, _06401_, _06398_);
  nand (_06403_, _06082_, _03188_);
  nand (_06404_, _06403_, _05848_);
  or (_06405_, _06404_, _06402_);
  and (_06406_, _06405_, _05849_);
  or (_06407_, _06406_, _04533_);
  not (_06408_, _04531_);
  not (_06409_, _04533_);
  not (_06410_, _06069_);
  or (_06411_, _06003_, _05311_);
  or (_06412_, _06018_, _05313_);
  and (_06413_, _06412_, _06016_);
  nand (_06414_, _06413_, _06411_);
  or (_06415_, _06003_, _05319_);
  or (_06416_, _06018_, _05317_);
  and (_06417_, _06416_, _06015_);
  nand (_06418_, _06417_, _06415_);
  nand (_06419_, _06418_, _06414_);
  nand (_06420_, _06419_, _05992_);
  or (_06421_, _06003_, _05331_);
  or (_06422_, _06018_, _05333_);
  and (_06423_, _06422_, _06016_);
  nand (_06424_, _06423_, _06421_);
  or (_06425_, _06003_, _05327_);
  or (_06426_, _06018_, _05325_);
  and (_06427_, _06426_, _06015_);
  nand (_06428_, _06427_, _06425_);
  nand (_06429_, _06428_, _06424_);
  nand (_06430_, _06429_, _06033_);
  and (_06431_, _06430_, _05982_);
  and (_06432_, _06431_, _06420_);
  or (_06433_, _06003_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_06434_, _06018_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_06435_, _06434_, _06433_);
  nand (_06436_, _06435_, _06015_);
  or (_06437_, _06003_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_06438_, _06018_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_06439_, _06438_, _06437_);
  nand (_06440_, _06439_, _06016_);
  nand (_06441_, _06440_, _06436_);
  nand (_06442_, _06441_, _05992_);
  or (_06443_, _06003_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_06444_, _06018_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_06445_, _06444_, _06443_);
  nand (_06446_, _06445_, _06015_);
  or (_06447_, _06003_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_06448_, _06018_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_06449_, _06448_, _06447_);
  nand (_06450_, _06449_, _06016_);
  nand (_06451_, _06450_, _06446_);
  nand (_06452_, _06451_, _06033_);
  and (_06453_, _06452_, _06046_);
  and (_06454_, _06453_, _06442_);
  or (_06455_, _06454_, _06432_);
  not (_06456_, _06455_);
  or (_06457_, _06003_, _04017_);
  or (_06458_, _06018_, _04347_);
  and (_06459_, _06458_, _06016_);
  nand (_06460_, _06459_, _06457_);
  or (_06461_, _06003_, _04355_);
  or (_06462_, _06018_, _04352_);
  and (_06463_, _06462_, _06015_);
  nand (_06464_, _06463_, _06461_);
  nand (_06465_, _06464_, _06460_);
  nand (_06466_, _06465_, _05992_);
  or (_06467_, _06003_, _04368_);
  or (_06468_, _06018_, _04370_);
  and (_06469_, _06468_, _06016_);
  nand (_06470_, _06469_, _06467_);
  or (_06471_, _06003_, _04364_);
  or (_06472_, _06018_, _04362_);
  and (_06473_, _06472_, _06015_);
  nand (_06474_, _06473_, _06471_);
  nand (_06475_, _06474_, _06470_);
  nand (_06476_, _06475_, _06033_);
  and (_06477_, _06476_, _05982_);
  and (_06478_, _06477_, _06466_);
  or (_06479_, _06003_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_06480_, _06018_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_06481_, _06480_, _06479_);
  nand (_06482_, _06481_, _06015_);
  or (_06483_, _06003_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_06484_, _06018_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_06485_, _06484_, _06483_);
  nand (_06486_, _06485_, _06016_);
  nand (_06487_, _06486_, _06482_);
  nand (_06488_, _06487_, _05992_);
  or (_06489_, _06003_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_06490_, _06018_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_06491_, _06490_, _06489_);
  nand (_06492_, _06491_, _06015_);
  or (_06493_, _06003_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_06494_, _06018_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_06495_, _06494_, _06493_);
  nand (_06496_, _06495_, _06016_);
  nand (_06497_, _06496_, _06492_);
  nand (_06498_, _06497_, _06033_);
  and (_06499_, _06498_, _06046_);
  and (_06500_, _06499_, _06488_);
  or (_06501_, _06500_, _06478_);
  or (_06502_, _06003_, _04563_);
  or (_06503_, _06018_, _04565_);
  and (_06504_, _06503_, _06016_);
  nand (_06505_, _06504_, _06502_);
  or (_06506_, _06003_, _04571_);
  or (_06507_, _06018_, _04569_);
  and (_06508_, _06507_, _06015_);
  nand (_06509_, _06508_, _06506_);
  nand (_06510_, _06509_, _06505_);
  nand (_06511_, _06510_, _05992_);
  or (_06512_, _06003_, _04584_);
  or (_06513_, _06018_, _04586_);
  and (_06514_, _06513_, _06016_);
  nand (_06515_, _06514_, _06512_);
  or (_06516_, _06003_, _04580_);
  or (_06517_, _06018_, _04578_);
  and (_06518_, _06517_, _06015_);
  nand (_06519_, _06518_, _06516_);
  nand (_06520_, _06519_, _06515_);
  nand (_06521_, _06520_, _06033_);
  and (_06522_, _06521_, _05982_);
  and (_06523_, _06522_, _06511_);
  or (_06524_, _06003_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_06525_, _06018_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_06526_, _06525_, _06524_);
  nand (_06527_, _06526_, _06015_);
  or (_06528_, _06003_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_06529_, _06018_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_06530_, _06529_, _06528_);
  nand (_06531_, _06530_, _06016_);
  nand (_06532_, _06531_, _06527_);
  nand (_06533_, _06532_, _05992_);
  or (_06534_, _06003_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_06535_, _06018_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_06536_, _06535_, _06534_);
  nand (_06537_, _06536_, _06015_);
  or (_06538_, _06003_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_06539_, _06018_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_06540_, _06539_, _06538_);
  nand (_06541_, _06540_, _06016_);
  nand (_06542_, _06541_, _06537_);
  nand (_06543_, _06542_, _06033_);
  and (_06544_, _06543_, _06046_);
  and (_06545_, _06544_, _06533_);
  or (_06546_, _06545_, _06523_);
  nor (_06547_, _06546_, _06501_);
  or (_06548_, _06003_, _04953_);
  or (_06549_, _06018_, _04955_);
  and (_06550_, _06549_, _06016_);
  nand (_06551_, _06550_, _06548_);
  or (_06552_, _06003_, _04961_);
  or (_06553_, _06018_, _04959_);
  and (_06554_, _06553_, _06015_);
  nand (_06555_, _06554_, _06552_);
  nand (_06556_, _06555_, _06551_);
  nand (_06557_, _06556_, _05992_);
  or (_06558_, _06003_, _04973_);
  or (_06559_, _06018_, _04975_);
  and (_06560_, _06559_, _06016_);
  nand (_06561_, _06560_, _06558_);
  or (_06562_, _06003_, _04969_);
  or (_06563_, _06018_, _04967_);
  and (_06564_, _06563_, _06015_);
  nand (_06565_, _06564_, _06562_);
  nand (_06566_, _06565_, _06561_);
  nand (_06567_, _06566_, _06033_);
  and (_06568_, _06567_, _05982_);
  and (_06569_, _06568_, _06557_);
  or (_06570_, _06003_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_06571_, _06018_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_06572_, _06571_, _06570_);
  nand (_06573_, _06572_, _06015_);
  or (_06574_, _06003_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_06575_, _06018_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_06576_, _06575_, _06574_);
  nand (_06577_, _06576_, _06016_);
  nand (_06578_, _06577_, _06573_);
  nand (_06579_, _06578_, _05992_);
  or (_06580_, _06003_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_06581_, _06018_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_06582_, _06581_, _06580_);
  nand (_06583_, _06582_, _06015_);
  or (_06584_, _06003_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_06585_, _06018_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_06586_, _06585_, _06584_);
  nand (_06587_, _06586_, _06016_);
  nand (_06588_, _06587_, _06583_);
  nand (_06589_, _06588_, _06033_);
  and (_06590_, _06589_, _06046_);
  and (_06591_, _06590_, _06579_);
  or (_06592_, _06591_, _06569_);
  or (_06593_, _06003_, _04819_);
  or (_06594_, _06018_, _04821_);
  and (_06595_, _06594_, _06016_);
  nand (_06596_, _06595_, _06593_);
  or (_06597_, _06003_, _04827_);
  or (_06598_, _06018_, _04825_);
  and (_06599_, _06598_, _06015_);
  nand (_06600_, _06599_, _06597_);
  nand (_06601_, _06600_, _06596_);
  nand (_06602_, _06601_, _05992_);
  or (_06603_, _06003_, _04839_);
  or (_06604_, _06018_, _04841_);
  and (_06605_, _06604_, _06016_);
  nand (_06606_, _06605_, _06603_);
  or (_06607_, _06003_, _04835_);
  or (_06608_, _06018_, _04833_);
  and (_06609_, _06608_, _06015_);
  nand (_06610_, _06609_, _06607_);
  nand (_06611_, _06610_, _06606_);
  nand (_06612_, _06611_, _06033_);
  and (_06613_, _06612_, _05982_);
  and (_06614_, _06613_, _06602_);
  or (_06615_, _06003_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_06616_, _06018_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_06617_, _06616_, _06615_);
  nand (_06618_, _06617_, _06015_);
  or (_06619_, _06003_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_06620_, _06018_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_06621_, _06620_, _06619_);
  nand (_06622_, _06621_, _06016_);
  nand (_06623_, _06622_, _06618_);
  nand (_06624_, _06623_, _05992_);
  or (_06625_, _06003_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_06626_, _06018_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_06627_, _06626_, _06625_);
  nand (_06628_, _06627_, _06015_);
  or (_06629_, _06003_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_06630_, _06018_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_06631_, _06630_, _06629_);
  nand (_06632_, _06631_, _06016_);
  nand (_06633_, _06632_, _06628_);
  nand (_06634_, _06633_, _06033_);
  and (_06635_, _06634_, _06046_);
  and (_06636_, _06635_, _06624_);
  or (_06637_, _06636_, _06614_);
  nor (_06638_, _06637_, _06592_);
  and (_06639_, _06638_, _06547_);
  or (_06640_, _06003_, _05413_);
  or (_06641_, _06018_, _05415_);
  and (_06642_, _06641_, _06016_);
  nand (_06643_, _06642_, _06640_);
  or (_06644_, _06003_, _05421_);
  or (_06645_, _06018_, _05419_);
  and (_06646_, _06645_, _06015_);
  nand (_06647_, _06646_, _06644_);
  nand (_06648_, _06647_, _06643_);
  nand (_06649_, _06648_, _05992_);
  or (_06650_, _06003_, _05433_);
  or (_06651_, _06018_, _05435_);
  and (_06652_, _06651_, _06016_);
  nand (_06653_, _06652_, _06650_);
  or (_06654_, _06003_, _05429_);
  or (_06655_, _06018_, _05427_);
  and (_06656_, _06655_, _06015_);
  nand (_06657_, _06656_, _06654_);
  nand (_06658_, _06657_, _06653_);
  nand (_06659_, _06658_, _06033_);
  and (_06660_, _06659_, _05982_);
  and (_06661_, _06660_, _06649_);
  or (_06662_, _06003_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_06663_, _06018_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_06664_, _06663_, _06662_);
  nand (_06665_, _06664_, _06015_);
  or (_06666_, _06003_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_06667_, _06018_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_06668_, _06667_, _06666_);
  nand (_06669_, _06668_, _06016_);
  nand (_06670_, _06669_, _06665_);
  nand (_06671_, _06670_, _05992_);
  or (_06672_, _06003_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_06673_, _06018_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_06674_, _06673_, _06672_);
  nand (_06675_, _06674_, _06015_);
  or (_06676_, _06003_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_06677_, _06018_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_06678_, _06677_, _06676_);
  nand (_06679_, _06678_, _06016_);
  nand (_06680_, _06679_, _06675_);
  nand (_06681_, _06680_, _06033_);
  and (_06682_, _06681_, _06046_);
  and (_06683_, _06682_, _06671_);
  or (_06684_, _06683_, _06661_);
  or (_06685_, _06003_, _05721_);
  or (_06686_, _06018_, _05723_);
  and (_06687_, _06686_, _06016_);
  nand (_06688_, _06687_, _06685_);
  or (_06689_, _06003_, _05729_);
  or (_06690_, _06018_, _05727_);
  and (_06691_, _06690_, _06015_);
  nand (_06692_, _06691_, _06689_);
  nand (_06693_, _06692_, _06688_);
  nand (_06694_, _06693_, _05992_);
  or (_06696_, _06003_, _05741_);
  or (_06697_, _06018_, _05743_);
  and (_06698_, _06697_, _06016_);
  nand (_06699_, _06698_, _06696_);
  or (_06700_, _06003_, _05737_);
  or (_06701_, _06018_, _05735_);
  and (_06702_, _06701_, _06015_);
  nand (_06703_, _06702_, _06700_);
  nand (_06704_, _06703_, _06699_);
  nand (_06705_, _06704_, _06033_);
  and (_06706_, _06705_, _05982_);
  and (_06707_, _06706_, _06694_);
  or (_06708_, _06003_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_06709_, _06018_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_06710_, _06709_, _06708_);
  nand (_06711_, _06710_, _06015_);
  or (_06712_, _06003_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_06713_, _06018_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_06714_, _06713_, _06712_);
  nand (_06715_, _06714_, _06016_);
  nand (_06716_, _06715_, _06711_);
  nand (_06717_, _06716_, _05992_);
  or (_06718_, _06003_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_06719_, _06018_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_06720_, _06719_, _06718_);
  nand (_06721_, _06720_, _06015_);
  or (_06722_, _06003_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_06723_, _06018_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_06724_, _06723_, _06722_);
  nand (_06725_, _06724_, _06016_);
  nand (_06726_, _06725_, _06721_);
  nand (_06727_, _06726_, _06033_);
  and (_06728_, _06727_, _06046_);
  and (_06729_, _06728_, _06717_);
  or (_06730_, _06729_, _06707_);
  nor (_06731_, _06730_, _06684_);
  and (_06732_, _06731_, _06639_);
  and (_06733_, _06732_, _06456_);
  nor (_06734_, _06733_, _06410_);
  and (_06735_, _06733_, _06410_);
  or (_06736_, _06735_, _06734_);
  or (_06737_, _06736_, _06409_);
  and (_06738_, _06737_, _06408_);
  and (_06739_, _06738_, _06407_);
  and (_06740_, _05964_, _04531_);
  or (_06741_, _06740_, _03629_);
  or (_06742_, _06741_, _06739_);
  and (_06743_, _02909_, \oc8051_golden_model_1.PC [2]);
  and (_06744_, _06743_, \oc8051_golden_model_1.PC [3]);
  and (_06745_, _06744_, _06078_);
  and (_06746_, _06745_, \oc8051_golden_model_1.PC [7]);
  nor (_06747_, _06745_, \oc8051_golden_model_1.PC [7]);
  nor (_06748_, _06747_, _06746_);
  not (_06749_, _06748_);
  nand (_06750_, _06749_, _03629_);
  and (_06751_, _06750_, _06742_);
  or (_06752_, _06751_, _03198_);
  and (_06753_, _06143_, _03198_);
  nor (_06754_, _06753_, _04539_);
  and (_06755_, _06754_, _06752_);
  and (_06756_, _05936_, _04539_);
  nor (_06757_, _04320_, _03960_);
  not (_06758_, _06757_);
  nor (_06759_, _06758_, _06756_);
  not (_06760_, _06759_);
  nor (_06761_, _06760_, _06755_);
  not (_06762_, _05469_);
  not (_06763_, _05777_);
  and (_06764_, _04405_, _04378_);
  and (_06765_, _06764_, _04620_);
  nor (_06766_, _04875_, _05005_);
  and (_06767_, _06766_, _06765_);
  and (_06768_, _06767_, _06763_);
  and (_06769_, _06768_, _06762_);
  and (_06770_, _05363_, _05204_);
  nor (_06771_, _05363_, _05204_);
  nor (_06772_, _06771_, _06770_);
  and (_06773_, _06772_, _06769_);
  nor (_06774_, _06769_, _05204_);
  nor (_06775_, _06774_, _06773_);
  and (_06776_, _06775_, _06758_);
  nor (_06777_, _06776_, _04547_);
  not (_06778_, _06777_);
  nor (_06779_, _06778_, _06761_);
  not (_06780_, _04547_);
  nor (_06781_, _06775_, _06780_);
  nor (_06782_, _06781_, _04552_);
  not (_06783_, _06782_);
  nor (_06784_, _06783_, _06779_);
  not (_06785_, _04552_);
  and (_06786_, _06546_, _06501_);
  and (_06787_, _06637_, _06592_);
  and (_06788_, _06787_, _06786_);
  and (_06789_, _06730_, _06684_);
  and (_06790_, _06789_, _06788_);
  and (_06791_, _06790_, _06455_);
  nor (_06792_, _06791_, _06410_);
  and (_06793_, _06791_, _06410_);
  or (_06794_, _06793_, _06792_);
  nor (_06795_, _06794_, _06785_);
  nor (_06796_, _06795_, _03448_);
  not (_06797_, _06796_);
  nor (_06798_, _06797_, _06784_);
  nor (_06799_, _06798_, _05832_);
  nor (_06800_, _06799_, _04797_);
  or (_06801_, _06800_, _05143_);
  and (_06802_, _06801_, _05142_);
  not (_06803_, \oc8051_golden_model_1.PC [15]);
  and (_06804_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and (_06805_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_06806_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_06807_, _06806_, _06805_);
  and (_06808_, _06807_, _06080_);
  and (_06809_, _06808_, _06804_);
  and (_06810_, _06809_, \oc8051_golden_model_1.PC [14]);
  and (_06811_, _06810_, _06803_);
  nor (_06812_, _06810_, _06803_);
  or (_06813_, _06812_, _06811_);
  not (_06814_, _06813_);
  nor (_06815_, _06814_, _03629_);
  and (_06816_, _06807_, _06746_);
  and (_06817_, _06816_, _06804_);
  and (_06818_, _06817_, \oc8051_golden_model_1.PC [14]);
  and (_06819_, _06818_, _06803_);
  nor (_06820_, _06818_, _06803_);
  or (_06821_, _06820_, _06819_);
  and (_06822_, _06821_, _03629_);
  or (_06823_, _06822_, _06815_);
  and (_06824_, _06823_, _05137_);
  and (_06825_, _06824_, _05140_);
  or (_40565_, _06825_, _06802_);
  not (_06826_, \oc8051_golden_model_1.B [7]);
  nor (_06827_, _43000_, _06826_);
  not (_06828_, _03790_);
  nor (_06829_, _05248_, _06826_);
  not (_06830_, _05248_);
  nor (_06831_, _06830_, _05204_);
  or (_06832_, _06831_, _06829_);
  and (_06833_, _04058_, _03168_);
  not (_06834_, _06833_);
  and (_06835_, _04750_, _03168_);
  not (_06836_, _06835_);
  and (_06837_, _06836_, _04477_);
  and (_06838_, _06837_, _06834_);
  or (_06839_, _06838_, _06832_);
  not (_06840_, _03719_);
  nor (_06841_, _05910_, _06826_);
  and (_06842_, _05952_, _05910_);
  or (_06843_, _06842_, _06841_);
  and (_06844_, _06843_, _03714_);
  and (_06845_, _05964_, _05248_);
  or (_06846_, _06845_, _06829_);
  or (_06847_, _06846_, _04081_);
  and (_06848_, _05248_, \oc8051_golden_model_1.ACC [7]);
  or (_06849_, _06848_, _06829_);
  and (_06850_, _06849_, _04409_);
  nor (_06851_, _04409_, _06826_);
  or (_06852_, _06851_, _03610_);
  or (_06853_, _06852_, _06850_);
  and (_06854_, _06853_, _04055_);
  and (_06855_, _06854_, _06847_);
  and (_06856_, _06095_, _05910_);
  or (_06857_, _06856_, _06841_);
  and (_06858_, _06857_, _03715_);
  or (_06859_, _06858_, _03723_);
  or (_06860_, _06859_, _06855_);
  or (_06861_, _06832_, _03996_);
  and (_06862_, _06861_, _06860_);
  or (_06863_, _06862_, _03729_);
  or (_06864_, _06849_, _03737_);
  and (_06865_, _06864_, _03736_);
  and (_06866_, _06865_, _06863_);
  or (_06867_, _06866_, _06844_);
  and (_06868_, _06867_, _06840_);
  and (_06869_, _03603_, _03751_);
  or (_06870_, _06841_, _06138_);
  and (_06871_, _06870_, _03719_);
  and (_06872_, _06871_, _06857_);
  or (_06873_, _06872_, _06869_);
  or (_06874_, _06873_, _06868_);
  not (_06875_, _06869_);
  and (_06876_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_06877_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_06878_, _06877_, _06876_);
  and (_06879_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_06880_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_06881_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_06882_, _06881_, _06880_);
  nor (_06883_, _06882_, _06878_);
  and (_06884_, _06883_, _06879_);
  nor (_06885_, _06884_, _06878_);
  and (_06886_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_06887_, _06886_, _06881_);
  and (_06888_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_06889_, _06888_, _06876_);
  nor (_06890_, _06889_, _06887_);
  not (_06891_, _06890_);
  nor (_06892_, _06891_, _06885_);
  and (_06893_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_06894_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_06895_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_06896_, _06895_, _06894_);
  nor (_06897_, _06895_, _06894_);
  nor (_06898_, _06897_, _06896_);
  and (_06899_, _06898_, _06893_);
  nor (_06900_, _06898_, _06893_);
  nor (_06901_, _06900_, _06899_);
  and (_06902_, _06891_, _06885_);
  nor (_06903_, _06902_, _06892_);
  and (_06904_, _06903_, _06901_);
  nor (_06905_, _06904_, _06892_);
  not (_06906_, _06881_);
  and (_06907_, _06886_, _06906_);
  and (_06908_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_06909_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_06910_, _06909_, _06894_);
  and (_06911_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_06912_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_06913_, _06912_, _06911_);
  nor (_06914_, _06913_, _06910_);
  and (_06915_, _06914_, _06908_);
  nor (_06916_, _06914_, _06908_);
  nor (_06917_, _06916_, _06915_);
  and (_06918_, _06917_, _06907_);
  nor (_06919_, _06917_, _06907_);
  nor (_06920_, _06919_, _06918_);
  not (_06921_, _06920_);
  nor (_06922_, _06921_, _06905_);
  and (_06923_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_06924_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_06925_, _06924_, _06923_);
  nor (_06926_, _06899_, _06896_);
  and (_06927_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_06928_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_06929_, _06928_, _06927_);
  nor (_06930_, _06928_, _06927_);
  nor (_06931_, _06930_, _06929_);
  not (_06932_, _06931_);
  nor (_06933_, _06932_, _06926_);
  and (_06934_, _06932_, _06926_);
  nor (_06935_, _06934_, _06933_);
  and (_06936_, _06935_, _06925_);
  nor (_06937_, _06935_, _06925_);
  nor (_06938_, _06937_, _06936_);
  and (_06939_, _06921_, _06905_);
  nor (_06940_, _06939_, _06922_);
  and (_06941_, _06940_, _06938_);
  nor (_06942_, _06941_, _06922_);
  nor (_06943_, _06915_, _06910_);
  and (_06944_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_06945_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_06946_, _06945_, _06944_);
  nor (_06947_, _06945_, _06944_);
  nor (_06948_, _06947_, _06946_);
  not (_06949_, _06948_);
  nor (_06950_, _06949_, _06943_);
  and (_06951_, _06949_, _06943_);
  nor (_06952_, _06951_, _06950_);
  and (_06953_, _06952_, _06929_);
  nor (_06954_, _06952_, _06929_);
  nor (_06955_, _06954_, _06953_);
  nor (_06956_, _06918_, _06887_);
  and (_06957_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_06958_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_06959_, _06958_, _06909_);
  nor (_06960_, _06958_, _06909_);
  nor (_06961_, _06960_, _06959_);
  and (_06962_, _06961_, _06957_);
  nor (_06963_, _06961_, _06957_);
  nor (_06964_, _06963_, _06962_);
  not (_06965_, _06964_);
  nor (_06966_, _06965_, _06956_);
  and (_06967_, _06965_, _06956_);
  nor (_06968_, _06967_, _06966_);
  and (_06969_, _06968_, _06955_);
  nor (_06970_, _06968_, _06955_);
  nor (_06971_, _06970_, _06969_);
  not (_06972_, _06971_);
  nor (_06973_, _06972_, _06942_);
  nor (_06974_, _06936_, _06933_);
  not (_06975_, _06974_);
  and (_06976_, _06972_, _06942_);
  nor (_06977_, _06976_, _06973_);
  and (_06978_, _06977_, _06975_);
  nor (_06979_, _06978_, _06973_);
  nor (_06980_, _06953_, _06950_);
  not (_06981_, _06980_);
  nor (_06982_, _06969_, _06966_);
  not (_06983_, _06982_);
  and (_06984_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_06985_, _06984_, _06909_);
  and (_06986_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_06987_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_06988_, _06987_, _06986_);
  nor (_06989_, _06988_, _06985_);
  nor (_06990_, _06962_, _06959_);
  and (_06991_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_06992_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_06993_, _06992_, _06991_);
  nor (_06994_, _06992_, _06991_);
  nor (_06995_, _06994_, _06993_);
  not (_06996_, _06995_);
  nor (_06997_, _06996_, _06990_);
  and (_06998_, _06996_, _06990_);
  nor (_06999_, _06998_, _06997_);
  and (_07000_, _06999_, _06946_);
  nor (_07001_, _06999_, _06946_);
  nor (_07002_, _07001_, _07000_);
  and (_07003_, _07002_, _06989_);
  nor (_07004_, _07002_, _06989_);
  nor (_07005_, _07004_, _07003_);
  and (_07006_, _07005_, _06983_);
  nor (_07007_, _07005_, _06983_);
  nor (_07008_, _07007_, _07006_);
  and (_07009_, _07008_, _06981_);
  nor (_07010_, _07008_, _06981_);
  nor (_07011_, _07010_, _07009_);
  not (_07012_, _07011_);
  nor (_07013_, _07012_, _06979_);
  nor (_07014_, _07009_, _07006_);
  nor (_07015_, _07000_, _06997_);
  not (_07016_, _07015_);
  and (_07017_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_07018_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_07019_, _07018_, _07017_);
  nor (_07020_, _07018_, _07017_);
  nor (_07021_, _07020_, _07019_);
  and (_07022_, _07021_, _06985_);
  nor (_07023_, _07021_, _06985_);
  nor (_07024_, _07023_, _07022_);
  and (_07025_, _07024_, _06993_);
  nor (_07026_, _07024_, _06993_);
  nor (_07027_, _07026_, _07025_);
  and (_07028_, _07027_, _06984_);
  nor (_07029_, _07027_, _06984_);
  nor (_07030_, _07029_, _07028_);
  and (_07031_, _07030_, _07003_);
  nor (_07032_, _07030_, _07003_);
  nor (_07033_, _07032_, _07031_);
  and (_07034_, _07033_, _07016_);
  nor (_07035_, _07033_, _07016_);
  nor (_07036_, _07035_, _07034_);
  not (_07037_, _07036_);
  nor (_07038_, _07037_, _07014_);
  and (_07039_, _07037_, _07014_);
  nor (_07040_, _07039_, _07038_);
  and (_07041_, _07040_, _07013_);
  nor (_07042_, _07034_, _07031_);
  nor (_07043_, _07025_, _07022_);
  not (_07044_, _07043_);
  and (_07045_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_07046_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_07047_, _07046_, _07045_);
  nor (_07048_, _07046_, _07045_);
  nor (_07049_, _07048_, _07047_);
  and (_07050_, _07049_, _07019_);
  nor (_07051_, _07049_, _07019_);
  nor (_07052_, _07051_, _07050_);
  and (_07053_, _07052_, _07028_);
  nor (_07054_, _07052_, _07028_);
  nor (_07055_, _07054_, _07053_);
  and (_07056_, _07055_, _07044_);
  nor (_07057_, _07055_, _07044_);
  nor (_07058_, _07057_, _07056_);
  not (_07059_, _07058_);
  nor (_07060_, _07059_, _07042_);
  and (_07061_, _07059_, _07042_);
  nor (_07062_, _07061_, _07060_);
  and (_07063_, _07062_, _07038_);
  nor (_07064_, _07062_, _07038_);
  nor (_07065_, _07064_, _07063_);
  and (_07066_, _07065_, _07041_);
  nor (_07067_, _07065_, _07041_);
  nor (_07068_, _07067_, _07066_);
  and (_07069_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_07070_, _07069_, _06881_);
  and (_07071_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_07072_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_07073_, _07072_, _06877_);
  nor (_07074_, _07073_, _07070_);
  and (_07075_, _07074_, _07071_);
  nor (_07076_, _07075_, _07070_);
  not (_07077_, _07076_);
  nor (_07078_, _06883_, _06879_);
  nor (_07079_, _07078_, _06884_);
  and (_07080_, _07079_, _07077_);
  and (_07081_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_07082_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_07083_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_07084_, _07083_, _07082_);
  nor (_07085_, _07083_, _07082_);
  nor (_07086_, _07085_, _07084_);
  and (_07087_, _07086_, _07081_);
  nor (_07088_, _07086_, _07081_);
  nor (_07089_, _07088_, _07087_);
  nor (_07090_, _07079_, _07077_);
  nor (_07091_, _07090_, _07080_);
  and (_07092_, _07091_, _07089_);
  nor (_07093_, _07092_, _07080_);
  nor (_07094_, _06903_, _06901_);
  nor (_07095_, _07094_, _06904_);
  not (_07096_, _07095_);
  nor (_07097_, _07096_, _07093_);
  and (_07098_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_07099_, _07098_, _06924_);
  nor (_07100_, _07087_, _07084_);
  nor (_07101_, _06924_, _06923_);
  nor (_07102_, _07101_, _06925_);
  not (_07103_, _07102_);
  nor (_07104_, _07103_, _07100_);
  and (_07105_, _07103_, _07100_);
  nor (_07106_, _07105_, _07104_);
  and (_07107_, _07106_, _07099_);
  nor (_07108_, _07106_, _07099_);
  nor (_07109_, _07108_, _07107_);
  and (_07110_, _07096_, _07093_);
  nor (_07111_, _07110_, _07097_);
  and (_07112_, _07111_, _07109_);
  nor (_07113_, _07112_, _07097_);
  nor (_07114_, _06940_, _06938_);
  nor (_07115_, _07114_, _06941_);
  not (_07116_, _07115_);
  nor (_07117_, _07116_, _07113_);
  nor (_07118_, _07107_, _07104_);
  not (_07119_, _07118_);
  and (_07120_, _07116_, _07113_);
  nor (_07121_, _07120_, _07117_);
  and (_07122_, _07121_, _07119_);
  nor (_07123_, _07122_, _07117_);
  nor (_07124_, _06977_, _06975_);
  nor (_07125_, _07124_, _06978_);
  not (_07126_, _07125_);
  nor (_07127_, _07126_, _07123_);
  and (_07128_, _07012_, _06979_);
  nor (_07129_, _07128_, _07013_);
  and (_07130_, _07129_, _07127_);
  nor (_07131_, _07040_, _07013_);
  nor (_07132_, _07131_, _07041_);
  and (_07133_, _07132_, _07130_);
  and (_07134_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_07135_, _07134_, _07069_);
  and (_07136_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_07137_, _07134_, _07069_);
  nor (_07138_, _07137_, _07135_);
  and (_07139_, _07138_, _07136_);
  nor (_07140_, _07139_, _07135_);
  not (_07141_, _07140_);
  nor (_07142_, _07074_, _07071_);
  nor (_07143_, _07142_, _07075_);
  and (_07144_, _07143_, _07141_);
  and (_07145_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_07146_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_07147_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_07148_, _07147_, _07146_);
  nor (_07149_, _07147_, _07146_);
  nor (_07150_, _07149_, _07148_);
  and (_07151_, _07150_, _07145_);
  nor (_07152_, _07150_, _07145_);
  nor (_07153_, _07152_, _07151_);
  nor (_07154_, _07143_, _07141_);
  nor (_07155_, _07154_, _07144_);
  and (_07156_, _07155_, _07153_);
  nor (_07157_, _07156_, _07144_);
  not (_07158_, _07157_);
  nor (_07159_, _07091_, _07089_);
  nor (_07160_, _07159_, _07092_);
  and (_07161_, _07160_, _07158_);
  nor (_07162_, _07151_, _07148_);
  and (_07163_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_07164_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_07165_, _07164_, _07163_);
  nor (_07166_, _07165_, _07099_);
  not (_07167_, _07166_);
  nor (_07168_, _07167_, _07162_);
  and (_07169_, _07167_, _07162_);
  nor (_07170_, _07169_, _07168_);
  nor (_07171_, _07160_, _07158_);
  nor (_07172_, _07171_, _07161_);
  and (_07173_, _07172_, _07170_);
  nor (_07174_, _07173_, _07161_);
  nor (_07175_, _07111_, _07109_);
  nor (_07176_, _07175_, _07112_);
  not (_07177_, _07176_);
  nor (_07178_, _07177_, _07174_);
  and (_07179_, _07177_, _07174_);
  nor (_07180_, _07179_, _07178_);
  and (_07181_, _07180_, _07168_);
  nor (_07182_, _07181_, _07178_);
  nor (_07183_, _07121_, _07119_);
  nor (_07184_, _07183_, _07122_);
  not (_07185_, _07184_);
  nor (_07186_, _07185_, _07182_);
  and (_07187_, _07126_, _07123_);
  nor (_07188_, _07187_, _07127_);
  and (_07189_, _07188_, _07186_);
  nor (_07190_, _07129_, _07127_);
  nor (_07191_, _07190_, _07130_);
  and (_07192_, _07191_, _07189_);
  nor (_07193_, _07191_, _07189_);
  nor (_07194_, _07193_, _07192_);
  and (_07195_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_07196_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_07197_, _07196_, _07195_);
  and (_07198_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_07199_, _07196_, _07195_);
  nor (_07200_, _07199_, _07197_);
  and (_07201_, _07200_, _07198_);
  nor (_07202_, _07201_, _07197_);
  not (_07203_, _07202_);
  nor (_07204_, _07138_, _07136_);
  nor (_07205_, _07204_, _07139_);
  and (_07206_, _07205_, _07203_);
  and (_07207_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_07208_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_07209_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_07210_, _07209_, _07208_);
  nor (_07211_, _07209_, _07208_);
  nor (_07212_, _07211_, _07210_);
  and (_07213_, _07212_, _07207_);
  nor (_07214_, _07212_, _07207_);
  nor (_07215_, _07214_, _07213_);
  nor (_07216_, _07205_, _07203_);
  nor (_07217_, _07216_, _07206_);
  and (_07218_, _07217_, _07215_);
  nor (_07219_, _07218_, _07206_);
  not (_07220_, _07219_);
  nor (_07221_, _07155_, _07153_);
  nor (_07222_, _07221_, _07156_);
  and (_07223_, _07222_, _07220_);
  not (_07224_, _07098_);
  nor (_07225_, _07213_, _07210_);
  nor (_07226_, _07225_, _07224_);
  and (_07227_, _07225_, _07224_);
  nor (_07228_, _07227_, _07226_);
  nor (_07229_, _07222_, _07220_);
  nor (_07230_, _07229_, _07223_);
  and (_07231_, _07230_, _07228_);
  nor (_07232_, _07231_, _07223_);
  not (_07233_, _07232_);
  nor (_07234_, _07172_, _07170_);
  nor (_07235_, _07234_, _07173_);
  and (_07236_, _07235_, _07233_);
  nor (_07237_, _07235_, _07233_);
  nor (_07238_, _07237_, _07236_);
  and (_07239_, _07238_, _07226_);
  nor (_07240_, _07239_, _07236_);
  nor (_07241_, _07180_, _07168_);
  nor (_07242_, _07241_, _07181_);
  not (_07243_, _07242_);
  nor (_07244_, _07243_, _07240_);
  and (_07245_, _07185_, _07182_);
  nor (_07246_, _07245_, _07186_);
  and (_07247_, _07246_, _07244_);
  nor (_07248_, _07188_, _07186_);
  nor (_07249_, _07248_, _07189_);
  and (_07250_, _07249_, _07247_);
  nor (_07251_, _07249_, _07247_);
  nor (_07252_, _07251_, _07250_);
  and (_07253_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_07254_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_07255_, _07254_, _07253_);
  and (_07256_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07257_, _07254_, _07253_);
  nor (_07258_, _07257_, _07255_);
  and (_07259_, _07258_, _07256_);
  nor (_07260_, _07259_, _07255_);
  not (_07261_, _07260_);
  nor (_07262_, _07200_, _07198_);
  nor (_07263_, _07262_, _07201_);
  and (_07264_, _07263_, _07261_);
  and (_07265_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_07266_, _07265_, _07209_);
  and (_07267_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_07268_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_07269_, _07268_, _07267_);
  nor (_07270_, _07269_, _07266_);
  nor (_07271_, _07263_, _07261_);
  nor (_07272_, _07271_, _07264_);
  and (_07273_, _07272_, _07270_);
  nor (_07274_, _07273_, _07264_);
  not (_07275_, _07274_);
  nor (_07276_, _07217_, _07215_);
  nor (_07277_, _07276_, _07218_);
  and (_07278_, _07277_, _07275_);
  nor (_07279_, _07277_, _07275_);
  nor (_07280_, _07279_, _07278_);
  and (_07281_, _07280_, _07266_);
  nor (_07282_, _07281_, _07278_);
  not (_07283_, _07282_);
  nor (_07284_, _07230_, _07228_);
  nor (_07285_, _07284_, _07231_);
  and (_07286_, _07285_, _07283_);
  nor (_07287_, _07238_, _07226_);
  nor (_07288_, _07287_, _07239_);
  and (_07289_, _07288_, _07286_);
  and (_07290_, _07243_, _07240_);
  nor (_07291_, _07290_, _07244_);
  and (_07292_, _07291_, _07289_);
  nor (_07293_, _07246_, _07244_);
  nor (_07294_, _07293_, _07247_);
  nor (_07295_, _07294_, _07292_);
  and (_07296_, _07294_, _07292_);
  not (_07297_, _07296_);
  and (_07298_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_07299_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_07300_, _07299_, _07298_);
  and (_07301_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_07302_, _07299_, _07298_);
  nor (_07303_, _07302_, _07300_);
  and (_07304_, _07303_, _07301_);
  nor (_07305_, _07304_, _07300_);
  not (_07306_, _07305_);
  nor (_07307_, _07258_, _07256_);
  nor (_07308_, _07307_, _07259_);
  and (_07309_, _07308_, _07306_);
  nor (_07310_, _07308_, _07306_);
  nor (_07311_, _07310_, _07309_);
  and (_07312_, _07311_, _07265_);
  nor (_07313_, _07312_, _07309_);
  not (_07314_, _07313_);
  nor (_07315_, _07272_, _07270_);
  nor (_07316_, _07315_, _07273_);
  and (_07317_, _07316_, _07314_);
  nor (_07318_, _07280_, _07266_);
  nor (_07319_, _07318_, _07281_);
  and (_07320_, _07319_, _07317_);
  nor (_07321_, _07285_, _07283_);
  nor (_07322_, _07321_, _07286_);
  and (_07323_, _07322_, _07320_);
  nor (_07324_, _07288_, _07286_);
  nor (_07325_, _07324_, _07289_);
  and (_07326_, _07325_, _07323_);
  nor (_07327_, _07291_, _07289_);
  nor (_07328_, _07327_, _07292_);
  and (_07329_, _07328_, _07326_);
  and (_07330_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_07331_, _07330_, _07299_);
  nor (_07332_, _07303_, _07301_);
  nor (_07333_, _07332_, _07304_);
  and (_07334_, _07333_, _07331_);
  nor (_07335_, _07311_, _07265_);
  nor (_07336_, _07335_, _07312_);
  and (_07337_, _07336_, _07334_);
  nor (_07338_, _07316_, _07314_);
  nor (_07339_, _07338_, _07317_);
  and (_07340_, _07339_, _07337_);
  nor (_07341_, _07319_, _07317_);
  nor (_07342_, _07341_, _07320_);
  and (_07343_, _07342_, _07340_);
  nor (_07344_, _07322_, _07320_);
  nor (_07345_, _07344_, _07323_);
  and (_07346_, _07345_, _07343_);
  nor (_07347_, _07325_, _07323_);
  nor (_07348_, _07347_, _07326_);
  and (_07349_, _07348_, _07346_);
  nor (_07350_, _07328_, _07326_);
  nor (_07351_, _07350_, _07329_);
  and (_07352_, _07351_, _07349_);
  nor (_07353_, _07352_, _07329_);
  and (_07354_, _07353_, _07297_);
  nor (_07355_, _07354_, _07295_);
  and (_07356_, _07355_, _07252_);
  nor (_07357_, _07356_, _07250_);
  not (_07358_, _07357_);
  and (_07359_, _07358_, _07194_);
  nor (_07360_, _07359_, _07192_);
  not (_07361_, _07360_);
  nor (_07362_, _07132_, _07130_);
  nor (_07363_, _07362_, _07133_);
  and (_07364_, _07363_, _07361_);
  nor (_07365_, _07364_, _07133_);
  not (_07366_, _07365_);
  and (_07367_, _07366_, _07068_);
  nor (_07368_, _07367_, _07066_);
  not (_07369_, _07368_);
  and (_07370_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_07371_, _07370_);
  nor (_07372_, _07371_, _07018_);
  nor (_07373_, _07372_, _07050_);
  nor (_07374_, _07056_, _07053_);
  nor (_07375_, _07374_, _07373_);
  and (_07376_, _07374_, _07373_);
  nor (_07377_, _07376_, _07375_);
  not (_07378_, _07377_);
  nor (_07379_, _07063_, _07060_);
  and (_07380_, _07379_, _07378_);
  nor (_07381_, _07379_, _07378_);
  nor (_07382_, _07381_, _07380_);
  and (_07383_, _07382_, _07369_);
  or (_07384_, _07375_, _07047_);
  or (_07385_, _07384_, _07381_);
  or (_07386_, _07385_, _07383_);
  or (_07387_, _07386_, _06875_);
  and (_07388_, _07387_, _03710_);
  and (_07389_, _07388_, _06874_);
  not (_07390_, _06838_);
  not (_07391_, _05910_);
  nor (_07392_, _05938_, _07391_);
  or (_07393_, _07392_, _06841_);
  and (_07394_, _07393_, _03505_);
  or (_07395_, _07394_, _07390_);
  or (_07396_, _07395_, _07389_);
  and (_07397_, _07396_, _06839_);
  or (_07398_, _07397_, _04481_);
  and (_07399_, _06069_, _05248_);
  not (_07400_, _04481_);
  or (_07401_, _06829_, _07400_);
  or (_07402_, _07401_, _07399_);
  and (_07403_, _07402_, _03589_);
  and (_07404_, _07403_, _07398_);
  and (_07405_, _03603_, _03168_);
  nor (_07406_, _06363_, _06830_);
  or (_07407_, _07406_, _06829_);
  and (_07408_, _07407_, _03222_);
  or (_07409_, _07408_, _07405_);
  or (_07410_, _07409_, _07404_);
  not (_07411_, _07405_);
  not (_07412_, \oc8051_golden_model_1.B [1]);
  nor (_07413_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_07414_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and (_07415_, _07414_, _07413_);
  and (_07416_, _07415_, _07412_);
  nor (_07417_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not (_07418_, \oc8051_golden_model_1.B [0]);
  and (_07419_, _07418_, \oc8051_golden_model_1.ACC [7]);
  and (_07420_, _07419_, _07417_);
  and (_07421_, _07420_, _07416_);
  or (_07422_, _07418_, \oc8051_golden_model_1.ACC [7]);
  and (_07423_, _07422_, _07417_);
  and (_07424_, _07423_, _07416_);
  or (_07425_, _07424_, _06075_);
  not (_07426_, \oc8051_golden_model_1.B [2]);
  not (_07427_, \oc8051_golden_model_1.B [3]);
  nor (_07428_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_07429_, _07428_, _07413_);
  and (_07430_, _07429_, _07427_);
  and (_07431_, _07430_, _07426_);
  not (_07432_, _07431_);
  not (_07433_, \oc8051_golden_model_1.ACC [6]);
  and (_07434_, \oc8051_golden_model_1.B [0], _07433_);
  nor (_07435_, _07434_, _06075_);
  nor (_07436_, _07435_, _07412_);
  nor (_07437_, _07436_, _07432_);
  nor (_07438_, _07437_, _07425_);
  nor (_07439_, _07438_, _07421_);
  and (_07440_, _07437_, \oc8051_golden_model_1.B [0]);
  nor (_07441_, _07440_, _07433_);
  and (_07442_, _07441_, _07412_);
  nor (_07443_, _07441_, _07412_);
  nor (_07444_, _07443_, _07442_);
  nor (_07445_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_07446_, _07445_, _07069_);
  nor (_07447_, _07446_, \oc8051_golden_model_1.ACC [4]);
  nor (_07448_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and (_07449_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_07450_, _07449_, _07418_);
  nor (_07451_, _07450_, _07448_);
  nor (_07452_, _07451_, _07447_);
  not (_07453_, _07452_);
  and (_07454_, _07453_, _07444_);
  nor (_07455_, _07439_, \oc8051_golden_model_1.B [2]);
  nor (_07456_, _07455_, _07442_);
  not (_07457_, _07456_);
  nor (_07458_, _07457_, _07454_);
  and (_07459_, \oc8051_golden_model_1.B [2], _06075_);
  nor (_07460_, _07459_, \oc8051_golden_model_1.B [7]);
  and (_07461_, _07460_, _07415_);
  not (_07462_, _07461_);
  nor (_07463_, _07462_, _07458_);
  nor (_07464_, _07463_, _07439_);
  nor (_07465_, _07464_, _07421_);
  and (_07466_, _07429_, \oc8051_golden_model_1.ACC [7]);
  nor (_07467_, _07466_, _07430_);
  nor (_07468_, _07453_, _07444_);
  nor (_07469_, _07468_, _07454_);
  not (_07470_, _07469_);
  and (_07471_, _07470_, _07463_);
  nor (_07472_, _07463_, _07441_);
  nor (_07473_, _07472_, _07471_);
  and (_07474_, _07473_, _07426_);
  nor (_07475_, _07473_, _07426_);
  nor (_07476_, _07475_, _07474_);
  not (_07477_, _07476_);
  not (_07478_, \oc8051_golden_model_1.ACC [5]);
  nor (_07479_, _07463_, _07478_);
  and (_07480_, _07463_, _07446_);
  or (_07481_, _07480_, _07479_);
  and (_07482_, _07481_, _07412_);
  nor (_07483_, _07481_, _07412_);
  not (_07484_, \oc8051_golden_model_1.ACC [4]);
  and (_07485_, \oc8051_golden_model_1.B [0], _07484_);
  nor (_07486_, _07485_, _07483_);
  nor (_07487_, _07486_, _07482_);
  nor (_07488_, _07487_, _07477_);
  nor (_07489_, _07465_, \oc8051_golden_model_1.B [3]);
  nor (_07490_, _07489_, _07474_);
  not (_07491_, _07490_);
  nor (_07492_, _07491_, _07488_);
  nor (_07493_, _07492_, _07467_);
  nor (_07494_, _07493_, _07465_);
  nor (_07495_, _07494_, _07421_);
  not (_07496_, _07493_);
  and (_07497_, _07487_, _07477_);
  nor (_07498_, _07497_, _07488_);
  nor (_07499_, _07498_, _07496_);
  nor (_07500_, _07493_, _07473_);
  nor (_07501_, _07500_, _07499_);
  and (_07502_, _07501_, _07427_);
  nor (_07503_, _07501_, _07427_);
  nor (_07504_, _07503_, _07502_);
  not (_07505_, _07504_);
  nor (_07506_, _07493_, _07481_);
  nor (_07507_, _07483_, _07482_);
  and (_07508_, _07507_, _07485_);
  nor (_07509_, _07507_, _07485_);
  nor (_07510_, _07509_, _07508_);
  and (_07511_, _07510_, _07493_);
  or (_07512_, _07511_, _07506_);
  nor (_07513_, _07512_, \oc8051_golden_model_1.B [2]);
  and (_07514_, _07512_, \oc8051_golden_model_1.B [2]);
  nor (_07515_, _07493_, _07484_);
  nor (_07516_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_07517_, _07516_, _07195_);
  and (_07518_, _07493_, _07517_);
  or (_07519_, _07518_, _07515_);
  and (_07520_, _07519_, _07412_);
  nor (_07521_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_07522_, _07521_, _07253_);
  nor (_07523_, _07522_, \oc8051_golden_model_1.ACC [2]);
  nor (_07524_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_07525_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_07526_, _07525_, _07418_);
  nor (_07527_, _07526_, _07524_);
  nor (_07528_, _07527_, _07523_);
  not (_07529_, _07528_);
  nor (_07530_, _07519_, _07412_);
  nor (_07531_, _07530_, _07520_);
  and (_07532_, _07531_, _07529_);
  nor (_07533_, _07532_, _07520_);
  nor (_07534_, _07533_, _07514_);
  nor (_07535_, _07534_, _07513_);
  nor (_07536_, _07535_, _07505_);
  nor (_07537_, _07495_, \oc8051_golden_model_1.B [4]);
  nor (_07538_, _07537_, _07502_);
  not (_07539_, _07538_);
  nor (_07540_, _07539_, _07536_);
  not (_07541_, \oc8051_golden_model_1.B [5]);
  and (_07542_, _07428_, _07541_);
  and (_07543_, \oc8051_golden_model_1.B [4], _06075_);
  not (_07544_, _07543_);
  and (_07545_, _07544_, _07542_);
  not (_07546_, _07545_);
  nor (_07547_, _07546_, _07540_);
  nor (_07548_, _07547_, _07495_);
  nor (_07549_, _07548_, _07421_);
  not (_07550_, \oc8051_golden_model_1.B [4]);
  and (_07551_, _07535_, _07505_);
  nor (_07552_, _07551_, _07536_);
  not (_07553_, _07552_);
  and (_07554_, _07553_, _07547_);
  nor (_07555_, _07547_, _07501_);
  nor (_07556_, _07555_, _07554_);
  and (_07557_, _07556_, _07550_);
  nor (_07558_, _07556_, _07550_);
  nor (_07559_, _07558_, _07557_);
  not (_07560_, _07559_);
  nor (_07561_, _07547_, _07512_);
  nor (_07562_, _07514_, _07513_);
  and (_07563_, _07562_, _07533_);
  nor (_07564_, _07562_, _07533_);
  nor (_07565_, _07564_, _07563_);
  not (_07566_, _07565_);
  and (_07567_, _07566_, _07547_);
  nor (_07568_, _07567_, _07561_);
  nor (_07569_, _07568_, \oc8051_golden_model_1.B [3]);
  and (_07570_, _07568_, \oc8051_golden_model_1.B [3]);
  nor (_07571_, _07531_, _07529_);
  nor (_07572_, _07571_, _07532_);
  not (_07573_, _07572_);
  and (_07574_, _07573_, _07547_);
  nor (_07575_, _07547_, _07519_);
  nor (_07576_, _07575_, _07574_);
  and (_07577_, _07576_, _07426_);
  not (_07578_, \oc8051_golden_model_1.ACC [3]);
  nor (_07579_, _07547_, _07578_);
  and (_07580_, _07547_, _07522_);
  or (_07581_, _07580_, _07579_);
  and (_07582_, _07581_, _07412_);
  nor (_07583_, _07581_, _07412_);
  not (_07584_, \oc8051_golden_model_1.ACC [2]);
  and (_07585_, \oc8051_golden_model_1.B [0], _07584_);
  nor (_07586_, _07585_, _07583_);
  nor (_07587_, _07586_, _07582_);
  nor (_07588_, _07576_, _07426_);
  nor (_07589_, _07588_, _07577_);
  not (_07590_, _07589_);
  nor (_07591_, _07590_, _07587_);
  nor (_07592_, _07591_, _07577_);
  nor (_07593_, _07592_, _07570_);
  nor (_07594_, _07593_, _07569_);
  nor (_07595_, _07594_, _07560_);
  nor (_07596_, _07549_, \oc8051_golden_model_1.B [5]);
  nor (_07597_, _07596_, _07557_);
  not (_07598_, _07597_);
  nor (_07599_, _07598_, _07595_);
  not (_07600_, _07599_);
  not (_07601_, _07428_);
  and (_07602_, \oc8051_golden_model_1.B [5], _06075_);
  nor (_07603_, _07602_, _07601_);
  and (_07604_, _07603_, _07600_);
  nor (_07605_, _07604_, _07549_);
  nor (_07606_, _07605_, _07421_);
  nor (_07607_, _07606_, \oc8051_golden_model_1.B [6]);
  and (_07608_, \oc8051_golden_model_1.B [6], _06075_);
  not (_07609_, _07604_);
  and (_07610_, _07594_, _07560_);
  nor (_07611_, _07610_, _07595_);
  nor (_07612_, _07611_, _07609_);
  nor (_07613_, _07604_, _07556_);
  nor (_07614_, _07613_, _07612_);
  and (_07615_, _07614_, _07541_);
  nor (_07616_, _07614_, _07541_);
  nor (_07617_, _07616_, _07615_);
  not (_07618_, _07617_);
  nor (_07619_, _07570_, _07569_);
  nor (_07620_, _07619_, _07592_);
  and (_07621_, _07619_, _07592_);
  or (_07622_, _07621_, _07620_);
  nor (_07623_, _07622_, _07609_);
  and (_07624_, _07609_, _07568_);
  nor (_07625_, _07624_, _07623_);
  and (_07626_, _07625_, _07550_);
  nor (_07627_, _07625_, _07550_);
  and (_07628_, _07590_, _07587_);
  nor (_07629_, _07628_, _07591_);
  nor (_07630_, _07629_, _07609_);
  nor (_07631_, _07604_, _07576_);
  nor (_07632_, _07631_, _07630_);
  and (_07633_, _07632_, _07427_);
  nor (_07634_, _07583_, _07582_);
  nor (_07635_, _07634_, _07585_);
  and (_07636_, _07634_, _07585_);
  or (_07637_, _07636_, _07635_);
  nor (_07638_, _07637_, _07609_);
  nor (_07639_, _07604_, _07581_);
  nor (_07640_, _07639_, _07638_);
  and (_07641_, _07640_, _07426_);
  nor (_07642_, _07640_, _07426_);
  nor (_07643_, _07604_, _07584_);
  nor (_07644_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07645_, _07644_, _07298_);
  and (_07646_, _07604_, _07645_);
  or (_07647_, _07646_, _07643_);
  and (_07648_, _07647_, _07412_);
  and (_07649_, \oc8051_golden_model_1.B [0], _03274_);
  not (_07650_, _07649_);
  nor (_07651_, _07647_, _07412_);
  nor (_07652_, _07651_, _07648_);
  and (_07653_, _07652_, _07650_);
  nor (_07654_, _07653_, _07648_);
  nor (_07655_, _07654_, _07642_);
  nor (_07656_, _07655_, _07641_);
  nor (_07657_, _07632_, _07427_);
  nor (_07658_, _07657_, _07633_);
  not (_07659_, _07658_);
  nor (_07660_, _07659_, _07656_);
  nor (_07661_, _07660_, _07633_);
  nor (_07662_, _07661_, _07627_);
  nor (_07663_, _07662_, _07626_);
  nor (_07664_, _07663_, _07618_);
  nor (_07665_, _07664_, _07615_);
  nor (_07666_, _07665_, _07608_);
  nor (_07667_, _07666_, _07607_);
  nor (_07668_, _07667_, \oc8051_golden_model_1.B [7]);
  nor (_07669_, _07668_, _07606_);
  or (_07670_, _07669_, _07421_);
  nor (_07671_, _07670_, \oc8051_golden_model_1.B [7]);
  nor (_07672_, _07671_, _07370_);
  not (_07673_, \oc8051_golden_model_1.B [6]);
  not (_07674_, _07668_);
  and (_07675_, _07663_, _07618_);
  nor (_07676_, _07675_, _07664_);
  nor (_07677_, _07676_, _07674_);
  nor (_07678_, _07668_, _07614_);
  nor (_07679_, _07678_, _07677_);
  nor (_07680_, _07679_, _07673_);
  not (_07681_, _07680_);
  nor (_07682_, _07681_, _07672_);
  nor (_07683_, _07642_, _07641_);
  and (_07684_, _07683_, _07654_);
  nor (_07685_, _07683_, _07654_);
  or (_07686_, _07685_, _07684_);
  and (_07687_, _07686_, _07668_);
  and (_07688_, _07674_, _07640_);
  nor (_07689_, _07688_, _07687_);
  nor (_07690_, _07689_, \oc8051_golden_model_1.B [3]);
  and (_07691_, _07689_, \oc8051_golden_model_1.B [3]);
  nor (_07692_, _07691_, _07690_);
  nor (_07693_, _07652_, _07650_);
  or (_07694_, _07693_, _07653_);
  and (_07695_, _07694_, _07668_);
  nor (_07696_, _07668_, _07647_);
  nor (_07697_, _07696_, _07695_);
  nor (_07698_, _07697_, _07426_);
  and (_07699_, _07697_, _07426_);
  nor (_07700_, _07699_, _07698_);
  and (_07701_, _07700_, _07692_);
  nor (_07702_, _07668_, \oc8051_golden_model_1.ACC [1]);
  and (_07703_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07704_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  or (_07705_, _07704_, _07703_);
  and (_07706_, _07668_, _07705_);
  nor (_07707_, _07706_, _07702_);
  and (_07708_, _07707_, _07412_);
  nor (_07709_, _07707_, _07412_);
  and (_07710_, _07418_, \oc8051_golden_model_1.ACC [0]);
  not (_07711_, _07710_);
  nor (_07712_, _07711_, _07709_);
  nor (_07713_, _07712_, _07708_);
  and (_07714_, _07713_, _07701_);
  not (_07715_, _07714_);
  and (_07716_, _07698_, _07692_);
  nor (_07717_, _07716_, _07691_);
  and (_07718_, _07717_, _07715_);
  and (_07719_, _07679_, _07673_);
  nor (_07720_, _07719_, _07680_);
  not (_07721_, _07720_);
  nor (_07722_, _07721_, _07672_);
  and (_07723_, _07659_, _07656_);
  or (_07724_, _07723_, _07660_);
  and (_07725_, _07724_, _07668_);
  nor (_07726_, _07668_, _07632_);
  nor (_07727_, _07726_, _07725_);
  nor (_07728_, _07727_, _07550_);
  and (_07729_, _07727_, _07550_);
  nor (_07730_, _07729_, _07728_);
  nor (_07731_, _07627_, _07626_);
  nor (_07732_, _07731_, _07661_);
  and (_07733_, _07731_, _07661_);
  or (_07734_, _07733_, _07732_);
  and (_07735_, _07734_, _07668_);
  and (_07736_, _07674_, _07625_);
  nor (_07737_, _07736_, _07735_);
  and (_07738_, _07737_, \oc8051_golden_model_1.B [5]);
  nor (_07739_, _07737_, \oc8051_golden_model_1.B [5]);
  nor (_07740_, _07739_, _07738_);
  and (_07741_, _07740_, _07730_);
  and (_07742_, _07741_, _07722_);
  not (_07743_, _07742_);
  nor (_07744_, _07743_, _07718_);
  and (_07745_, _07606_, \oc8051_golden_model_1.B [7]);
  and (_07746_, _07740_, _07728_);
  nor (_07747_, _07746_, _07738_);
  not (_07748_, _07747_);
  and (_07749_, _07748_, _07722_);
  or (_07750_, _07749_, _07745_);
  or (_07751_, _07750_, _07744_);
  nor (_07752_, _07751_, _07682_);
  and (_07753_, \oc8051_golden_model_1.B [0], _03335_);
  not (_07754_, _07753_);
  nor (_07755_, _07709_, _07708_);
  and (_07756_, _07755_, _07754_);
  and (_07757_, _07756_, _07711_);
  and (_07758_, _07757_, _07701_);
  and (_07759_, _07758_, _07742_);
  nor (_07760_, _07759_, _07752_);
  or (_07761_, _07760_, _07421_);
  and (_07762_, _07761_, _07670_);
  or (_07763_, _07762_, _07411_);
  and (_07764_, _07763_, _07410_);
  or (_07765_, _07764_, _03601_);
  not (_07766_, _03600_);
  and (_07767_, _06171_, _05248_);
  or (_07768_, _07767_, _06829_);
  or (_07769_, _07768_, _05886_);
  and (_07770_, _07769_, _07766_);
  and (_07771_, _07770_, _07765_);
  and (_07772_, _05884_, _05248_);
  or (_07773_, _07772_, _06829_);
  and (_07774_, _07773_, _03600_);
  or (_07775_, _07774_, _03780_);
  or (_07776_, _07775_, _07771_);
  not (_07777_, _03622_);
  not (_07778_, _03780_);
  and (_07779_, _06378_, _05248_);
  or (_07780_, _07779_, _06829_);
  or (_07781_, _07780_, _07778_);
  and (_07782_, _07781_, _07777_);
  and (_07783_, _07782_, _07776_);
  or (_07784_, _06829_, _05310_);
  and (_07785_, _07768_, _03622_);
  and (_07786_, _07785_, _07784_);
  or (_07787_, _07786_, _07783_);
  and (_07788_, _07787_, _06828_);
  and (_07789_, _06849_, _03790_);
  and (_07790_, _07789_, _07784_);
  or (_07791_, _07790_, _03624_);
  or (_07792_, _07791_, _07788_);
  not (_07793_, _03785_);
  nor (_07794_, _05882_, _06830_);
  not (_07795_, _03624_);
  or (_07796_, _06829_, _07795_);
  or (_07797_, _07796_, _07794_);
  and (_07798_, _07797_, _07793_);
  and (_07799_, _07798_, _07792_);
  nor (_07800_, _06377_, _06830_);
  or (_07801_, _07800_, _06829_);
  and (_07802_, _07801_, _03785_);
  or (_07803_, _07802_, _03815_);
  or (_07804_, _07803_, _07799_);
  or (_07805_, _06846_, _04246_);
  and (_07806_, _07805_, _03823_);
  and (_07807_, _07806_, _07804_);
  and (_07808_, _06843_, _03453_);
  or (_07809_, _07808_, _03447_);
  or (_07810_, _07809_, _07807_);
  and (_07811_, _05831_, _05248_);
  or (_07812_, _06829_, _03514_);
  or (_07813_, _07812_, _07811_);
  and (_07814_, _07813_, _43000_);
  and (_07815_, _07814_, _07810_);
  or (_07816_, _07815_, _06827_);
  and (_40566_, _07816_, _41806_);
  nor (_07817_, _43000_, _06075_);
  not (_07818_, _05363_);
  and (_07819_, _06769_, \oc8051_golden_model_1.PSW [7]);
  and (_07820_, _07819_, _07818_);
  nor (_07821_, _07820_, _05204_);
  and (_07822_, _07820_, _05204_);
  nor (_07823_, _07822_, _07821_);
  and (_07824_, _07823_, \oc8051_golden_model_1.ACC [7]);
  nor (_07825_, _07823_, \oc8051_golden_model_1.ACC [7]);
  nor (_07826_, _07825_, _07824_);
  nor (_07827_, _07819_, _07818_);
  nor (_07828_, _07827_, _07820_);
  and (_07829_, _07828_, \oc8051_golden_model_1.ACC [6]);
  nor (_07830_, _07828_, _07433_);
  and (_07831_, _07828_, _07433_);
  nor (_07832_, _07831_, _07830_);
  and (_07833_, _06765_, \oc8051_golden_model_1.PSW [7]);
  and (_07834_, _07833_, _06766_);
  and (_07835_, _07834_, _06763_);
  nor (_07836_, _07835_, _06762_);
  nor (_07837_, _07836_, _07819_);
  and (_07838_, _07837_, \oc8051_golden_model_1.ACC [5]);
  nor (_07839_, _07837_, _07478_);
  and (_07840_, _07837_, _07478_);
  nor (_07841_, _07840_, _07839_);
  nor (_07842_, _07834_, _06763_);
  nor (_07843_, _07842_, _07835_);
  and (_07844_, _07843_, \oc8051_golden_model_1.ACC [4]);
  nor (_07845_, _07843_, _07484_);
  and (_07846_, _07843_, _07484_);
  nor (_07847_, _07846_, _07845_);
  not (_07848_, _05005_);
  not (_07849_, _04875_);
  and (_07850_, _06765_, _07849_);
  and (_07851_, _07850_, \oc8051_golden_model_1.PSW [7]);
  nor (_07852_, _07851_, _07848_);
  nor (_07853_, _07852_, _07834_);
  and (_07854_, _07853_, \oc8051_golden_model_1.ACC [3]);
  nor (_07855_, _07853_, _07578_);
  and (_07856_, _07853_, _07578_);
  nor (_07857_, _07856_, _07855_);
  nor (_07858_, _07833_, _07849_);
  nor (_07859_, _07858_, _07851_);
  and (_07860_, _07859_, \oc8051_golden_model_1.ACC [2]);
  nor (_07861_, _07859_, _07584_);
  and (_07862_, _07859_, _07584_);
  nor (_07863_, _07862_, _07861_);
  and (_07864_, _04620_, \oc8051_golden_model_1.PSW [7]);
  nor (_07865_, _07864_, _06764_);
  nor (_07866_, _07865_, _07833_);
  and (_07867_, _07866_, \oc8051_golden_model_1.ACC [1]);
  and (_07868_, _07866_, _03274_);
  nor (_07869_, _07866_, _03274_);
  nor (_07870_, _07869_, _07868_);
  not (_07871_, \oc8051_golden_model_1.PSW [7]);
  and (_07872_, _04634_, _07871_);
  nor (_07873_, _07872_, _07864_);
  and (_07874_, _07873_, \oc8051_golden_model_1.ACC [0]);
  not (_07875_, _07874_);
  nor (_07876_, _07875_, _07870_);
  nor (_07877_, _07876_, _07867_);
  nor (_07878_, _07877_, _07863_);
  nor (_07879_, _07878_, _07860_);
  nor (_07880_, _07879_, _07857_);
  nor (_07881_, _07880_, _07854_);
  nor (_07882_, _07881_, _07847_);
  nor (_07883_, _07882_, _07844_);
  nor (_07884_, _07883_, _07841_);
  nor (_07885_, _07884_, _07838_);
  nor (_07886_, _07885_, _07832_);
  nor (_07887_, _07886_, _07829_);
  nor (_07888_, _07887_, _07826_);
  and (_07889_, _07887_, _07826_);
  nor (_07890_, _07889_, _07888_);
  and (_07891_, _03494_, _03187_);
  not (_07892_, _07891_);
  and (_07893_, _04066_, _03187_);
  and (_07894_, _03493_, _03611_);
  nor (_07895_, _07894_, _03489_);
  nor (_07896_, _07895_, _04207_);
  nor (_07897_, _07896_, _07893_);
  and (_07898_, _07897_, _07892_);
  or (_07899_, _07898_, _07890_);
  nor (_07900_, _05254_, _06075_);
  and (_07901_, _05884_, _05254_);
  nor (_07902_, _07901_, _07900_);
  nand (_07903_, _07902_, _03600_);
  and (_07904_, _03603_, _03181_);
  not (_07905_, _07904_);
  or (_07906_, _06378_, _03779_);
  and (_07907_, _07906_, _07905_);
  not (_07908_, _05254_);
  nor (_07909_, _07908_, _05204_);
  nor (_07910_, _07909_, _07900_);
  nand (_07911_, _07910_, _07390_);
  not (_07912_, _03248_);
  and (_07913_, _03603_, _03223_);
  not (_07914_, _07913_);
  and (_07915_, _05210_, \oc8051_golden_model_1.PSW [7]);
  and (_07916_, _07915_, _05261_);
  and (_07917_, _07916_, _05237_);
  and (_07918_, _07917_, _05112_);
  nor (_07919_, _07918_, _03446_);
  and (_07920_, _07918_, _03446_);
  nor (_07921_, _07920_, _07919_);
  and (_07922_, _07921_, \oc8051_golden_model_1.ACC [7]);
  nor (_07923_, _07921_, \oc8051_golden_model_1.ACC [7]);
  nor (_07924_, _07923_, _07922_);
  nor (_07925_, _07917_, _05112_);
  nor (_07926_, _07925_, _07918_);
  nor (_07927_, _07926_, _07433_);
  and (_07928_, _07926_, _07433_);
  and (_07929_, _07916_, _05218_);
  nor (_07930_, _07929_, _05226_);
  nor (_07931_, _07930_, _07917_);
  and (_07932_, _07931_, _07478_);
  nor (_07933_, _07931_, _07478_);
  nor (_07934_, _07916_, _05218_);
  nor (_07935_, _07934_, _07929_);
  nor (_07936_, _07935_, _07484_);
  nor (_07937_, _07936_, _07933_);
  nor (_07938_, _07937_, _07932_);
  nor (_07939_, _07933_, _07932_);
  and (_07940_, _07935_, _07484_);
  nor (_07941_, _07940_, _07936_);
  and (_07942_, _07941_, _07939_);
  not (_07943_, _07942_);
  nor (_07944_, _05937_, _03756_);
  nor (_07945_, _07944_, _07916_);
  nor (_07946_, _07945_, _07578_);
  and (_07947_, _07945_, _07578_);
  nor (_07948_, _07947_, _07946_);
  nor (_07949_, _07915_, _04800_);
  nor (_07950_, _07949_, _05937_);
  nor (_07951_, _07950_, _07584_);
  and (_07952_, _07950_, _07584_);
  nor (_07953_, _07952_, _07951_);
  and (_07954_, _07953_, _07948_);
  nor (_07955_, _04048_, _07871_);
  nor (_07956_, _07955_, _03415_);
  nor (_07957_, _07956_, _07915_);
  nor (_07958_, _07957_, _03274_);
  and (_07959_, _07957_, _03274_);
  and (_07960_, _04048_, _07871_);
  nor (_07961_, _07960_, _07955_);
  nor (_07962_, _07961_, _03335_);
  not (_07963_, _07962_);
  nor (_07964_, _07963_, _07959_);
  nor (_07965_, _07964_, _07958_);
  and (_07966_, _07965_, _07954_);
  not (_07967_, _07966_);
  and (_07968_, _07952_, _07948_);
  nor (_07969_, _07968_, _07947_);
  and (_07970_, _07969_, _07967_);
  not (_07971_, _07954_);
  nor (_07972_, _07959_, _07958_);
  and (_07973_, _07961_, _03335_);
  nor (_07974_, _07962_, _07973_);
  nand (_07975_, _07974_, _07972_);
  nor (_07976_, _07975_, _07971_);
  nor (_07977_, _07976_, _07970_);
  nor (_07978_, _07977_, _07943_);
  nor (_07979_, _07978_, _07938_);
  nor (_07980_, _07979_, _07928_);
  or (_07981_, _07980_, _07927_);
  or (_07982_, _07981_, _07924_);
  nand (_07983_, _07981_, _07924_);
  and (_07984_, _07983_, _07982_);
  or (_07985_, _07984_, _07914_);
  and (_07986_, _06791_, \oc8051_golden_model_1.PSW [7]);
  nor (_07987_, _07986_, _06410_);
  and (_07988_, _07986_, _06410_);
  nor (_07989_, _07988_, _07987_);
  and (_07990_, _07989_, \oc8051_golden_model_1.ACC [7]);
  nor (_07991_, _07989_, \oc8051_golden_model_1.ACC [7]);
  nor (_07992_, _07991_, _07990_);
  not (_07993_, _07992_);
  and (_07994_, _06790_, \oc8051_golden_model_1.PSW [7]);
  nor (_07995_, _07994_, _06455_);
  nor (_07996_, _07995_, _07986_);
  nor (_07997_, _07996_, _07433_);
  and (_07998_, _07996_, _07433_);
  and (_07999_, _06788_, _06730_);
  and (_08000_, _07999_, \oc8051_golden_model_1.PSW [7]);
  nor (_08001_, _08000_, _06684_);
  nor (_08002_, _08001_, _07994_);
  and (_08003_, _08002_, _07478_);
  nor (_08004_, _08002_, _07478_);
  and (_08005_, _06786_, \oc8051_golden_model_1.PSW [7]);
  and (_08006_, _08005_, _06787_);
  nor (_08007_, _08006_, _06730_);
  nor (_08008_, _08007_, _08000_);
  nor (_08009_, _08008_, _07484_);
  nor (_08010_, _08009_, _08004_);
  nor (_08011_, _08010_, _08003_);
  nor (_08012_, _08004_, _08003_);
  and (_08013_, _08008_, _07484_);
  nor (_08014_, _08013_, _08009_);
  and (_08015_, _08014_, _08012_);
  and (_08016_, _06786_, _06637_);
  and (_08017_, _08016_, \oc8051_golden_model_1.PSW [7]);
  nor (_08018_, _08017_, _06592_);
  nor (_08019_, _08018_, _08006_);
  nor (_08020_, _08019_, _07578_);
  and (_08021_, _08019_, _07578_);
  nor (_08022_, _08021_, _08020_);
  nor (_08023_, _08005_, _06637_);
  nor (_08024_, _08023_, _08017_);
  nor (_08025_, _08024_, _07584_);
  and (_08026_, _08024_, _07584_);
  nor (_08027_, _08026_, _08025_);
  and (_08028_, _08027_, _08022_);
  and (_08029_, _06546_, \oc8051_golden_model_1.PSW [7]);
  nor (_08030_, _08029_, _06501_);
  nor (_08031_, _08030_, _08005_);
  nor (_08032_, _08031_, _03274_);
  and (_08033_, _08031_, _03274_);
  nor (_08034_, _06546_, \oc8051_golden_model_1.PSW [7]);
  nor (_08035_, _08034_, _08029_);
  and (_08036_, _08035_, _03335_);
  nor (_08037_, _08036_, _08033_);
  or (_08038_, _08037_, _08032_);
  and (_08039_, _08038_, _08028_);
  and (_08040_, _08025_, _08022_);
  or (_08041_, _08040_, _08020_);
  nor (_08042_, _08041_, _08039_);
  not (_08043_, _08042_);
  and (_08044_, _08043_, _08015_);
  nor (_08045_, _08044_, _08011_);
  nor (_08046_, _08045_, _07998_);
  or (_08047_, _08046_, _07997_);
  and (_08048_, _08047_, _07993_);
  nor (_08049_, _08047_, _07993_);
  nor (_08050_, _08049_, _08048_);
  nor (_08051_, _03511_, _03247_);
  nand (_08052_, _08051_, _08050_);
  and (_08053_, _04058_, _03223_);
  not (_08054_, _08053_);
  and (_08055_, _04474_, _03223_);
  nor (_08056_, _04750_, _03595_);
  nor (_08057_, _08056_, _03247_);
  nor (_08058_, _08057_, _08055_);
  and (_08059_, _08058_, _08054_);
  not (_08060_, _08059_);
  not (_08061_, _04759_);
  nor (_08062_, _04751_, _03985_);
  and (_08063_, _08062_, _08061_);
  not (_08064_, _08063_);
  nand (_08065_, _08064_, _05204_);
  and (_08066_, _03603_, _03725_);
  not (_08067_, _08066_);
  or (_08068_, _08067_, _06069_);
  and (_08069_, _04081_, _03235_);
  nor (_08070_, _07894_, _03595_);
  nor (_08071_, _08070_, _03234_);
  nor (_08072_, _08071_, _04067_);
  nor (_08073_, _03511_, _03234_);
  nor (_08074_, _08073_, _03726_);
  and (_08075_, _08074_, _08072_);
  and (_08076_, _03494_, _03725_);
  not (_08077_, _08076_);
  and (_08078_, _08077_, _08075_);
  not (_08079_, _08078_);
  nand (_08080_, _08079_, _05204_);
  nor (_08081_, _04064_, _06075_);
  and (_08082_, _04064_, _06075_);
  nor (_08083_, _08082_, _08081_);
  nand (_08084_, _08083_, _08078_);
  and (_08085_, _08084_, _08080_);
  or (_08086_, _08085_, _08066_);
  and (_08087_, _08086_, _08069_);
  and (_08088_, _08087_, _08068_);
  and (_08089_, _03603_, _03609_);
  and (_08090_, _05964_, _05254_);
  nor (_08091_, _08090_, _07900_);
  nor (_08092_, _08091_, _04081_);
  or (_08093_, _08092_, _08089_);
  or (_08094_, _08093_, _08088_);
  nor (_08095_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_08096_, _08095_, _07578_);
  and (_08097_, _08096_, _07449_);
  and (_08098_, _08097_, \oc8051_golden_model_1.ACC [6]);
  and (_08099_, _08098_, \oc8051_golden_model_1.ACC [7]);
  nor (_08100_, _08098_, \oc8051_golden_model_1.ACC [7]);
  nor (_08101_, _08100_, _08099_);
  and (_08102_, _08096_, \oc8051_golden_model_1.ACC [4]);
  nor (_08103_, _08102_, \oc8051_golden_model_1.ACC [5]);
  nor (_08104_, _08103_, _08097_);
  nor (_08105_, _08097_, \oc8051_golden_model_1.ACC [6]);
  nor (_08106_, _08105_, _08098_);
  nor (_08107_, _08106_, _08104_);
  not (_08108_, _08107_);
  and (_08109_, _08108_, _08101_);
  nor (_08110_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_08111_, _08110_, _08107_);
  nor (_08112_, _08111_, _08101_);
  nor (_08113_, _08112_, _08109_);
  not (_08114_, _08113_);
  nand (_08115_, _08114_, _08089_);
  and (_08116_, _08115_, _03730_);
  and (_08117_, _08116_, _08094_);
  nor (_08118_, _05903_, _06075_);
  and (_08119_, _06095_, _05903_);
  nor (_08120_, _08119_, _08118_);
  nor (_08121_, _08120_, _04055_);
  nor (_08122_, _07910_, _03996_);
  or (_08123_, _08122_, _08064_);
  or (_08124_, _08123_, _08121_);
  or (_08125_, _08124_, _08117_);
  and (_08126_, _08125_, _08065_);
  or (_08127_, _08126_, _04443_);
  not (_08128_, _04443_);
  or (_08129_, _06069_, _08128_);
  and (_08130_, _08129_, _03737_);
  and (_08131_, _08130_, _08127_);
  and (_08132_, _03603_, _03507_);
  nor (_08133_, _06133_, _03737_);
  or (_08134_, _08133_, _08132_);
  or (_08135_, _08134_, _08131_);
  nand (_08136_, _08132_, _07578_);
  and (_08137_, _08136_, _08135_);
  or (_08138_, _08137_, _03714_);
  and (_08139_, _05952_, _05903_);
  nor (_08140_, _08139_, _08118_);
  nand (_08141_, _08140_, _03714_);
  and (_08142_, _08141_, _06840_);
  and (_08143_, _08142_, _08138_);
  and (_08144_, _08119_, _06138_);
  nor (_08145_, _08144_, _08118_);
  nor (_08146_, _08145_, _06840_);
  or (_08147_, _08146_, _06869_);
  or (_08148_, _08147_, _08143_);
  nor (_08149_, _07348_, _07346_);
  nor (_08150_, _08149_, _07349_);
  or (_08151_, _08150_, _06875_);
  and (_08152_, _08151_, _08148_);
  or (_08153_, _08152_, _08060_);
  not (_08154_, _07826_);
  nor (_08155_, _07845_, _07839_);
  nor (_08156_, _08155_, _07840_);
  and (_08157_, _07847_, _07841_);
  not (_08158_, _08157_);
  and (_08159_, _07863_, _07857_);
  nor (_08160_, _07873_, _03335_);
  not (_08161_, _08160_);
  nor (_08162_, _08161_, _07868_);
  nor (_08163_, _08162_, _07869_);
  and (_08164_, _08163_, _08159_);
  not (_08165_, _08164_);
  and (_08166_, _07862_, _07857_);
  nor (_08167_, _08166_, _07856_);
  and (_08168_, _08167_, _08165_);
  and (_08169_, _07873_, _03335_);
  nor (_08170_, _08160_, _08169_);
  and (_08171_, _08170_, _07870_);
  and (_08172_, _08171_, _08159_);
  nor (_08173_, _08172_, _08168_);
  nor (_08174_, _08173_, _08158_);
  nor (_08175_, _08174_, _08156_);
  nor (_08176_, _08175_, _07831_);
  or (_08177_, _08176_, _07830_);
  and (_08178_, _08177_, _08154_);
  nor (_08179_, _08177_, _08154_);
  or (_08180_, _08179_, _08178_);
  or (_08181_, _08180_, _08059_);
  and (_08182_, _08181_, _08153_);
  or (_08183_, _08182_, _08051_);
  and (_08184_, _08183_, _03766_);
  and (_08185_, _08184_, _08052_);
  nor (_08186_, _07913_, _03761_);
  not (_08187_, _08186_);
  and (_08188_, _06133_, _06075_);
  nor (_08189_, _06133_, _06075_);
  nor (_08190_, _08189_, _08188_);
  not (_08191_, _08190_);
  and (_08192_, _05293_, \oc8051_golden_model_1.P0INREG [6]);
  and (_08193_, _05266_, \oc8051_golden_model_1.P1INREG [6]);
  not (_08194_, _08193_);
  and (_08195_, _05235_, \oc8051_golden_model_1.P2INREG [6]);
  and (_08196_, _05239_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_08197_, _08196_, _08195_);
  and (_08198_, _08197_, _08194_);
  nand (_08199_, _08198_, _05398_);
  nor (_08200_, _08199_, _08192_);
  and (_08201_, _08200_, _05391_);
  and (_08202_, _08201_, _05381_);
  and (_08203_, _08202_, _05364_);
  and (_08204_, _08203_, \oc8051_golden_model_1.ACC [6]);
  nor (_08205_, _08203_, \oc8051_golden_model_1.ACC [6]);
  nor (_08206_, _08205_, _08204_);
  and (_08207_, _05293_, \oc8051_golden_model_1.P0INREG [5]);
  and (_08208_, _05266_, \oc8051_golden_model_1.P1INREG [5]);
  not (_08209_, _08208_);
  and (_08210_, _05235_, \oc8051_golden_model_1.P2INREG [5]);
  and (_08211_, _05239_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_08212_, _08211_, _08210_);
  and (_08213_, _08212_, _08209_);
  nand (_08214_, _08213_, _05506_);
  nor (_08215_, _08214_, _08207_);
  and (_08216_, _08215_, _05497_);
  and (_08217_, _08216_, _05491_);
  and (_08218_, _08217_, _05470_);
  and (_08219_, _08218_, \oc8051_golden_model_1.ACC [5]);
  nor (_08220_, _08218_, \oc8051_golden_model_1.ACC [5]);
  and (_08221_, _05266_, \oc8051_golden_model_1.P1INREG [4]);
  not (_08222_, _08221_);
  not (_08223_, _05799_);
  and (_08224_, _05235_, \oc8051_golden_model_1.P2INREG [4]);
  and (_08225_, _05239_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_08226_, _08225_, _08224_);
  and (_08227_, _08226_, _08223_);
  and (_08228_, _08227_, _08222_);
  and (_08229_, _05293_, \oc8051_golden_model_1.P0INREG [4]);
  not (_08230_, _08229_);
  and (_08231_, _08230_, _05819_);
  and (_08232_, _08231_, _05814_);
  and (_08233_, _08232_, _08228_);
  and (_08234_, _08233_, _05796_);
  and (_08235_, _08234_, _05778_);
  and (_08236_, _08235_, \oc8051_golden_model_1.ACC [4]);
  and (_08237_, _05293_, \oc8051_golden_model_1.P0INREG [3]);
  and (_08238_, _05266_, \oc8051_golden_model_1.P1INREG [3]);
  not (_08239_, _08238_);
  and (_08240_, _05235_, \oc8051_golden_model_1.P2INREG [3]);
  and (_08241_, _05239_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_08242_, _08241_, _08240_);
  and (_08243_, _08242_, _08239_);
  nand (_08244_, _08243_, _05555_);
  nor (_08245_, _08244_, _08237_);
  and (_08246_, _08245_, _05546_);
  and (_08247_, _08246_, _05540_);
  and (_08248_, _08247_, _05519_);
  and (_08249_, _08248_, \oc8051_golden_model_1.ACC [3]);
  nor (_08250_, _08248_, \oc8051_golden_model_1.ACC [3]);
  and (_08251_, _05235_, \oc8051_golden_model_1.P2INREG [2]);
  and (_08252_, _05239_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_08253_, _08252_, _08251_);
  and (_08254_, _05293_, \oc8051_golden_model_1.P0INREG [2]);
  and (_08255_, _05266_, \oc8051_golden_model_1.P1INREG [2]);
  nor (_08256_, _08255_, _08254_);
  and (_08257_, _08256_, _08253_);
  and (_08258_, _08257_, _05674_);
  and (_08259_, _08258_, _05715_);
  and (_08260_, _08259_, _05668_);
  and (_08261_, _08260_, \oc8051_golden_model_1.ACC [2]);
  and (_08262_, _05235_, \oc8051_golden_model_1.P2INREG [1]);
  and (_08263_, _05239_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_08264_, _08263_, _08262_);
  and (_08265_, _05293_, \oc8051_golden_model_1.P0INREG [1]);
  and (_08266_, _05266_, \oc8051_golden_model_1.P1INREG [1]);
  nor (_08267_, _08266_, _08265_);
  and (_08268_, _08267_, _08264_);
  and (_08269_, _08268_, _05574_);
  and (_08270_, _08269_, _05615_);
  and (_08271_, _08270_, _05568_);
  and (_08272_, _08271_, \oc8051_golden_model_1.ACC [1]);
  nor (_08273_, _08271_, \oc8051_golden_model_1.ACC [1]);
  and (_08274_, _05293_, \oc8051_golden_model_1.P0INREG [0]);
  and (_08275_, _05266_, \oc8051_golden_model_1.P1INREG [0]);
  not (_08276_, _08275_);
  and (_08277_, _05235_, \oc8051_golden_model_1.P2INREG [0]);
  and (_08278_, _05239_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_08279_, _08278_, _08277_);
  and (_08280_, _08279_, _08276_);
  nand (_08281_, _08280_, _05655_);
  nor (_08282_, _08281_, _08274_);
  and (_08283_, _08282_, _05646_);
  and (_08284_, _08283_, _05640_);
  and (_08285_, _08284_, _05619_);
  nor (_08286_, _08285_, \oc8051_golden_model_1.ACC [0]);
  nor (_08287_, _08286_, _08273_);
  or (_08288_, _08287_, _08272_);
  nor (_08289_, _08260_, \oc8051_golden_model_1.ACC [2]);
  nor (_08290_, _08289_, _08261_);
  and (_08291_, _08290_, _08288_);
  nor (_08292_, _08291_, _08261_);
  nor (_08293_, _08292_, _08250_);
  or (_08294_, _08293_, _08249_);
  nor (_08295_, _08235_, \oc8051_golden_model_1.ACC [4]);
  nor (_08296_, _08295_, _08236_);
  and (_08297_, _08296_, _08294_);
  nor (_08298_, _08297_, _08236_);
  nor (_08299_, _08298_, _08220_);
  or (_08300_, _08299_, _08219_);
  and (_08301_, _08300_, _08206_);
  nor (_08302_, _08301_, _08204_);
  and (_08303_, _08302_, _08191_);
  nor (_08304_, _08302_, _08191_);
  nor (_08305_, _08304_, _08303_);
  nor (_08306_, _08300_, _08206_);
  nor (_08307_, _08306_, _08301_);
  nor (_08308_, _08219_, _08220_);
  nor (_08309_, _08308_, _08298_);
  and (_08310_, _08308_, _08298_);
  or (_08311_, _08310_, _08309_);
  nor (_08312_, _08296_, _08294_);
  nor (_08313_, _08312_, _08297_);
  nor (_08314_, _08249_, _08250_);
  and (_08315_, _08314_, _08290_);
  nor (_08316_, _08272_, _08273_);
  and (_08317_, _08285_, \oc8051_golden_model_1.ACC [0]);
  nor (_08318_, _08317_, _08286_);
  and (_08319_, _08318_, _08316_);
  and (_08320_, _08319_, _08315_);
  and (_08321_, _08320_, \oc8051_golden_model_1.PSW [7]);
  not (_08322_, _08321_);
  nor (_08323_, _08322_, _08313_);
  not (_08324_, _08323_);
  nor (_08325_, _08324_, _08311_);
  not (_08326_, _08325_);
  nor (_08327_, _08326_, _08307_);
  nor (_08328_, _08327_, _08305_);
  and (_08329_, _08327_, _08305_);
  nor (_08330_, _08329_, _08328_);
  nand (_08331_, _08330_, _07914_);
  and (_08332_, _08331_, _08187_);
  or (_08333_, _08332_, _08185_);
  and (_08334_, _08333_, _07985_);
  or (_08335_, _08334_, _07912_);
  nand (_08336_, _03446_, _07912_);
  and (_08337_, _08336_, _03710_);
  and (_08338_, _08337_, _08335_);
  not (_08339_, _05903_);
  nor (_08340_, _05938_, _08339_);
  nor (_08341_, _08340_, _08118_);
  nor (_08342_, _08341_, _03710_);
  or (_08343_, _08342_, _07390_);
  or (_08344_, _08343_, _08338_);
  and (_08345_, _08344_, _07911_);
  or (_08346_, _08345_, _04481_);
  and (_08347_, _06069_, _05254_);
  nor (_08348_, _08347_, _07900_);
  nand (_08349_, _08348_, _04481_);
  and (_08350_, _08349_, _03589_);
  and (_08351_, _08350_, _08346_);
  nor (_08352_, _06363_, _07908_);
  nor (_08353_, _08352_, _07900_);
  nor (_08354_, _08353_, _03589_);
  or (_08355_, _08354_, _07405_);
  or (_08356_, _08355_, _08351_);
  or (_08357_, _07424_, _07411_);
  and (_08358_, _08357_, _08356_);
  or (_08359_, _08358_, _03216_);
  nand (_08360_, _03446_, _03216_);
  and (_08361_, _08360_, _08359_);
  or (_08362_, _08361_, _03601_);
  and (_08363_, _03603_, _03176_);
  not (_08364_, _08363_);
  and (_08365_, _06171_, _05254_);
  nor (_08366_, _08365_, _07900_);
  nand (_08367_, _08366_, _03601_);
  and (_08368_, _08367_, _08364_);
  and (_08369_, _08368_, _08362_);
  nor (_08370_, _08364_, _03446_);
  and (_08371_, _04474_, _03181_);
  or (_08372_, _08371_, _08370_);
  or (_08373_, _08372_, _08369_);
  and (_08374_, _05204_, _06075_);
  nor (_08375_, _05204_, _06075_);
  nor (_08376_, _08375_, _08374_);
  not (_08377_, _08371_);
  or (_08378_, _08377_, _08376_);
  not (_08379_, _04181_);
  and (_08380_, _03595_, _03181_);
  and (_08381_, _07894_, _03181_);
  nor (_08382_, _08381_, _08380_);
  and (_08383_, _08382_, _08379_);
  and (_08384_, _08383_, _08378_);
  and (_08385_, _08384_, _08373_);
  and (_08386_, _03494_, _03181_);
  nor (_08387_, _08386_, _04181_);
  nand (_08388_, _08387_, _08382_);
  or (_08389_, _08386_, _08376_);
  and (_08390_, _08389_, _08388_);
  or (_08391_, _08390_, _08385_);
  nor (_08392_, _03511_, _04175_);
  not (_08393_, _08392_);
  not (_08394_, _08386_);
  or (_08395_, _08394_, _08376_);
  and (_08396_, _08395_, _08393_);
  and (_08397_, _08396_, _08391_);
  nor (_08398_, _06069_, \oc8051_golden_model_1.ACC [7]);
  and (_08399_, _06069_, \oc8051_golden_model_1.ACC [7]);
  nor (_08400_, _08399_, _08398_);
  and (_08401_, _08392_, _08400_);
  or (_08402_, _08401_, _03778_);
  or (_08403_, _08402_, _08397_);
  and (_08404_, _08403_, _07907_);
  nor (_08405_, _03446_, _06075_);
  and (_08406_, _03446_, _06075_);
  nor (_08407_, _08406_, _08405_);
  and (_08408_, _08407_, _07904_);
  or (_08409_, _08408_, _03600_);
  or (_08410_, _08409_, _08404_);
  and (_08411_, _08410_, _07903_);
  or (_08412_, _08411_, _03780_);
  or (_08413_, _07900_, _07778_);
  not (_08414_, _04198_);
  and (_08415_, _03489_, _03191_);
  nor (_08416_, _08415_, _04315_);
  and (_08417_, _08416_, _08414_);
  and (_08418_, _08417_, _08413_);
  and (_08419_, _08418_, _08412_);
  nor (_08420_, _03511_, _04193_);
  not (_08421_, _08417_);
  and (_08422_, _08421_, _08375_);
  or (_08423_, _08422_, _08420_);
  or (_08424_, _08423_, _08419_);
  not (_08425_, _08420_);
  or (_08426_, _08425_, _08399_);
  and (_08427_, _08426_, _03789_);
  and (_08428_, _08427_, _08424_);
  and (_08429_, _03603_, _03191_);
  nor (_08430_, _08429_, _03788_);
  not (_08431_, _08430_);
  or (_08432_, _08429_, _06376_);
  and (_08433_, _08432_, _08431_);
  or (_08434_, _08433_, _08428_);
  not (_08435_, _08429_);
  or (_08436_, _08435_, _08405_);
  and (_08437_, _08436_, _07777_);
  and (_08438_, _08437_, _08434_);
  or (_08439_, _08366_, _06377_);
  nor (_08440_, _08439_, _07777_);
  and (_08441_, _03489_, _03200_);
  or (_08442_, _08441_, _08440_);
  or (_08443_, _08442_, _08438_);
  and (_08444_, _03493_, _03200_);
  nor (_08445_, _08444_, _08374_);
  and (_08446_, _03200_, _02962_);
  not (_08447_, _08446_);
  or (_08448_, _08447_, _08445_);
  and (_08449_, _08448_, _08443_);
  nor (_08450_, _03511_, _04190_);
  not (_08451_, _08374_);
  and (_08452_, _08444_, _08451_);
  or (_08453_, _08452_, _08450_);
  or (_08454_, _08453_, _08449_);
  nand (_08455_, _08450_, _08398_);
  and (_08456_, _08455_, _03784_);
  and (_08457_, _08456_, _08454_);
  and (_08458_, _03603_, _03200_);
  nor (_08459_, _08458_, _03783_);
  not (_08460_, _08459_);
  not (_08461_, _08458_);
  nand (_08462_, _08461_, _06377_);
  and (_08463_, _08462_, _08460_);
  or (_08464_, _08463_, _08457_);
  nand (_08465_, _08458_, _08406_);
  and (_08466_, _08465_, _07795_);
  and (_08467_, _08466_, _08464_);
  not (_08468_, _07898_);
  nor (_08469_, _05882_, _07908_);
  nor (_08470_, _08469_, _07900_);
  nor (_08471_, _08470_, _07795_);
  or (_08472_, _08471_, _08468_);
  or (_08473_, _08472_, _08467_);
  and (_08474_, _08473_, _07899_);
  nor (_08475_, _03511_, _04207_);
  or (_08476_, _08475_, _08474_);
  not (_08477_, _08475_);
  and (_08478_, _07996_, \oc8051_golden_model_1.ACC [6]);
  nor (_08479_, _07997_, _07998_);
  and (_08480_, _08002_, \oc8051_golden_model_1.ACC [5]);
  and (_08481_, _08008_, \oc8051_golden_model_1.ACC [4]);
  and (_08482_, _08019_, \oc8051_golden_model_1.ACC [3]);
  and (_08483_, _08024_, \oc8051_golden_model_1.ACC [2]);
  and (_08484_, _08031_, \oc8051_golden_model_1.ACC [1]);
  nor (_08485_, _08032_, _08033_);
  and (_08486_, _08035_, \oc8051_golden_model_1.ACC [0]);
  not (_08487_, _08486_);
  nor (_08488_, _08487_, _08485_);
  nor (_08489_, _08488_, _08484_);
  nor (_08490_, _08489_, _08027_);
  nor (_08491_, _08490_, _08483_);
  nor (_08492_, _08491_, _08022_);
  nor (_08493_, _08492_, _08482_);
  nor (_08494_, _08493_, _08014_);
  nor (_08495_, _08494_, _08481_);
  nor (_08496_, _08495_, _08012_);
  nor (_08497_, _08496_, _08480_);
  nor (_08498_, _08497_, _08479_);
  nor (_08499_, _08498_, _08478_);
  nor (_08500_, _08499_, _07992_);
  and (_08501_, _08499_, _07992_);
  nor (_08502_, _08501_, _08500_);
  or (_08503_, _08502_, _08477_);
  and (_08504_, _08503_, _03777_);
  and (_08505_, _08504_, _08476_);
  and (_08506_, _03603_, _03187_);
  nor (_08507_, _08506_, _03776_);
  not (_08508_, _08507_);
  not (_08509_, _08203_);
  not (_08510_, _08248_);
  not (_08511_, _08260_);
  not (_08512_, _08271_);
  nor (_08513_, _08285_, _07871_);
  and (_08514_, _08513_, _08512_);
  and (_08515_, _08514_, _08511_);
  and (_08516_, _08515_, _08510_);
  nor (_08517_, _08235_, _08218_);
  and (_08518_, _08517_, _08516_);
  and (_08519_, _08518_, _08509_);
  nor (_08520_, _08519_, _06133_);
  and (_08521_, _08519_, _06133_);
  nor (_08522_, _08521_, _08520_);
  and (_08523_, _08522_, \oc8051_golden_model_1.ACC [7]);
  nor (_08524_, _08522_, \oc8051_golden_model_1.ACC [7]);
  nor (_08525_, _08524_, _08523_);
  nor (_08526_, _08518_, _08509_);
  nor (_08527_, _08526_, _08519_);
  and (_08528_, _08527_, \oc8051_golden_model_1.ACC [6]);
  and (_08529_, _08527_, _07433_);
  nor (_08530_, _08527_, _07433_);
  nor (_08531_, _08530_, _08529_);
  not (_08532_, _08218_);
  not (_08533_, _08235_);
  and (_08534_, _08516_, _08533_);
  nor (_08535_, _08534_, _08532_);
  nor (_08536_, _08535_, _08518_);
  and (_08537_, _08536_, \oc8051_golden_model_1.ACC [5]);
  and (_08538_, _08536_, _07478_);
  nor (_08539_, _08536_, _07478_);
  nor (_08540_, _08539_, _08538_);
  nor (_08541_, _08516_, _08533_);
  nor (_08542_, _08541_, _08534_);
  and (_08543_, _08542_, \oc8051_golden_model_1.ACC [4]);
  nor (_08544_, _08542_, _07484_);
  and (_08545_, _08542_, _07484_);
  nor (_08546_, _08545_, _08544_);
  nor (_08547_, _08515_, _08510_);
  nor (_08548_, _08547_, _08516_);
  and (_08549_, _08548_, \oc8051_golden_model_1.ACC [3]);
  nor (_08550_, _08548_, _07578_);
  and (_08551_, _08548_, _07578_);
  nor (_08552_, _08551_, _08550_);
  nor (_08553_, _08514_, _08511_);
  nor (_08554_, _08553_, _08515_);
  and (_08555_, _08554_, \oc8051_golden_model_1.ACC [2]);
  nor (_08556_, _08554_, _07584_);
  and (_08557_, _08554_, _07584_);
  nor (_08558_, _08557_, _08556_);
  nor (_08559_, _08513_, _08512_);
  nor (_08560_, _08559_, _08514_);
  and (_08561_, _08560_, \oc8051_golden_model_1.ACC [1]);
  and (_08562_, _08560_, _03274_);
  nor (_08563_, _08560_, _03274_);
  nor (_08564_, _08563_, _08562_);
  and (_08565_, _08285_, _07871_);
  nor (_08566_, _08565_, _08513_);
  and (_08567_, _08566_, \oc8051_golden_model_1.ACC [0]);
  not (_08568_, _08567_);
  nor (_08569_, _08568_, _08564_);
  nor (_08570_, _08569_, _08561_);
  nor (_08571_, _08570_, _08558_);
  nor (_08572_, _08571_, _08555_);
  nor (_08573_, _08572_, _08552_);
  nor (_08574_, _08573_, _08549_);
  nor (_08575_, _08574_, _08546_);
  nor (_08576_, _08575_, _08543_);
  nor (_08577_, _08576_, _08540_);
  nor (_08578_, _08577_, _08537_);
  nor (_08579_, _08578_, _08531_);
  nor (_08580_, _08579_, _08528_);
  nor (_08581_, _08580_, _08525_);
  and (_08582_, _08580_, _08525_);
  nor (_08583_, _08582_, _08581_);
  or (_08584_, _08583_, _08506_);
  and (_08585_, _08584_, _08508_);
  or (_08586_, _08585_, _08505_);
  and (_08587_, _03599_, _03187_);
  not (_08588_, _08587_);
  not (_08589_, _08506_);
  and (_08590_, _07926_, \oc8051_golden_model_1.ACC [6]);
  nor (_08591_, _07927_, _07928_);
  and (_08592_, _07931_, \oc8051_golden_model_1.ACC [5]);
  and (_08593_, _07935_, \oc8051_golden_model_1.ACC [4]);
  and (_08594_, _07945_, \oc8051_golden_model_1.ACC [3]);
  and (_08595_, _07950_, \oc8051_golden_model_1.ACC [2]);
  and (_08596_, _07957_, \oc8051_golden_model_1.ACC [1]);
  and (_08597_, _07961_, \oc8051_golden_model_1.ACC [0]);
  not (_08598_, _08597_);
  nor (_08599_, _08598_, _07972_);
  nor (_08600_, _08599_, _08596_);
  nor (_08601_, _08600_, _07953_);
  nor (_08602_, _08601_, _08595_);
  nor (_08603_, _08602_, _07948_);
  nor (_08604_, _08603_, _08594_);
  nor (_08605_, _08604_, _07941_);
  nor (_08606_, _08605_, _08593_);
  nor (_08607_, _08606_, _07939_);
  nor (_08608_, _08607_, _08592_);
  nor (_08609_, _08608_, _08591_);
  nor (_08610_, _08609_, _08590_);
  nor (_08611_, _08610_, _07924_);
  and (_08612_, _08610_, _07924_);
  nor (_08613_, _08612_, _08611_);
  or (_08614_, _08613_, _08589_);
  and (_08615_, _08614_, _08588_);
  and (_08616_, _08615_, _08586_);
  nand (_08617_, _03202_, _02962_);
  not (_08618_, _08617_);
  and (_08619_, _08587_, \oc8051_golden_model_1.ACC [6]);
  nor (_08620_, _03511_, _03949_);
  or (_08621_, _08620_, _08619_);
  or (_08622_, _08621_, _08618_);
  or (_08623_, _08622_, _08616_);
  not (_08624_, _08620_);
  and (_08625_, _06455_, \oc8051_golden_model_1.ACC [6]);
  nor (_08626_, _06455_, \oc8051_golden_model_1.ACC [6]);
  nor (_08627_, _08626_, _08625_);
  and (_08628_, _06684_, \oc8051_golden_model_1.ACC [5]);
  nor (_08629_, _06684_, \oc8051_golden_model_1.ACC [5]);
  nor (_08630_, _08629_, _08628_);
  not (_08631_, _08630_);
  and (_08632_, _06730_, \oc8051_golden_model_1.ACC [4]);
  nor (_08633_, _06730_, \oc8051_golden_model_1.ACC [4]);
  nor (_08634_, _08633_, _08632_);
  and (_08635_, _06592_, \oc8051_golden_model_1.ACC [3]);
  nor (_08636_, _06591_, _06569_);
  and (_08637_, _08636_, _07578_);
  and (_08638_, _06637_, \oc8051_golden_model_1.ACC [2]);
  nor (_08639_, _06637_, \oc8051_golden_model_1.ACC [2]);
  nor (_08640_, _08639_, _08638_);
  not (_08641_, _08640_);
  and (_08642_, _06501_, \oc8051_golden_model_1.ACC [1]);
  nor (_08643_, _06501_, \oc8051_golden_model_1.ACC [1]);
  nor (_08644_, _08643_, _08642_);
  and (_08645_, _06546_, \oc8051_golden_model_1.ACC [0]);
  and (_08646_, _08645_, _08644_);
  nor (_08647_, _08646_, _08642_);
  nor (_08648_, _08647_, _08641_);
  nor (_08649_, _08648_, _08638_);
  nor (_08650_, _08649_, _08637_);
  or (_08651_, _08650_, _08635_);
  and (_08652_, _08651_, _08634_);
  nor (_08653_, _08652_, _08632_);
  nor (_08654_, _08653_, _08631_);
  or (_08655_, _08654_, _08628_);
  and (_08656_, _08655_, _08627_);
  nor (_08657_, _08656_, _08625_);
  nor (_08658_, _08657_, _08400_);
  and (_08659_, _08657_, _08400_);
  or (_08660_, _08659_, _08658_);
  or (_08661_, _08660_, _08624_);
  nor (_08662_, _05363_, _07433_);
  and (_08663_, _05363_, _07433_);
  nor (_08664_, _08663_, _08662_);
  nor (_08665_, _05469_, _07478_);
  and (_08666_, _05469_, _07478_);
  nor (_08667_, _05777_, _07484_);
  and (_08668_, _05777_, _07484_);
  nor (_08669_, _08668_, _08667_);
  not (_08670_, _08669_);
  nor (_08671_, _05005_, _07578_);
  not (_08672_, _08671_);
  and (_08673_, _05005_, _07578_);
  nor (_08674_, _04875_, _07584_);
  and (_08675_, _04875_, _07584_);
  nor (_08676_, _08675_, _08674_);
  not (_08677_, _08676_);
  and (_08678_, _06764_, \oc8051_golden_model_1.ACC [1]);
  and (_08679_, _04406_, _03274_);
  nor (_08680_, _08679_, _08678_);
  and (_08681_, _04620_, \oc8051_golden_model_1.ACC [0]);
  and (_08682_, _08681_, _08680_);
  nor (_08683_, _08682_, _08678_);
  nor (_08684_, _08683_, _08677_);
  nor (_08685_, _08684_, _08674_);
  or (_08686_, _08685_, _08673_);
  and (_08687_, _08686_, _08672_);
  nor (_08688_, _08687_, _08670_);
  nor (_08689_, _08688_, _08667_);
  nor (_08690_, _08689_, _08666_);
  or (_08691_, _08690_, _08665_);
  and (_08692_, _08691_, _08664_);
  nor (_08693_, _08692_, _08662_);
  nor (_08694_, _08693_, _08376_);
  and (_08695_, _08693_, _08376_);
  or (_08696_, _08695_, _08694_);
  or (_08697_, _08696_, _08617_);
  and (_08698_, _08697_, _03518_);
  and (_08699_, _08698_, _08661_);
  and (_08700_, _08699_, _08623_);
  and (_08701_, _03603_, _03202_);
  nor (_08702_, _08701_, _03517_);
  not (_08703_, _08702_);
  nor (_08704_, _08203_, _07433_);
  nor (_08705_, _08218_, _07478_);
  nor (_08706_, _08235_, _07484_);
  not (_08707_, _08296_);
  nor (_08708_, _08260_, _07584_);
  nor (_08709_, _08271_, _03274_);
  nor (_08710_, _08285_, _03335_);
  not (_08711_, _08710_);
  nor (_08712_, _08711_, _08316_);
  nor (_08713_, _08712_, _08709_);
  nor (_08714_, _08713_, _08290_);
  nor (_08715_, _08714_, _08708_);
  nor (_08716_, _08715_, _08248_);
  or (_08717_, _08716_, \oc8051_golden_model_1.ACC [3]);
  nand (_08718_, _08715_, _08248_);
  and (_08719_, _08718_, _08717_);
  and (_08720_, _08719_, _08707_);
  nor (_08721_, _08720_, _08706_);
  nor (_08722_, _08721_, _08308_);
  nor (_08723_, _08722_, _08705_);
  nor (_08724_, _08723_, _08206_);
  nor (_08725_, _08724_, _08704_);
  nor (_08726_, _08725_, _08190_);
  and (_08727_, _08725_, _08190_);
  or (_08728_, _08727_, _08726_);
  or (_08729_, _08728_, _08701_);
  and (_08730_, _08729_, _08703_);
  or (_08731_, _08730_, _08700_);
  and (_08732_, _03599_, _03202_);
  not (_08733_, _08732_);
  not (_08734_, _08701_);
  nor (_08735_, _03549_, _07433_);
  and (_08736_, _03549_, _07433_);
  or (_08737_, _08736_, _08735_);
  not (_08738_, _08737_);
  nor (_08739_, _03860_, _07478_);
  and (_08740_, _03860_, _07478_);
  nor (_08741_, _03486_, _07484_);
  and (_08742_, _03486_, _07484_);
  nor (_08743_, _08742_, _08741_);
  nor (_08744_, _03581_, _07578_);
  and (_08745_, _03581_, _07578_);
  nor (_08746_, _03904_, _07584_);
  and (_08747_, _03904_, _07584_);
  nor (_08748_, _08747_, _08746_);
  not (_08749_, _08748_);
  nor (_08750_, _03414_, _03274_);
  nor (_08751_, _04048_, _03335_);
  and (_08752_, _03414_, _03274_);
  nor (_08753_, _08752_, _08750_);
  and (_08754_, _08753_, _08751_);
  nor (_08755_, _08754_, _08750_);
  nor (_08756_, _08755_, _08749_);
  nor (_08757_, _08756_, _08746_);
  nor (_08758_, _08757_, _08745_);
  or (_08759_, _08758_, _08744_);
  and (_08760_, _08759_, _08743_);
  nor (_08761_, _08760_, _08741_);
  nor (_08762_, _08761_, _08740_);
  or (_08763_, _08762_, _08739_);
  and (_08764_, _08763_, _08738_);
  nor (_08765_, _08764_, _08735_);
  nor (_08766_, _08765_, _08407_);
  and (_08767_, _08765_, _08407_);
  or (_08768_, _08767_, _08766_);
  or (_08769_, _08768_, _08734_);
  and (_08770_, _08769_, _08733_);
  and (_08771_, _08770_, _08731_);
  and (_08772_, _08732_, \oc8051_golden_model_1.ACC [6]);
  or (_08773_, _08772_, _03815_);
  or (_08774_, _08773_, _08771_);
  and (_08775_, _03603_, _03197_);
  not (_08776_, _08775_);
  nand (_08777_, _08091_, _03815_);
  and (_08778_, _08777_, _08776_);
  and (_08779_, _08778_, _08774_);
  and (_08780_, _03599_, _03197_);
  nor (_08781_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08782_, _08781_, _07524_);
  and (_08783_, _08782_, _07448_);
  and (_08784_, _08783_, _07433_);
  nor (_08785_, _08784_, _06075_);
  and (_08786_, _08784_, _06075_);
  nor (_08787_, _08786_, _08785_);
  not (_08788_, _08787_);
  and (_08789_, _08788_, _08775_);
  or (_08790_, _08789_, _08780_);
  or (_08791_, _08790_, _08779_);
  nand (_08792_, _08780_, _07871_);
  and (_08793_, _08792_, _03823_);
  and (_08794_, _08793_, _08791_);
  nor (_08795_, _08140_, _03823_);
  or (_08796_, _08795_, _03447_);
  or (_08797_, _08796_, _08794_);
  and (_08798_, _03603_, _03195_);
  not (_08799_, _08798_);
  and (_08800_, _05831_, _05254_);
  nor (_08801_, _08800_, _07900_);
  nand (_08802_, _08801_, _03447_);
  and (_08803_, _08802_, _08799_);
  and (_08804_, _08803_, _08797_);
  and (_08805_, _03599_, _03195_);
  and (_08806_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08807_, _08806_, _07525_);
  nor (_08808_, _08807_, _07484_);
  and (_08809_, _08808_, \oc8051_golden_model_1.ACC [5]);
  and (_08810_, _08809_, \oc8051_golden_model_1.ACC [6]);
  nor (_08811_, _08810_, \oc8051_golden_model_1.ACC [7]);
  and (_08812_, _08810_, \oc8051_golden_model_1.ACC [7]);
  nor (_08813_, _08812_, _08811_);
  and (_08814_, _08813_, _08798_);
  or (_08815_, _08814_, _08805_);
  or (_08816_, _08815_, _08804_);
  nand (_08817_, _08805_, _03335_);
  and (_08818_, _08817_, _43000_);
  and (_08819_, _08818_, _08816_);
  or (_08820_, _08819_, _07817_);
  and (_40567_, _08820_, _41806_);
  not (_08821_, \oc8051_golden_model_1.DPL [7]);
  nor (_08822_, _43000_, _08821_);
  nor (_08823_, _05303_, _08821_);
  not (_08824_, _05303_);
  nor (_08825_, _06377_, _08824_);
  or (_08826_, _08825_, _08823_);
  and (_08827_, _08826_, _03785_);
  not (_08828_, _03602_);
  nor (_08829_, _08824_, _05204_);
  or (_08830_, _08829_, _08823_);
  or (_08831_, _08830_, _06838_);
  not (_08832_, _03625_);
  and (_08833_, _05964_, _05303_);
  or (_08834_, _08833_, _08823_);
  or (_08835_, _08834_, _04081_);
  and (_08836_, _05303_, \oc8051_golden_model_1.ACC [7]);
  or (_08837_, _08836_, _08823_);
  and (_08838_, _08837_, _04409_);
  nor (_08839_, _04409_, _08821_);
  or (_08840_, _08839_, _03610_);
  or (_08841_, _08840_, _08838_);
  and (_08842_, _08841_, _03996_);
  and (_08843_, _08842_, _08835_);
  and (_08844_, _08830_, _03723_);
  or (_08845_, _08844_, _03729_);
  or (_08846_, _08845_, _08843_);
  nor (_08847_, _03237_, _03215_);
  not (_08848_, _08847_);
  or (_08849_, _08837_, _03737_);
  and (_08850_, _08849_, _08848_);
  and (_08851_, _08850_, _08846_);
  and (_08852_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_08853_, _08852_, \oc8051_golden_model_1.DPL [2]);
  and (_08854_, _08853_, \oc8051_golden_model_1.DPL [3]);
  and (_08855_, _08854_, \oc8051_golden_model_1.DPL [4]);
  and (_08856_, _08855_, \oc8051_golden_model_1.DPL [5]);
  and (_08857_, _08856_, \oc8051_golden_model_1.DPL [6]);
  nor (_08858_, _08857_, \oc8051_golden_model_1.DPL [7]);
  and (_08859_, _08857_, \oc8051_golden_model_1.DPL [7]);
  nor (_08860_, _08859_, _08858_);
  and (_08861_, _08860_, _08847_);
  or (_08862_, _08861_, _08851_);
  and (_08863_, _08862_, _08832_);
  nor (_08864_, _05881_, _08832_);
  or (_08865_, _08864_, _07390_);
  or (_08866_, _08865_, _08863_);
  and (_08867_, _08866_, _08831_);
  or (_08868_, _08867_, _04481_);
  and (_08869_, _06069_, _05303_);
  or (_08870_, _08823_, _07400_);
  or (_08871_, _08870_, _08869_);
  and (_08872_, _08871_, _03589_);
  and (_08873_, _08872_, _08868_);
  nor (_08874_, _06363_, _08824_);
  or (_08875_, _08874_, _08823_);
  and (_08876_, _08875_, _03222_);
  or (_08877_, _08876_, _08873_);
  or (_08878_, _08877_, _08828_);
  and (_08879_, _05884_, _05303_);
  or (_08880_, _08823_, _07766_);
  or (_08881_, _08880_, _08879_);
  and (_08882_, _06171_, _05303_);
  or (_08883_, _08882_, _08823_);
  or (_08884_, _08883_, _05886_);
  and (_08885_, _08884_, _07778_);
  and (_08886_, _08885_, _08881_);
  and (_08887_, _08886_, _08878_);
  and (_08888_, _06378_, _05303_);
  or (_08889_, _08888_, _08823_);
  and (_08890_, _08889_, _03780_);
  or (_08891_, _08890_, _08887_);
  and (_08892_, _08891_, _07777_);
  or (_08893_, _08823_, _05310_);
  and (_08894_, _08883_, _03622_);
  and (_08895_, _08894_, _08893_);
  or (_08896_, _08895_, _08892_);
  and (_08897_, _08896_, _06828_);
  and (_08898_, _08837_, _03790_);
  and (_08899_, _08898_, _08893_);
  or (_08900_, _08899_, _03624_);
  or (_08901_, _08900_, _08897_);
  nor (_08902_, _05882_, _08824_);
  or (_08903_, _08823_, _07795_);
  or (_08904_, _08903_, _08902_);
  and (_08905_, _08904_, _07793_);
  and (_08906_, _08905_, _08901_);
  or (_08907_, _08906_, _08827_);
  and (_08908_, _08907_, _04246_);
  and (_08909_, _08834_, _03815_);
  or (_08910_, _08909_, _03447_);
  or (_08911_, _08910_, _08908_);
  and (_08912_, _05831_, _05303_);
  or (_08913_, _08823_, _03514_);
  or (_08914_, _08913_, _08912_);
  and (_08915_, _08914_, _43000_);
  and (_08916_, _08915_, _08911_);
  or (_08917_, _08916_, _08822_);
  and (_40568_, _08917_, _41806_);
  not (_08918_, \oc8051_golden_model_1.DPH [7]);
  nor (_08919_, _43000_, _08918_);
  nor (_08920_, _05297_, _08918_);
  not (_08921_, _05297_);
  nor (_08922_, _06377_, _08921_);
  or (_08923_, _08922_, _08920_);
  and (_08924_, _08923_, _03785_);
  nor (_08925_, _08921_, _05204_);
  or (_08926_, _08925_, _08920_);
  or (_08927_, _08926_, _06838_);
  and (_08928_, _05964_, _05297_);
  or (_08929_, _08928_, _08920_);
  or (_08930_, _08929_, _04081_);
  and (_08931_, _05297_, \oc8051_golden_model_1.ACC [7]);
  or (_08933_, _08931_, _08920_);
  and (_08934_, _08933_, _04409_);
  nor (_08935_, _04409_, _08918_);
  or (_08936_, _08935_, _03610_);
  or (_08937_, _08936_, _08934_);
  and (_08938_, _08937_, _03996_);
  and (_08939_, _08938_, _08930_);
  and (_08940_, _08926_, _03723_);
  or (_08941_, _08940_, _03729_);
  or (_08942_, _08941_, _08939_);
  or (_08944_, _08933_, _03737_);
  and (_08945_, _08944_, _08848_);
  and (_08946_, _08945_, _08942_);
  and (_08947_, _08859_, \oc8051_golden_model_1.DPH [0]);
  and (_08948_, _08947_, \oc8051_golden_model_1.DPH [1]);
  and (_08949_, _08948_, \oc8051_golden_model_1.DPH [2]);
  and (_08950_, _08949_, \oc8051_golden_model_1.DPH [3]);
  and (_08951_, _08950_, \oc8051_golden_model_1.DPH [4]);
  and (_08952_, _08951_, \oc8051_golden_model_1.DPH [5]);
  and (_08953_, _08952_, \oc8051_golden_model_1.DPH [6]);
  nor (_08955_, _08953_, _08918_);
  and (_08956_, _08953_, _08918_);
  or (_08957_, _08956_, _08955_);
  and (_08958_, _08957_, _08847_);
  or (_08959_, _08958_, _08946_);
  and (_08960_, _08959_, _08832_);
  nor (_08961_, _08832_, _03446_);
  or (_08962_, _08961_, _07390_);
  or (_08963_, _08962_, _08960_);
  and (_08964_, _08963_, _08927_);
  or (_08966_, _08964_, _04481_);
  and (_08967_, _06069_, _05297_);
  or (_08968_, _08920_, _07400_);
  or (_08969_, _08968_, _08967_);
  and (_08970_, _08969_, _03589_);
  and (_08971_, _08970_, _08966_);
  nor (_08972_, _06363_, _08921_);
  or (_08973_, _08972_, _08920_);
  and (_08974_, _08973_, _03222_);
  or (_08975_, _08974_, _08971_);
  or (_08977_, _08975_, _08828_);
  and (_08978_, _05884_, _05297_);
  or (_08979_, _08920_, _07766_);
  or (_08980_, _08979_, _08978_);
  and (_08981_, _06171_, _05297_);
  or (_08982_, _08981_, _08920_);
  or (_08983_, _08982_, _05886_);
  and (_08984_, _08983_, _07778_);
  and (_08985_, _08984_, _08980_);
  and (_08986_, _08985_, _08977_);
  and (_08988_, _06378_, _05297_);
  or (_08989_, _08988_, _08920_);
  and (_08990_, _08989_, _03780_);
  or (_08991_, _08990_, _08986_);
  and (_08992_, _08991_, _07777_);
  or (_08993_, _08920_, _05310_);
  and (_08994_, _08982_, _03622_);
  and (_08995_, _08994_, _08993_);
  or (_08996_, _08995_, _08992_);
  and (_08997_, _08996_, _06828_);
  and (_08999_, _08933_, _03790_);
  and (_09000_, _08999_, _08993_);
  or (_09001_, _09000_, _03624_);
  or (_09002_, _09001_, _08997_);
  nor (_09003_, _05882_, _08921_);
  or (_09004_, _08920_, _07795_);
  or (_09005_, _09004_, _09003_);
  and (_09006_, _09005_, _07793_);
  and (_09007_, _09006_, _09002_);
  or (_09008_, _09007_, _08924_);
  and (_09009_, _09008_, _04246_);
  and (_09010_, _08929_, _03815_);
  or (_09011_, _09010_, _03447_);
  or (_09012_, _09011_, _09009_);
  and (_09013_, _05831_, _05297_);
  or (_09014_, _08920_, _03514_);
  or (_09015_, _09014_, _09013_);
  and (_09016_, _09015_, _43000_);
  and (_09017_, _09016_, _09012_);
  or (_09018_, _09017_, _08919_);
  and (_40569_, _09018_, _41806_);
  not (_09019_, \oc8051_golden_model_1.IE [7]);
  nor (_09020_, _05229_, _09019_);
  not (_09021_, _05229_);
  nor (_09022_, _09021_, _05204_);
  nor (_09023_, _09022_, _09020_);
  and (_09024_, _09023_, _07390_);
  nor (_09025_, _05924_, _09019_);
  and (_09026_, _05952_, _05924_);
  nor (_09027_, _09026_, _09025_);
  nor (_09028_, _09027_, _03736_);
  not (_09029_, _04409_);
  and (_09030_, _05229_, \oc8051_golden_model_1.ACC [7]);
  nor (_09031_, _09030_, _09020_);
  nor (_09032_, _09031_, _09029_);
  nor (_09033_, _04409_, _09019_);
  or (_09034_, _09033_, _09032_);
  and (_09035_, _09034_, _04081_);
  and (_09036_, _05964_, _05229_);
  nor (_09037_, _09036_, _09020_);
  nor (_09038_, _09037_, _04081_);
  or (_09039_, _09038_, _09035_);
  and (_09040_, _09039_, _04055_);
  and (_09041_, _06095_, _05924_);
  nor (_09042_, _09041_, _09025_);
  nor (_09043_, _09042_, _04055_);
  or (_09044_, _09043_, _03723_);
  or (_09045_, _09044_, _09040_);
  nand (_09046_, _09023_, _03723_);
  and (_09047_, _09046_, _09045_);
  and (_09048_, _09047_, _03737_);
  nor (_09049_, _09031_, _03737_);
  or (_09050_, _09049_, _09048_);
  and (_09051_, _09050_, _03736_);
  nor (_09052_, _09051_, _09028_);
  nor (_09053_, _09052_, _03719_);
  nor (_09054_, _09025_, _06138_);
  or (_09055_, _09042_, _06840_);
  nor (_09056_, _09055_, _09054_);
  nor (_09057_, _09056_, _09053_);
  nor (_09058_, _09057_, _03505_);
  not (_09059_, _05924_);
  nor (_09060_, _05938_, _09059_);
  nor (_09061_, _09060_, _09025_);
  nor (_09062_, _09061_, _03710_);
  nor (_09063_, _09062_, _07390_);
  not (_09064_, _09063_);
  nor (_09065_, _09064_, _09058_);
  nor (_09066_, _09065_, _09024_);
  nor (_09067_, _09066_, _04481_);
  and (_09068_, _06069_, _05229_);
  nor (_09069_, _09020_, _07400_);
  not (_09070_, _09069_);
  nor (_09071_, _09070_, _09068_);
  nor (_09072_, _09071_, _03222_);
  not (_09073_, _09072_);
  nor (_09074_, _09073_, _09067_);
  nor (_09075_, _06363_, _09021_);
  nor (_09076_, _09075_, _09020_);
  nor (_09077_, _09076_, _03589_);
  or (_09078_, _09077_, _08828_);
  or (_09079_, _09078_, _09074_);
  and (_09080_, _05884_, _05229_);
  or (_09081_, _09020_, _07766_);
  or (_09082_, _09081_, _09080_);
  and (_09083_, _06171_, _05229_);
  nor (_09084_, _09083_, _09020_);
  and (_09085_, _09084_, _03601_);
  nor (_09086_, _09085_, _03780_);
  and (_09087_, _09086_, _09082_);
  and (_09088_, _09087_, _09079_);
  and (_09089_, _06378_, _05229_);
  nor (_09090_, _09089_, _09020_);
  nor (_09091_, _09090_, _07778_);
  nor (_09092_, _09091_, _09088_);
  nor (_09093_, _09092_, _03622_);
  nor (_09094_, _09020_, _05310_);
  not (_09095_, _09094_);
  nor (_09096_, _09084_, _07777_);
  and (_09097_, _09096_, _09095_);
  nor (_09098_, _09097_, _09093_);
  nor (_09099_, _09098_, _03790_);
  nor (_09100_, _09031_, _06828_);
  and (_09101_, _09100_, _09095_);
  or (_09102_, _09101_, _09099_);
  and (_09103_, _09102_, _07795_);
  nor (_09104_, _05882_, _09021_);
  nor (_09105_, _09104_, _09020_);
  nor (_09106_, _09105_, _07795_);
  or (_09107_, _09106_, _09103_);
  and (_09108_, _09107_, _07793_);
  nor (_09109_, _06377_, _09021_);
  nor (_09110_, _09109_, _09020_);
  nor (_09111_, _09110_, _07793_);
  or (_09112_, _09111_, _09108_);
  and (_09113_, _09112_, _04246_);
  nor (_09114_, _09037_, _04246_);
  or (_09115_, _09114_, _09113_);
  and (_09116_, _09115_, _03823_);
  nor (_09117_, _09027_, _03823_);
  or (_09118_, _09117_, _09116_);
  and (_09119_, _09118_, _03514_);
  and (_09120_, _05831_, _05229_);
  nor (_09121_, _09120_, _09020_);
  nor (_09122_, _09121_, _03514_);
  or (_09123_, _09122_, _09119_);
  or (_09124_, _09123_, _43004_);
  or (_09125_, _43000_, \oc8051_golden_model_1.IE [7]);
  and (_09126_, _09125_, _41806_);
  and (_40571_, _09126_, _09124_);
  not (_09127_, \oc8051_golden_model_1.IP [7]);
  nor (_09128_, _05251_, _09127_);
  not (_09129_, _05251_);
  nor (_09130_, _09129_, _05204_);
  nor (_09131_, _09130_, _09128_);
  and (_09132_, _09131_, _07390_);
  nor (_09133_, _05908_, _09127_);
  and (_09134_, _05952_, _05908_);
  nor (_09135_, _09134_, _09133_);
  nor (_09136_, _09135_, _03736_);
  and (_09137_, _05251_, \oc8051_golden_model_1.ACC [7]);
  nor (_09138_, _09137_, _09128_);
  nor (_09139_, _09138_, _09029_);
  nor (_09140_, _04409_, _09127_);
  or (_09141_, _09140_, _09139_);
  and (_09142_, _09141_, _04081_);
  and (_09143_, _05964_, _05251_);
  nor (_09144_, _09143_, _09128_);
  nor (_09145_, _09144_, _04081_);
  or (_09146_, _09145_, _09142_);
  and (_09147_, _09146_, _04055_);
  and (_09148_, _06095_, _05908_);
  nor (_09149_, _09148_, _09133_);
  nor (_09150_, _09149_, _04055_);
  or (_09151_, _09150_, _03723_);
  or (_09152_, _09151_, _09147_);
  nand (_09153_, _09131_, _03723_);
  and (_09154_, _09153_, _09152_);
  and (_09155_, _09154_, _03737_);
  nor (_09156_, _09138_, _03737_);
  or (_09157_, _09156_, _09155_);
  and (_09158_, _09157_, _03736_);
  nor (_09159_, _09158_, _09136_);
  nor (_09160_, _09159_, _03719_);
  nor (_09161_, _09133_, _06138_);
  or (_09162_, _09149_, _06840_);
  nor (_09163_, _09162_, _09161_);
  nor (_09164_, _09163_, _09160_);
  nor (_09165_, _09164_, _03505_);
  not (_09166_, _05908_);
  nor (_09167_, _05938_, _09166_);
  nor (_09168_, _09167_, _09133_);
  nor (_09169_, _09168_, _03710_);
  nor (_09170_, _09169_, _07390_);
  not (_09171_, _09170_);
  nor (_09172_, _09171_, _09165_);
  nor (_09173_, _09172_, _09132_);
  nor (_09174_, _09173_, _04481_);
  and (_09175_, _06069_, _05251_);
  nor (_09176_, _09128_, _07400_);
  not (_09177_, _09176_);
  nor (_09178_, _09177_, _09175_);
  nor (_09179_, _09178_, _03222_);
  not (_09180_, _09179_);
  nor (_09181_, _09180_, _09174_);
  nor (_09182_, _06363_, _09129_);
  nor (_09183_, _09182_, _09128_);
  nor (_09184_, _09183_, _03589_);
  or (_09185_, _09184_, _08828_);
  or (_09186_, _09185_, _09181_);
  and (_09187_, _05884_, _05251_);
  or (_09188_, _09128_, _07766_);
  or (_09189_, _09188_, _09187_);
  and (_09190_, _06171_, _05251_);
  nor (_09191_, _09190_, _09128_);
  and (_09192_, _09191_, _03601_);
  nor (_09193_, _09192_, _03780_);
  and (_09194_, _09193_, _09189_);
  and (_09195_, _09194_, _09186_);
  and (_09196_, _06378_, _05251_);
  nor (_09197_, _09196_, _09128_);
  nor (_09198_, _09197_, _07778_);
  nor (_09199_, _09198_, _09195_);
  nor (_09200_, _09199_, _03622_);
  nor (_09201_, _09128_, _05310_);
  not (_09202_, _09201_);
  nor (_09203_, _09191_, _07777_);
  and (_09204_, _09203_, _09202_);
  nor (_09205_, _09204_, _09200_);
  nor (_09206_, _09205_, _03790_);
  nor (_09207_, _09138_, _06828_);
  and (_09208_, _09207_, _09202_);
  or (_09209_, _09208_, _09206_);
  and (_09210_, _09209_, _07795_);
  nor (_09211_, _05882_, _09129_);
  nor (_09212_, _09211_, _09128_);
  nor (_09213_, _09212_, _07795_);
  or (_09214_, _09213_, _09210_);
  and (_09215_, _09214_, _07793_);
  nor (_09216_, _06377_, _09129_);
  nor (_09217_, _09216_, _09128_);
  nor (_09218_, _09217_, _07793_);
  or (_09219_, _09218_, _09215_);
  and (_09220_, _09219_, _04246_);
  nor (_09221_, _09144_, _04246_);
  or (_09222_, _09221_, _09220_);
  and (_09223_, _09222_, _03823_);
  nor (_09224_, _09135_, _03823_);
  or (_09225_, _09224_, _09223_);
  and (_09226_, _09225_, _03514_);
  and (_09227_, _05831_, _05251_);
  nor (_09228_, _09227_, _09128_);
  nor (_09229_, _09228_, _03514_);
  or (_09230_, _09229_, _09226_);
  or (_09231_, _09230_, _43004_);
  or (_09232_, _43000_, \oc8051_golden_model_1.IP [7]);
  and (_09233_, _09232_, _41806_);
  and (_40572_, _09233_, _09231_);
  not (_09234_, \oc8051_golden_model_1.P0 [7]);
  nor (_09235_, _05293_, _09234_);
  not (_09236_, _05293_);
  nor (_09237_, _09236_, _05204_);
  or (_09238_, _09237_, _09235_);
  or (_09239_, _09238_, _06838_);
  nor (_09240_, _05209_, _09234_);
  and (_09241_, _05952_, _05209_);
  or (_09242_, _09241_, _09240_);
  and (_09243_, _09242_, _03714_);
  and (_09244_, _05964_, _05293_);
  or (_09245_, _09244_, _09235_);
  or (_09246_, _09245_, _04081_);
  and (_09247_, _05293_, \oc8051_golden_model_1.ACC [7]);
  or (_09248_, _09247_, _09235_);
  and (_09249_, _09248_, _04409_);
  nor (_09250_, _04409_, _09234_);
  or (_09251_, _09250_, _03610_);
  or (_09252_, _09251_, _09249_);
  and (_09253_, _09252_, _04055_);
  and (_09254_, _09253_, _09246_);
  and (_09255_, _06095_, _05209_);
  or (_09256_, _09255_, _09240_);
  and (_09257_, _09256_, _03715_);
  or (_09258_, _09257_, _03723_);
  or (_09259_, _09258_, _09254_);
  or (_09260_, _09238_, _03996_);
  and (_09261_, _09260_, _09259_);
  or (_09262_, _09261_, _03729_);
  or (_09263_, _09248_, _03737_);
  and (_09264_, _09263_, _03736_);
  and (_09265_, _09264_, _09262_);
  or (_09266_, _09265_, _09243_);
  and (_09267_, _09266_, _06840_);
  or (_09268_, _09240_, _06138_);
  and (_09269_, _09268_, _03719_);
  and (_09270_, _09269_, _09256_);
  or (_09271_, _09270_, _09267_);
  and (_09272_, _09271_, _03710_);
  or (_09273_, _05952_, _05937_);
  and (_09274_, _09273_, _05209_);
  or (_09275_, _09274_, _09240_);
  and (_09276_, _09275_, _03505_);
  or (_09277_, _09276_, _07390_);
  or (_09278_, _09277_, _09272_);
  and (_09279_, _09278_, _09239_);
  or (_09280_, _09279_, _04481_);
  and (_09281_, _06069_, _05293_);
  or (_09282_, _09235_, _07400_);
  or (_09283_, _09282_, _09281_);
  and (_09284_, _09283_, _03589_);
  and (_09285_, _09284_, _09280_);
  and (_09286_, _06340_, \oc8051_golden_model_1.P1 [7]);
  and (_09287_, _06343_, \oc8051_golden_model_1.P0 [7]);
  and (_09288_, _06346_, \oc8051_golden_model_1.P2 [7]);
  and (_09289_, _06348_, \oc8051_golden_model_1.P3 [7]);
  or (_09290_, _09289_, _09288_);
  or (_09291_, _09290_, _09287_);
  nor (_09292_, _09291_, _09286_);
  and (_09293_, _09292_, _06358_);
  and (_09294_, _09293_, _06339_);
  nand (_09295_, _09294_, _06326_);
  or (_09296_, _09295_, _06172_);
  and (_09297_, _09296_, _05293_);
  or (_09298_, _09297_, _09235_);
  and (_09299_, _09298_, _03222_);
  or (_09300_, _09299_, _08828_);
  or (_09301_, _09300_, _09285_);
  and (_09302_, _05884_, _05293_);
  or (_09303_, _09235_, _07766_);
  or (_09304_, _09303_, _09302_);
  and (_09305_, _06171_, _05293_);
  or (_09306_, _09305_, _09235_);
  or (_09307_, _09306_, _05886_);
  and (_09308_, _09307_, _07778_);
  and (_09309_, _09308_, _09304_);
  and (_09310_, _09309_, _09301_);
  and (_09311_, _06378_, _05293_);
  or (_09312_, _09311_, _09235_);
  and (_09313_, _09312_, _03780_);
  or (_09314_, _09313_, _09310_);
  and (_09315_, _09314_, _07777_);
  or (_09316_, _09235_, _05310_);
  and (_09317_, _09306_, _03622_);
  and (_09318_, _09317_, _09316_);
  or (_09319_, _09318_, _09315_);
  and (_09320_, _09319_, _06828_);
  and (_09321_, _09248_, _03790_);
  and (_09322_, _09321_, _09316_);
  or (_09323_, _09322_, _03624_);
  or (_09324_, _09323_, _09320_);
  nor (_09325_, _05882_, _09236_);
  or (_09326_, _09235_, _07795_);
  or (_09327_, _09326_, _09325_);
  and (_09328_, _09327_, _07793_);
  and (_09329_, _09328_, _09324_);
  nor (_09330_, _06377_, _09236_);
  or (_09331_, _09330_, _09235_);
  and (_09332_, _09331_, _03785_);
  or (_09333_, _09332_, _03815_);
  or (_09334_, _09333_, _09329_);
  or (_09335_, _09245_, _04246_);
  and (_09336_, _09335_, _03823_);
  and (_09337_, _09336_, _09334_);
  and (_09338_, _09242_, _03453_);
  or (_09339_, _09338_, _03447_);
  or (_09340_, _09339_, _09337_);
  and (_09341_, _05831_, _05293_);
  or (_09342_, _09235_, _03514_);
  or (_09343_, _09342_, _09341_);
  and (_09344_, _09343_, _43000_);
  and (_09345_, _09344_, _09340_);
  nor (_09346_, _43000_, _09234_);
  or (_09347_, _09346_, rst);
  or (_40573_, _09347_, _09345_);
  not (_09348_, \oc8051_golden_model_1.P1 [7]);
  nor (_09349_, _43000_, _09348_);
  or (_09350_, _09349_, rst);
  nor (_09351_, _05266_, _09348_);
  not (_09352_, _05266_);
  nor (_09353_, _09352_, _05204_);
  or (_09354_, _09353_, _09351_);
  or (_09355_, _09354_, _06838_);
  nor (_09356_, _05916_, _09348_);
  and (_09357_, _05952_, _05916_);
  or (_09358_, _09357_, _09356_);
  and (_09359_, _09358_, _03714_);
  and (_09360_, _05964_, _05266_);
  or (_09361_, _09360_, _09351_);
  or (_09362_, _09361_, _04081_);
  and (_09363_, _05266_, \oc8051_golden_model_1.ACC [7]);
  or (_09364_, _09363_, _09351_);
  and (_09365_, _09364_, _04409_);
  nor (_09366_, _04409_, _09348_);
  or (_09367_, _09366_, _03610_);
  or (_09368_, _09367_, _09365_);
  and (_09369_, _09368_, _04055_);
  and (_09370_, _09369_, _09362_);
  and (_09371_, _06095_, _05916_);
  or (_09372_, _09371_, _09356_);
  and (_09373_, _09372_, _03715_);
  or (_09374_, _09373_, _03723_);
  or (_09375_, _09374_, _09370_);
  or (_09376_, _09354_, _03996_);
  and (_09377_, _09376_, _09375_);
  or (_09378_, _09377_, _03729_);
  or (_09379_, _09364_, _03737_);
  and (_09380_, _09379_, _03736_);
  and (_09381_, _09380_, _09378_);
  or (_09382_, _09381_, _09359_);
  and (_09383_, _09382_, _06840_);
  and (_09384_, _06139_, _05916_);
  or (_09385_, _09384_, _09356_);
  and (_09386_, _09385_, _03719_);
  or (_09387_, _09386_, _09383_);
  and (_09388_, _09387_, _03710_);
  and (_09389_, _09273_, _05916_);
  or (_09390_, _09389_, _09356_);
  and (_09391_, _09390_, _03505_);
  or (_09392_, _09391_, _07390_);
  or (_09393_, _09392_, _09388_);
  and (_09394_, _09393_, _09355_);
  or (_09395_, _09394_, _04481_);
  and (_09396_, _06069_, _05266_);
  or (_09397_, _09351_, _07400_);
  or (_09398_, _09397_, _09396_);
  and (_09399_, _09398_, _03589_);
  and (_09400_, _09399_, _09395_);
  and (_09401_, _09296_, _05266_);
  or (_09402_, _09401_, _09351_);
  and (_09403_, _09402_, _03222_);
  or (_09404_, _09403_, _08828_);
  or (_09405_, _09404_, _09400_);
  and (_09406_, _05884_, _05266_);
  or (_09407_, _09351_, _07766_);
  or (_09408_, _09407_, _09406_);
  and (_09409_, _06171_, _05266_);
  or (_09410_, _09409_, _09351_);
  or (_09411_, _09410_, _05886_);
  and (_09412_, _09411_, _07778_);
  and (_09413_, _09412_, _09408_);
  and (_09414_, _09413_, _09405_);
  and (_09415_, _06378_, _05266_);
  or (_09416_, _09415_, _09351_);
  and (_09417_, _09416_, _03780_);
  or (_09418_, _09417_, _09414_);
  and (_09419_, _09418_, _07777_);
  or (_09420_, _09351_, _05310_);
  and (_09421_, _09410_, _03622_);
  and (_09422_, _09421_, _09420_);
  or (_09423_, _09422_, _09419_);
  and (_09424_, _09423_, _06828_);
  and (_09425_, _09364_, _03790_);
  and (_09426_, _09425_, _09420_);
  or (_09427_, _09426_, _03624_);
  or (_09428_, _09427_, _09424_);
  nor (_09429_, _05882_, _09352_);
  or (_09430_, _09351_, _07795_);
  or (_09431_, _09430_, _09429_);
  and (_09432_, _09431_, _07793_);
  and (_09433_, _09432_, _09428_);
  nor (_09434_, _06377_, _09352_);
  or (_09435_, _09434_, _09351_);
  and (_09436_, _09435_, _03785_);
  or (_09437_, _09436_, _03815_);
  or (_09438_, _09437_, _09433_);
  or (_09439_, _09361_, _04246_);
  and (_09440_, _09439_, _03823_);
  and (_09441_, _09440_, _09438_);
  and (_09442_, _09358_, _03453_);
  or (_09443_, _09442_, _03447_);
  or (_09444_, _09443_, _09441_);
  and (_09445_, _05831_, _05266_);
  or (_09446_, _09351_, _03514_);
  or (_09447_, _09446_, _09445_);
  and (_09448_, _09447_, _43000_);
  and (_09449_, _09448_, _09444_);
  or (_40574_, _09449_, _09350_);
  not (_09450_, \oc8051_golden_model_1.P2 [7]);
  nor (_09451_, _43000_, _09450_);
  or (_09452_, _09451_, rst);
  nor (_09453_, _05235_, _09450_);
  not (_09454_, _05235_);
  nor (_09455_, _09454_, _05204_);
  or (_09456_, _09455_, _09453_);
  or (_09457_, _09456_, _06838_);
  nor (_09458_, _05918_, _09450_);
  and (_09459_, _05952_, _05918_);
  or (_09460_, _09459_, _09458_);
  and (_09461_, _09460_, _03714_);
  and (_09462_, _05964_, _05235_);
  or (_09463_, _09462_, _09453_);
  or (_09464_, _09463_, _04081_);
  and (_09465_, _05235_, \oc8051_golden_model_1.ACC [7]);
  or (_09466_, _09465_, _09453_);
  and (_09467_, _09466_, _04409_);
  nor (_09468_, _04409_, _09450_);
  or (_09469_, _09468_, _03610_);
  or (_09470_, _09469_, _09467_);
  and (_09471_, _09470_, _04055_);
  and (_09472_, _09471_, _09464_);
  and (_09473_, _06095_, _05918_);
  or (_09474_, _09473_, _09458_);
  and (_09475_, _09474_, _03715_);
  or (_09476_, _09475_, _03723_);
  or (_09477_, _09476_, _09472_);
  or (_09478_, _09456_, _03996_);
  and (_09479_, _09478_, _09477_);
  or (_09480_, _09479_, _03729_);
  or (_09481_, _09466_, _03737_);
  and (_09482_, _09481_, _03736_);
  and (_09483_, _09482_, _09480_);
  or (_09484_, _09483_, _09461_);
  and (_09485_, _09484_, _06840_);
  and (_09486_, _06139_, _05918_);
  or (_09487_, _09486_, _09458_);
  and (_09488_, _09487_, _03719_);
  or (_09489_, _09488_, _09485_);
  and (_09490_, _09489_, _03710_);
  and (_09491_, _09273_, _05918_);
  or (_09492_, _09491_, _09458_);
  and (_09493_, _09492_, _03505_);
  or (_09494_, _09493_, _07390_);
  or (_09495_, _09494_, _09490_);
  and (_09496_, _09495_, _09457_);
  or (_09497_, _09496_, _04481_);
  and (_09498_, _06069_, _05235_);
  or (_09499_, _09453_, _07400_);
  or (_09500_, _09499_, _09498_);
  and (_09501_, _09500_, _03589_);
  and (_09502_, _09501_, _09497_);
  and (_09503_, _09296_, _05235_);
  or (_09504_, _09503_, _09453_);
  and (_09505_, _09504_, _03222_);
  or (_09506_, _09505_, _08828_);
  or (_09507_, _09506_, _09502_);
  and (_09508_, _05884_, _05235_);
  or (_09509_, _09453_, _07766_);
  or (_09510_, _09509_, _09508_);
  and (_09511_, _06171_, _05235_);
  or (_09512_, _09511_, _09453_);
  or (_09513_, _09512_, _05886_);
  and (_09514_, _09513_, _07778_);
  and (_09515_, _09514_, _09510_);
  and (_09516_, _09515_, _09507_);
  and (_09517_, _06378_, _05235_);
  or (_09518_, _09517_, _09453_);
  and (_09519_, _09518_, _03780_);
  or (_09520_, _09519_, _09516_);
  and (_09521_, _09520_, _07777_);
  or (_09522_, _09453_, _05310_);
  and (_09523_, _09512_, _03622_);
  and (_09524_, _09523_, _09522_);
  or (_09525_, _09524_, _09521_);
  and (_09526_, _09525_, _06828_);
  and (_09527_, _09466_, _03790_);
  and (_09528_, _09527_, _09522_);
  or (_09529_, _09528_, _03624_);
  or (_09530_, _09529_, _09526_);
  nor (_09531_, _05882_, _09454_);
  or (_09532_, _09453_, _07795_);
  or (_09533_, _09532_, _09531_);
  and (_09534_, _09533_, _07793_);
  and (_09535_, _09534_, _09530_);
  nor (_09536_, _06377_, _09454_);
  or (_09537_, _09536_, _09453_);
  and (_09538_, _09537_, _03785_);
  or (_09539_, _09538_, _03815_);
  or (_09540_, _09539_, _09535_);
  or (_09541_, _09463_, _04246_);
  and (_09542_, _09541_, _03823_);
  and (_09543_, _09542_, _09540_);
  and (_09545_, _09460_, _03453_);
  or (_09546_, _09545_, _03447_);
  or (_09547_, _09546_, _09543_);
  and (_09548_, _05831_, _05235_);
  or (_09549_, _09453_, _03514_);
  or (_09550_, _09549_, _09548_);
  and (_09551_, _09550_, _43000_);
  and (_09552_, _09551_, _09547_);
  or (_40575_, _09552_, _09452_);
  not (_09553_, \oc8051_golden_model_1.P3 [7]);
  nor (_09554_, _43000_, _09553_);
  or (_09555_, _09554_, rst);
  nor (_09556_, _05239_, _09553_);
  not (_09557_, _05239_);
  nor (_09558_, _09557_, _05204_);
  or (_09559_, _09558_, _09556_);
  or (_09560_, _09559_, _06838_);
  nor (_09561_, _05929_, _09553_);
  and (_09562_, _05952_, _05929_);
  or (_09563_, _09562_, _09561_);
  and (_09565_, _09563_, _03714_);
  and (_09566_, _05964_, _05239_);
  or (_09567_, _09566_, _09556_);
  or (_09568_, _09567_, _04081_);
  and (_09569_, _05239_, \oc8051_golden_model_1.ACC [7]);
  or (_09570_, _09569_, _09556_);
  and (_09571_, _09570_, _04409_);
  nor (_09572_, _04409_, _09553_);
  or (_09573_, _09572_, _03610_);
  or (_09574_, _09573_, _09571_);
  and (_09575_, _09574_, _04055_);
  and (_09576_, _09575_, _09568_);
  and (_09577_, _06095_, _05929_);
  or (_09578_, _09577_, _09561_);
  and (_09579_, _09578_, _03715_);
  or (_09580_, _09579_, _03723_);
  or (_09581_, _09580_, _09576_);
  or (_09582_, _09559_, _03996_);
  and (_09583_, _09582_, _09581_);
  or (_09584_, _09583_, _03729_);
  or (_09585_, _09570_, _03737_);
  and (_09586_, _09585_, _03736_);
  and (_09587_, _09586_, _09584_);
  or (_09588_, _09587_, _09565_);
  and (_09589_, _09588_, _06840_);
  and (_09590_, _06139_, _05929_);
  or (_09591_, _09590_, _09561_);
  and (_09592_, _09591_, _03719_);
  or (_09593_, _09592_, _09589_);
  and (_09594_, _09593_, _03710_);
  and (_09595_, _09273_, _05929_);
  or (_09596_, _09595_, _09561_);
  and (_09597_, _09596_, _03505_);
  or (_09598_, _09597_, _07390_);
  or (_09599_, _09598_, _09594_);
  and (_09600_, _09599_, _09560_);
  or (_09601_, _09600_, _04481_);
  and (_09602_, _06069_, _05239_);
  or (_09603_, _09556_, _07400_);
  or (_09604_, _09603_, _09602_);
  and (_09605_, _09604_, _03589_);
  and (_09606_, _09605_, _09601_);
  and (_09607_, _09296_, _05239_);
  or (_09608_, _09607_, _09556_);
  and (_09609_, _09608_, _03222_);
  or (_09610_, _09609_, _08828_);
  or (_09611_, _09610_, _09606_);
  and (_09612_, _05884_, _05239_);
  or (_09613_, _09556_, _07766_);
  or (_09614_, _09613_, _09612_);
  and (_09615_, _06171_, _05239_);
  or (_09616_, _09615_, _09556_);
  or (_09617_, _09616_, _05886_);
  and (_09618_, _09617_, _07778_);
  and (_09619_, _09618_, _09614_);
  and (_09620_, _09619_, _09611_);
  and (_09621_, _06378_, _05239_);
  or (_09622_, _09621_, _09556_);
  and (_09623_, _09622_, _03780_);
  or (_09624_, _09623_, _09620_);
  and (_09625_, _09624_, _07777_);
  or (_09626_, _09556_, _05310_);
  and (_09627_, _09616_, _03622_);
  and (_09628_, _09627_, _09626_);
  or (_09629_, _09628_, _09625_);
  and (_09630_, _09629_, _06828_);
  and (_09631_, _09570_, _03790_);
  and (_09632_, _09631_, _09626_);
  or (_09633_, _09632_, _03624_);
  or (_09634_, _09633_, _09630_);
  nor (_09635_, _05882_, _09557_);
  or (_09636_, _09556_, _07795_);
  or (_09637_, _09636_, _09635_);
  and (_09638_, _09637_, _07793_);
  and (_09639_, _09638_, _09634_);
  nor (_09640_, _06377_, _09557_);
  or (_09641_, _09640_, _09556_);
  and (_09642_, _09641_, _03785_);
  or (_09643_, _09642_, _03815_);
  or (_09644_, _09643_, _09639_);
  or (_09645_, _09567_, _04246_);
  and (_09646_, _09645_, _03823_);
  and (_09647_, _09646_, _09644_);
  and (_09648_, _09563_, _03453_);
  or (_09649_, _09648_, _03447_);
  or (_09650_, _09649_, _09647_);
  and (_09651_, _05831_, _05239_);
  or (_09652_, _09556_, _03514_);
  or (_09653_, _09652_, _09651_);
  and (_09654_, _09653_, _43000_);
  and (_09655_, _09654_, _09650_);
  or (_40577_, _09655_, _09555_);
  and (_09656_, _08780_, \oc8051_golden_model_1.ACC [0]);
  nor (_09657_, _05245_, _07871_);
  and (_09658_, _06378_, _05245_);
  or (_09659_, _09658_, _09657_);
  and (_09660_, _09659_, _03780_);
  not (_09661_, _05245_);
  nor (_09662_, _06363_, _09661_);
  or (_09663_, _09662_, _09657_);
  and (_09664_, _09663_, _03222_);
  nor (_09665_, _09661_, _05204_);
  or (_09666_, _09665_, _09657_);
  or (_09667_, _09666_, _06838_);
  not (_09668_, _03752_);
  not (_09669_, _03753_);
  not (_09670_, _05302_);
  and (_09671_, _05927_, \oc8051_golden_model_1.TCON [2]);
  and (_09672_, _05910_, \oc8051_golden_model_1.B [2]);
  nor (_09673_, _09672_, _09671_);
  and (_09674_, _05908_, \oc8051_golden_model_1.IP [2]);
  not (_09675_, _09674_);
  and (_09676_, _05901_, \oc8051_golden_model_1.PSW [2]);
  and (_09677_, _05903_, \oc8051_golden_model_1.ACC [2]);
  nor (_09678_, _09677_, _09676_);
  and (_09679_, _09678_, _09675_);
  and (_09680_, _09679_, _09673_);
  and (_09681_, _05922_, \oc8051_golden_model_1.SCON [2]);
  and (_09682_, _05924_, \oc8051_golden_model_1.IE [2]);
  nor (_09683_, _09682_, _09681_);
  and (_09684_, _05209_, \oc8051_golden_model_1.P0INREG [2]);
  and (_09685_, _05918_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_09686_, _09685_, _09684_);
  and (_09687_, _05916_, \oc8051_golden_model_1.P1INREG [2]);
  and (_09688_, _05929_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_09689_, _09688_, _09687_);
  and (_09690_, _09689_, _09686_);
  and (_09691_, _09690_, _09683_);
  and (_09692_, _09691_, _09680_);
  and (_09693_, _09692_, _05668_);
  nor (_09694_, _09693_, _09670_);
  not (_09695_, _05216_);
  and (_09696_, _05901_, \oc8051_golden_model_1.PSW [1]);
  and (_09697_, _05910_, \oc8051_golden_model_1.B [1]);
  nor (_09698_, _09697_, _09696_);
  and (_09699_, _05908_, \oc8051_golden_model_1.IP [1]);
  and (_09700_, _05903_, \oc8051_golden_model_1.ACC [1]);
  nor (_09701_, _09700_, _09699_);
  and (_09702_, _09701_, _09698_);
  and (_09703_, _05929_, \oc8051_golden_model_1.P3INREG [1]);
  not (_09704_, _09703_);
  and (_09705_, _05209_, \oc8051_golden_model_1.P0INREG [1]);
  and (_09706_, _05918_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_09707_, _09706_, _09705_);
  and (_09708_, _09707_, _09704_);
  and (_09709_, _05922_, \oc8051_golden_model_1.SCON [1]);
  and (_09710_, _05924_, \oc8051_golden_model_1.IE [1]);
  nor (_09711_, _09710_, _09709_);
  and (_09712_, _05927_, \oc8051_golden_model_1.TCON [1]);
  and (_09713_, _05916_, \oc8051_golden_model_1.P1INREG [1]);
  nor (_09714_, _09713_, _09712_);
  and (_09715_, _09714_, _09711_);
  and (_09716_, _09715_, _09708_);
  and (_09717_, _09716_, _09702_);
  and (_09718_, _09717_, _05568_);
  nor (_09719_, _09718_, _09695_);
  nor (_09720_, _09719_, _09694_);
  and (_09721_, _05223_, _04800_);
  not (_09722_, _09721_);
  and (_09723_, _05901_, \oc8051_golden_model_1.PSW [4]);
  and (_09724_, _05910_, \oc8051_golden_model_1.B [4]);
  nor (_09725_, _09724_, _09723_);
  and (_09726_, _05908_, \oc8051_golden_model_1.IP [4]);
  and (_09727_, _05903_, \oc8051_golden_model_1.ACC [4]);
  nor (_09728_, _09727_, _09726_);
  and (_09729_, _09728_, _09725_);
  and (_09730_, _05922_, \oc8051_golden_model_1.SCON [4]);
  and (_09731_, _05924_, \oc8051_golden_model_1.IE [4]);
  nor (_09732_, _09731_, _09730_);
  and (_09733_, _05927_, \oc8051_golden_model_1.TCON [4]);
  and (_09734_, _05929_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_09735_, _09734_, _09733_);
  and (_09736_, _09735_, _09732_);
  and (_09737_, _05916_, \oc8051_golden_model_1.P1INREG [4]);
  not (_09738_, _09737_);
  and (_09739_, _05209_, \oc8051_golden_model_1.P0INREG [4]);
  and (_09740_, _05918_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_09741_, _09740_, _09739_);
  and (_09742_, _09741_, _09738_);
  and (_09743_, _09742_, _09736_);
  and (_09744_, _09743_, _09729_);
  and (_09745_, _09744_, _05778_);
  nor (_09746_, _09745_, _09722_);
  nor (_09747_, _05935_, _06094_);
  nor (_09748_, _09747_, _09746_);
  and (_09749_, _09748_, _09720_);
  not (_09750_, _05224_);
  and (_09751_, _05927_, \oc8051_golden_model_1.TCON [0]);
  and (_09752_, _05910_, \oc8051_golden_model_1.B [0]);
  nor (_09753_, _09752_, _09751_);
  and (_09754_, _05901_, \oc8051_golden_model_1.PSW [0]);
  not (_09755_, _09754_);
  and (_09756_, _05908_, \oc8051_golden_model_1.IP [0]);
  and (_09757_, _05903_, \oc8051_golden_model_1.ACC [0]);
  nor (_09758_, _09757_, _09756_);
  and (_09759_, _09758_, _09755_);
  and (_09760_, _09759_, _09753_);
  and (_09761_, _05922_, \oc8051_golden_model_1.SCON [0]);
  and (_09762_, _05924_, \oc8051_golden_model_1.IE [0]);
  nor (_09763_, _09762_, _09761_);
  and (_09764_, _05916_, \oc8051_golden_model_1.P1INREG [0]);
  and (_09765_, _05929_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_09766_, _09765_, _09764_);
  and (_09767_, _05209_, \oc8051_golden_model_1.P0INREG [0]);
  and (_09768_, _05918_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_09769_, _09768_, _09767_);
  and (_09770_, _09769_, _09766_);
  and (_09771_, _09770_, _09763_);
  and (_09772_, _09771_, _09760_);
  and (_09773_, _09772_, _05619_);
  nor (_09774_, _09773_, _09750_);
  and (_09775_, _05281_, _04800_);
  not (_09776_, _09775_);
  and (_09777_, _05927_, \oc8051_golden_model_1.TCON [6]);
  and (_09778_, _05910_, \oc8051_golden_model_1.B [6]);
  nor (_09779_, _09778_, _09777_);
  and (_09780_, _05901_, \oc8051_golden_model_1.PSW [6]);
  not (_09781_, _09780_);
  and (_09782_, _05908_, \oc8051_golden_model_1.IP [6]);
  and (_09783_, _05903_, \oc8051_golden_model_1.ACC [6]);
  nor (_09784_, _09783_, _09782_);
  and (_09785_, _09784_, _09781_);
  and (_09786_, _09785_, _09779_);
  and (_09787_, _05922_, \oc8051_golden_model_1.SCON [6]);
  and (_09788_, _05924_, \oc8051_golden_model_1.IE [6]);
  nor (_09789_, _09788_, _09787_);
  and (_09790_, _05209_, \oc8051_golden_model_1.P0INREG [6]);
  and (_09791_, _05918_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_09792_, _09791_, _09790_);
  and (_09793_, _05916_, \oc8051_golden_model_1.P1INREG [6]);
  and (_09794_, _05929_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_09795_, _09794_, _09793_);
  and (_09796_, _09795_, _09792_);
  and (_09797_, _09796_, _09789_);
  and (_09798_, _09797_, _09786_);
  and (_09799_, _09798_, _05364_);
  nor (_09800_, _09799_, _09776_);
  nor (_09801_, _09800_, _09774_);
  not (_09802_, _05296_);
  and (_09803_, _05901_, \oc8051_golden_model_1.PSW [3]);
  and (_09804_, _05910_, \oc8051_golden_model_1.B [3]);
  nor (_09805_, _09804_, _09803_);
  and (_09806_, _05908_, \oc8051_golden_model_1.IP [3]);
  and (_09807_, _05903_, \oc8051_golden_model_1.ACC [3]);
  nor (_09808_, _09807_, _09806_);
  and (_09809_, _09808_, _09805_);
  and (_09810_, _05929_, \oc8051_golden_model_1.P3INREG [3]);
  not (_09811_, _09810_);
  and (_09812_, _05916_, \oc8051_golden_model_1.P1INREG [3]);
  and (_09813_, _05918_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_09814_, _09813_, _09812_);
  and (_09815_, _09814_, _09811_);
  and (_09816_, _05922_, \oc8051_golden_model_1.SCON [3]);
  and (_09817_, _05924_, \oc8051_golden_model_1.IE [3]);
  nor (_09818_, _09817_, _09816_);
  and (_09819_, _05927_, \oc8051_golden_model_1.TCON [3]);
  and (_09820_, _05209_, \oc8051_golden_model_1.P0INREG [3]);
  nor (_09821_, _09820_, _09819_);
  and (_09822_, _09821_, _09818_);
  and (_09823_, _09822_, _09815_);
  and (_09824_, _09823_, _09809_);
  and (_09825_, _09824_, _05519_);
  nor (_09826_, _09825_, _09802_);
  and (_09827_, _05215_, _04800_);
  not (_09828_, _09827_);
  and (_09829_, _05922_, \oc8051_golden_model_1.SCON [5]);
  and (_09830_, _05924_, \oc8051_golden_model_1.IE [5]);
  nor (_09831_, _09830_, _09829_);
  and (_09832_, _05927_, \oc8051_golden_model_1.TCON [5]);
  and (_09833_, _05929_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_09834_, _09833_, _09832_);
  and (_09835_, _09834_, _09831_);
  and (_09836_, _05908_, \oc8051_golden_model_1.IP [5]);
  and (_09837_, _05903_, \oc8051_golden_model_1.ACC [5]);
  nor (_09838_, _09837_, _09836_);
  and (_09839_, _05901_, \oc8051_golden_model_1.PSW [5]);
  and (_09840_, _05910_, \oc8051_golden_model_1.B [5]);
  nor (_09841_, _09840_, _09839_);
  and (_09842_, _09841_, _09838_);
  and (_09843_, _05916_, \oc8051_golden_model_1.P1INREG [5]);
  and (_09844_, _05918_, \oc8051_golden_model_1.P2INREG [5]);
  and (_09845_, _05209_, \oc8051_golden_model_1.P0INREG [5]);
  or (_09846_, _09845_, _09844_);
  nor (_09847_, _09846_, _09843_);
  and (_09848_, _09847_, _09842_);
  and (_09849_, _09848_, _09835_);
  and (_09850_, _09849_, _05470_);
  nor (_09851_, _09850_, _09828_);
  nor (_09852_, _09851_, _09826_);
  and (_09853_, _09852_, _09801_);
  and (_09854_, _09853_, _09749_);
  nor (_09855_, _09854_, _09669_);
  not (_09856_, _03604_);
  not (_09857_, _08316_);
  nor (_09858_, _08317_, _09857_);
  or (_09859_, _09858_, _08273_);
  and (_09860_, _09859_, _08315_);
  and (_09861_, _08314_, _08289_);
  or (_09862_, _09861_, _08250_);
  or (_09863_, _09862_, _09860_);
  and (_09864_, _08308_, _08296_);
  and (_09865_, _08206_, _08191_);
  and (_09866_, _09865_, _09864_);
  and (_09867_, _09866_, _09863_);
  nor (_09868_, _08295_, _08220_);
  nor (_09869_, _09868_, _08219_);
  and (_09870_, _09869_, _09865_);
  nor (_09871_, _06133_, \oc8051_golden_model_1.ACC [7]);
  and (_09872_, _08205_, _08191_);
  or (_09873_, _09872_, _09871_);
  or (_09874_, _09873_, _09870_);
  or (_09875_, _09874_, _09867_);
  and (_09876_, _09866_, _08320_);
  nor (_09877_, _09876_, _04107_);
  and (_09878_, _09877_, _09875_);
  and (_09879_, _05964_, _05245_);
  or (_09880_, _09879_, _09657_);
  or (_09881_, _09880_, _04081_);
  not (_09882_, _08089_);
  and (_09883_, _05245_, \oc8051_golden_model_1.ACC [7]);
  or (_09884_, _09883_, _09657_);
  and (_09885_, _09884_, _04409_);
  nor (_09886_, _04409_, _07871_);
  or (_09887_, _09886_, _03610_);
  or (_09888_, _09887_, _09885_);
  and (_09889_, _09888_, _09882_);
  and (_09890_, _09889_, _09881_);
  nor (_09891_, _08099_, \oc8051_golden_model_1.PSW [7]);
  not (_09892_, _09891_);
  nor (_09893_, _09892_, _08109_);
  nor (_09894_, _09893_, _09882_);
  nor (_09895_, _03229_, _03215_);
  not (_09896_, _09895_);
  nand (_09897_, _09896_, _03730_);
  or (_09898_, _09897_, _09894_);
  or (_09899_, _09898_, _09890_);
  nor (_09900_, _05901_, _07871_);
  and (_09901_, _06095_, _05901_);
  or (_09902_, _09901_, _09900_);
  or (_09903_, _09902_, _04055_);
  or (_09904_, _09666_, _03996_);
  and (_09905_, _09904_, _09903_);
  and (_09906_, _09905_, _09899_);
  or (_09907_, _09906_, _03729_);
  or (_09908_, _09884_, _03737_);
  nor (_09909_, _03232_, _03215_);
  nor (_09910_, _09909_, _03714_);
  and (_09911_, _09910_, _09908_);
  and (_09912_, _09911_, _09907_);
  and (_09913_, _05952_, _05901_);
  or (_09914_, _09913_, _09900_);
  and (_09915_, _09914_, _03714_);
  or (_09916_, _09915_, _09912_);
  nor (_09917_, _03226_, _03219_);
  or (_09918_, _09917_, _09916_);
  nor (_09919_, _03511_, _03226_);
  not (_09920_, _09919_);
  not (_09921_, _09917_);
  nor (_09922_, _05005_, _03756_);
  and (_09923_, _04875_, _04800_);
  nor (_09924_, _09923_, _09922_);
  and (_09925_, _05005_, _03756_);
  nor (_09926_, _04875_, _04800_);
  nor (_09927_, _09926_, _09925_);
  and (_09928_, _09927_, _09924_);
  and (_09929_, _04406_, _03415_);
  and (_09930_, _06764_, _03414_);
  and (_09931_, _04620_, _04048_);
  or (_09932_, _09931_, _09929_);
  nor (_09933_, _09932_, _09930_);
  or (_09934_, _09933_, _09929_);
  and (_09935_, _09934_, _09928_);
  not (_09936_, _09923_);
  nor (_09937_, _09936_, _09922_);
  or (_09938_, _09937_, _09925_);
  or (_09939_, _09938_, _09935_);
  and (_09940_, _05204_, _03454_);
  not (_09941_, _09940_);
  and (_09942_, _09941_, _05205_);
  and (_09943_, _05363_, _03549_);
  nor (_09944_, _05363_, _03549_);
  or (_09945_, _09944_, _09943_);
  and (_09946_, _09945_, _09942_);
  and (_09947_, _05469_, _05226_);
  nor (_09948_, _05469_, _05226_);
  nor (_09949_, _09948_, _09947_);
  and (_09950_, _05777_, _03486_);
  nor (_09951_, _05777_, _03486_);
  or (_09952_, _09951_, _09950_);
  and (_09953_, _09952_, _09949_);
  and (_09954_, _09953_, _09946_);
  and (_09955_, _09954_, _09939_);
  and (_09956_, _05777_, _05218_);
  and (_09957_, _09949_, _09956_);
  or (_09958_, _09957_, _09947_);
  and (_09959_, _09958_, _09946_);
  and (_09960_, _05363_, _05112_);
  and (_09961_, _09942_, _09960_);
  or (_09962_, _09961_, _09940_);
  or (_09963_, _09962_, _09959_);
  nor (_09964_, _09963_, _09955_);
  and (_09965_, _04634_, _04188_);
  not (_09966_, _09965_);
  and (_09967_, _09933_, _09928_);
  and (_09968_, _09967_, _09966_);
  and (_09969_, _09968_, _09954_);
  nor (_09970_, _09969_, _09964_);
  or (_09971_, _09970_, _09921_);
  and (_09972_, _09971_, _09920_);
  and (_09973_, _09972_, _09918_);
  or (_09974_, _06592_, _03581_);
  or (_09975_, _06637_, _03904_);
  or (_09976_, _08636_, _03756_);
  and (_09977_, _09976_, _09974_);
  not (_09978_, _09977_);
  or (_09979_, _09978_, _09975_);
  nand (_09980_, _09979_, _09974_);
  nor (_09981_, _06501_, _03414_);
  nand (_09982_, _06501_, _03414_);
  and (_09983_, _06546_, _04048_);
  nor (_09984_, _09983_, _09981_);
  and (_09985_, _09984_, _09982_);
  or (_09986_, _09985_, _09981_);
  nand (_09987_, _06637_, _03904_);
  and (_09988_, _09987_, _09977_);
  and (_09989_, _09988_, _09975_);
  and (_09990_, _09989_, _09986_);
  or (_09991_, _09990_, _09980_);
  nand (_09992_, _06455_, _03549_);
  or (_09993_, _06455_, _03549_);
  nor (_09994_, _06069_, _03446_);
  nor (_09995_, _09994_, _06150_);
  and (_09996_, _09995_, _09993_);
  and (_09997_, _09996_, _09992_);
  nor (_09998_, _06730_, _03486_);
  not (_09999_, _09998_);
  nand (_10000_, _06684_, _03860_);
  and (_10001_, _10000_, _09999_);
  nor (_10002_, _06684_, _03860_);
  and (_10003_, _06730_, _03486_);
  nor (_10004_, _10003_, _10002_);
  and (_10005_, _10004_, _10001_);
  and (_10006_, _10005_, _09997_);
  and (_10007_, _10006_, _09991_);
  or (_10008_, _09998_, _10002_);
  and (_10009_, _09997_, _10008_);
  and (_10010_, _10009_, _10000_);
  nor (_10011_, _09993_, _06150_);
  or (_10012_, _10011_, _09994_);
  or (_10013_, _10012_, _10010_);
  or (_10014_, _10013_, _10007_);
  or (_10015_, _06546_, _04048_);
  and (_10016_, _09989_, _09985_);
  and (_10017_, _10016_, _10015_);
  nand (_10018_, _10017_, _10006_);
  and (_10019_, _10018_, _09919_);
  and (_10020_, _10019_, _10014_);
  or (_10021_, _10020_, _09973_);
  and (_10022_, _10021_, _04107_);
  or (_10023_, _10022_, _09878_);
  and (_10024_, _10023_, _09856_);
  nor (_10025_, _03226_, _03215_);
  nor (_10026_, _08740_, _08739_);
  nor (_10027_, _10026_, _08743_);
  nor (_10028_, _08738_, _08407_);
  and (_10029_, _10028_, _10027_);
  nor (_10030_, _08744_, _08745_);
  nor (_10031_, _10030_, _08748_);
  nor (_10032_, _03414_, \oc8051_golden_model_1.ACC [1]);
  and (_10033_, _03414_, \oc8051_golden_model_1.ACC [1]);
  and (_10034_, _04048_, \oc8051_golden_model_1.ACC [0]);
  nor (_10035_, _10034_, _10033_);
  or (_10036_, _10035_, _10032_);
  and (_10037_, _10036_, _10031_);
  nand (_10038_, _03581_, \oc8051_golden_model_1.ACC [3]);
  nor (_10039_, _03581_, \oc8051_golden_model_1.ACC [3]);
  nor (_10040_, _03904_, \oc8051_golden_model_1.ACC [2]);
  or (_10041_, _10040_, _10039_);
  and (_10042_, _10041_, _10038_);
  or (_10043_, _10042_, _10037_);
  and (_10044_, _10043_, _10029_);
  nand (_10045_, _03860_, \oc8051_golden_model_1.ACC [5]);
  nor (_10046_, _03860_, \oc8051_golden_model_1.ACC [5]);
  nor (_10047_, _03486_, \oc8051_golden_model_1.ACC [4]);
  or (_10048_, _10047_, _10046_);
  and (_10049_, _10048_, _10045_);
  and (_10050_, _10049_, _10028_);
  nor (_10051_, _03446_, \oc8051_golden_model_1.ACC [7]);
  or (_10052_, _03549_, \oc8051_golden_model_1.ACC [6]);
  nor (_10053_, _10052_, _08407_);
  or (_10054_, _10053_, _10051_);
  or (_10055_, _10054_, _10050_);
  or (_10056_, _10055_, _10044_);
  and (_10057_, _04048_, _03335_);
  nor (_10058_, _10057_, _08751_);
  nor (_10059_, _08753_, _10058_);
  and (_10060_, _10059_, _10031_);
  and (_10061_, _10060_, _10029_);
  nor (_10062_, _10061_, _09856_);
  and (_10063_, _10062_, _10056_);
  or (_10064_, _10063_, _10025_);
  or (_10065_, _10064_, _10024_);
  nand (_10066_, _10025_, \oc8051_golden_model_1.PSW [7]);
  and (_10067_, _10066_, _06840_);
  and (_10068_, _10067_, _10065_);
  or (_10069_, _09900_, _06138_);
  and (_10070_, _09902_, _03719_);
  and (_10071_, _10070_, _10069_);
  nor (_10072_, _10071_, _10068_);
  nor (_10073_, _10072_, _03718_);
  and (_10074_, _05918_, \oc8051_golden_model_1.P2 [2]);
  and (_10075_, _05929_, \oc8051_golden_model_1.P3 [2]);
  nor (_10076_, _10075_, _10074_);
  and (_10077_, _05209_, \oc8051_golden_model_1.P0 [2]);
  and (_10078_, _05916_, \oc8051_golden_model_1.P1 [2]);
  nor (_10079_, _10078_, _10077_);
  and (_10080_, _10079_, _10076_);
  and (_10081_, _10080_, _09683_);
  and (_10082_, _10081_, _09680_);
  and (_10083_, _10082_, _05668_);
  nor (_10084_, _10083_, _09670_);
  and (_10085_, _05209_, \oc8051_golden_model_1.P0 [1]);
  and (_10086_, _05916_, \oc8051_golden_model_1.P1 [1]);
  nor (_10087_, _10086_, _10085_);
  and (_10088_, _05929_, \oc8051_golden_model_1.P3 [1]);
  and (_10089_, _05918_, \oc8051_golden_model_1.P2 [1]);
  or (_10090_, _10089_, _10088_);
  nor (_10091_, _10090_, _09712_);
  and (_10092_, _10091_, _09702_);
  and (_10093_, _10092_, _09711_);
  and (_10094_, _10093_, _10087_);
  and (_10095_, _10094_, _05568_);
  nor (_10096_, _10095_, _09695_);
  nor (_10097_, _10096_, _10084_);
  and (_10098_, _05929_, \oc8051_golden_model_1.P3 [4]);
  not (_10099_, _10098_);
  and (_10100_, _05918_, \oc8051_golden_model_1.P2 [4]);
  nor (_10101_, _10100_, _09733_);
  and (_10102_, _10101_, _10099_);
  and (_10103_, _05209_, \oc8051_golden_model_1.P0 [4]);
  and (_10104_, _05916_, \oc8051_golden_model_1.P1 [4]);
  nor (_10105_, _10104_, _10103_);
  and (_10106_, _10105_, _09732_);
  and (_10107_, _10106_, _10102_);
  and (_10108_, _10107_, _09729_);
  and (_10109_, _10108_, _05778_);
  nor (_10110_, _09722_, _10109_);
  nor (_10111_, _10110_, _06137_);
  and (_10112_, _10111_, _10097_);
  and (_10113_, _05918_, \oc8051_golden_model_1.P2 [0]);
  and (_10114_, _05929_, \oc8051_golden_model_1.P3 [0]);
  nor (_10115_, _10114_, _10113_);
  and (_10116_, _05209_, \oc8051_golden_model_1.P0 [0]);
  and (_10117_, _05916_, \oc8051_golden_model_1.P1 [0]);
  nor (_10118_, _10117_, _10116_);
  and (_10119_, _10118_, _10115_);
  and (_10120_, _10119_, _09763_);
  and (_10121_, _10120_, _09760_);
  and (_10122_, _10121_, _05619_);
  nor (_10123_, _10122_, _09750_);
  and (_10124_, _05918_, \oc8051_golden_model_1.P2 [6]);
  and (_10125_, _05929_, \oc8051_golden_model_1.P3 [6]);
  nor (_10126_, _10125_, _10124_);
  and (_10127_, _05209_, \oc8051_golden_model_1.P0 [6]);
  and (_10128_, _05916_, \oc8051_golden_model_1.P1 [6]);
  nor (_10129_, _10128_, _10127_);
  and (_10130_, _10129_, _10126_);
  and (_10131_, _10130_, _09789_);
  and (_10132_, _10131_, _09786_);
  and (_10133_, _10132_, _05364_);
  nor (_10134_, _09776_, _10133_);
  nor (_10135_, _10134_, _10123_);
  and (_10136_, _05209_, \oc8051_golden_model_1.P0 [3]);
  and (_10137_, _05916_, \oc8051_golden_model_1.P1 [3]);
  nor (_10138_, _10137_, _10136_);
  and (_10139_, _05929_, \oc8051_golden_model_1.P3 [3]);
  and (_10140_, _05918_, \oc8051_golden_model_1.P2 [3]);
  or (_10141_, _10140_, _10139_);
  nor (_10142_, _10141_, _09819_);
  and (_10143_, _10142_, _09809_);
  and (_10144_, _10143_, _09818_);
  and (_10145_, _10144_, _10138_);
  and (_10146_, _10145_, _05519_);
  nor (_10147_, _10146_, _09802_);
  and (_10148_, _05209_, \oc8051_golden_model_1.P0 [5]);
  and (_10149_, _05916_, \oc8051_golden_model_1.P1 [5]);
  nor (_10150_, _10149_, _10148_);
  and (_10151_, _05929_, \oc8051_golden_model_1.P3 [5]);
  and (_10152_, _05918_, \oc8051_golden_model_1.P2 [5]);
  or (_10153_, _10152_, _10151_);
  nor (_10154_, _10153_, _09832_);
  and (_10155_, _10154_, _09842_);
  and (_10156_, _10155_, _09831_);
  and (_10157_, _10156_, _10150_);
  and (_10158_, _10157_, _05470_);
  nor (_10159_, _09828_, _10158_);
  nor (_10160_, _10159_, _10147_);
  and (_10161_, _10160_, _10135_);
  and (_10162_, _10161_, _10112_);
  and (_10163_, _03718_, \oc8051_golden_model_1.PSW [7]);
  and (_10164_, _10163_, _10162_);
  or (_10165_, _10164_, _10073_);
  nor (_10166_, _06869_, _03753_);
  and (_10167_, _10166_, _10165_);
  or (_10168_, _10167_, _09855_);
  and (_10169_, _10168_, _09668_);
  not (_10170_, _08058_);
  or (_10171_, _10162_, \oc8051_golden_model_1.PSW [7]);
  and (_10172_, _10171_, _03752_);
  or (_10173_, _10172_, _10170_);
  or (_10174_, _10173_, _10169_);
  and (_10175_, _07835_, _06762_);
  and (_10176_, _10175_, _06771_);
  and (_10177_, _07830_, _07826_);
  nor (_10178_, _10177_, _07824_);
  not (_10179_, _10178_);
  and (_10180_, _07832_, _07826_);
  not (_10181_, _10180_);
  nor (_10182_, _10181_, _08175_);
  nor (_10183_, _10182_, _10179_);
  or (_10184_, _10183_, _10176_);
  and (_10185_, _10184_, _08054_);
  or (_10186_, _10185_, _08059_);
  and (_10187_, _10186_, _10174_);
  and (_10188_, _10184_, _08053_);
  or (_10189_, _10188_, _08051_);
  or (_10190_, _10189_, _10187_);
  and (_10191_, _07997_, _07992_);
  nor (_10192_, _10191_, _07990_);
  not (_10193_, _10192_);
  and (_10194_, _08479_, _07992_);
  not (_10195_, _10194_);
  nor (_10196_, _10195_, _08045_);
  nor (_10197_, _10196_, _10193_);
  and (_10198_, _08000_, _06684_);
  and (_10199_, _10198_, _06455_);
  and (_10200_, _10199_, _06069_);
  not (_10201_, _08051_);
  or (_10202_, _10201_, _10200_);
  or (_10203_, _10202_, _10197_);
  and (_10204_, _10203_, _10190_);
  or (_10205_, _10204_, _03761_);
  and (_10206_, _08534_, _08532_);
  nand (_10207_, _10206_, _08509_);
  nor (_10208_, _10207_, _06133_);
  and (_10209_, _08530_, _08525_);
  nor (_10210_, _10209_, _08523_);
  nor (_10211_, _08544_, _08539_);
  nor (_10212_, _10211_, _08538_);
  and (_10213_, _08531_, _08525_);
  nand (_10214_, _10213_, _10212_);
  and (_10215_, _10214_, _10210_);
  and (_10216_, _08558_, _08552_);
  and (_10217_, _08566_, _03335_);
  nor (_10218_, _10217_, _08562_);
  or (_10219_, _10218_, _08563_);
  and (_10220_, _10219_, _10216_);
  and (_10221_, _08556_, _08552_);
  or (_10222_, _10221_, _08550_);
  nor (_10223_, _10222_, _10220_);
  and (_10224_, _08546_, _08540_);
  nand (_10225_, _10213_, _10224_);
  or (_10226_, _10225_, _10223_);
  and (_10227_, _10226_, _10215_);
  or (_10228_, _10227_, _10208_);
  or (_10229_, _10228_, _03766_);
  and (_10230_, _10229_, _07914_);
  and (_10231_, _10230_, _10205_);
  and (_10232_, _07916_, _05247_);
  and (_10233_, _07927_, _07924_);
  nor (_10234_, _10233_, _07922_);
  not (_10235_, _10234_);
  and (_10236_, _08591_, _07924_);
  not (_10237_, _10236_);
  nor (_10238_, _10237_, _07979_);
  nor (_10239_, _10238_, _10235_);
  or (_10240_, _10239_, _10232_);
  and (_10241_, _10240_, _07913_);
  or (_10242_, _10241_, _07390_);
  or (_10243_, _10242_, _10231_);
  and (_10244_, _10243_, _09667_);
  or (_10245_, _10244_, _04481_);
  and (_10246_, _06069_, _05245_);
  or (_10247_, _09657_, _07400_);
  or (_10248_, _10247_, _10246_);
  and (_10249_, _10248_, _03589_);
  and (_10250_, _10249_, _10245_);
  or (_10251_, _10250_, _09664_);
  nor (_10252_, _07405_, _03585_);
  and (_10253_, _10252_, _10251_);
  nor (_10254_, _10162_, _07871_);
  and (_10255_, _10254_, _03585_);
  or (_10256_, _10255_, _03601_);
  or (_10257_, _10256_, _10253_);
  and (_10258_, _06171_, _05245_);
  or (_10259_, _10258_, _09657_);
  or (_10260_, _10259_, _05886_);
  and (_10261_, _10260_, _10257_);
  or (_10262_, _10261_, _03584_);
  not (_10263_, _03584_);
  nand (_10264_, _10162_, _07871_);
  or (_10265_, _10264_, _10263_);
  and (_10266_, _10265_, _10262_);
  or (_10267_, _10266_, _03600_);
  and (_10268_, _05884_, _05245_);
  or (_10269_, _10268_, _09657_);
  or (_10270_, _10269_, _07766_);
  and (_10271_, _10270_, _07778_);
  and (_10272_, _10271_, _10267_);
  or (_10273_, _10272_, _09660_);
  and (_10274_, _10273_, _07777_);
  or (_10275_, _09657_, _05310_);
  and (_10276_, _10259_, _03622_);
  and (_10277_, _10276_, _10275_);
  or (_10278_, _10277_, _10274_);
  and (_10279_, _10278_, _06828_);
  and (_10280_, _09884_, _03790_);
  and (_10281_, _10280_, _10275_);
  or (_10282_, _10281_, _03624_);
  or (_10283_, _10282_, _10279_);
  nor (_10284_, _05882_, _09661_);
  or (_10285_, _09657_, _07795_);
  or (_10286_, _10285_, _10284_);
  and (_10287_, _10286_, _07793_);
  and (_10288_, _10287_, _10283_);
  nor (_10289_, _06377_, _09661_);
  or (_10290_, _10289_, _09657_);
  and (_10291_, _10290_, _03785_);
  or (_10292_, _10291_, _08468_);
  or (_10293_, _10292_, _10288_);
  nor (_10294_, _07823_, _06075_);
  or (_10295_, _10294_, _07888_);
  or (_10296_, _10295_, _10176_);
  or (_10297_, _10296_, _07898_);
  and (_10298_, _10297_, _10293_);
  or (_10299_, _10298_, _08475_);
  nor (_10300_, _07989_, _06075_);
  or (_10301_, _10300_, _08500_);
  or (_10302_, _08477_, _10200_);
  or (_10303_, _10302_, _10301_);
  and (_10304_, _10303_, _03777_);
  and (_10305_, _10304_, _10299_);
  nor (_10306_, _08522_, _06075_);
  or (_10307_, _10306_, _08581_);
  or (_10308_, _10307_, _10208_);
  and (_10309_, _10308_, _03776_);
  or (_10310_, _10309_, _08506_);
  or (_10311_, _10310_, _10305_);
  nor (_10312_, _07921_, _06075_);
  or (_10313_, _10312_, _08611_);
  or (_10314_, _10232_, _08589_);
  or (_10315_, _10314_, _10313_);
  and (_10316_, _10315_, _08588_);
  and (_10317_, _10316_, _10311_);
  nor (_10318_, _08070_, _03949_);
  and (_10319_, _04474_, _03202_);
  nor (_10320_, _10319_, _10318_);
  nor (_10321_, _04488_, _04066_);
  or (_10322_, _10321_, _03949_);
  nand (_10323_, _10322_, _10320_);
  and (_10324_, _08587_, \oc8051_golden_model_1.ACC [7]);
  or (_10325_, _10324_, _10323_);
  or (_10326_, _10325_, _10317_);
  and (_10327_, _04058_, _03202_);
  not (_10328_, _10327_);
  nor (_10329_, _08662_, _08375_);
  not (_10330_, _10329_);
  or (_10331_, _10330_, _08692_);
  and (_10332_, _10331_, _08451_);
  and (_10333_, _10332_, _10328_);
  or (_10334_, _10333_, _08617_);
  and (_10335_, _10334_, _10326_);
  and (_10336_, _10332_, _10327_);
  or (_10337_, _10336_, _08620_);
  or (_10338_, _10337_, _10335_);
  and (_10339_, _08656_, _08400_);
  nor (_10340_, _08625_, _08399_);
  nor (_10341_, _10340_, _08398_);
  or (_10342_, _10341_, _08624_);
  or (_10343_, _10342_, _10339_);
  and (_10344_, _10343_, _08702_);
  and (_10345_, _10344_, _10338_);
  not (_10346_, _08406_);
  not (_10347_, _08405_);
  nand (_10348_, _08765_, _10347_);
  and (_10349_, _10348_, _08701_);
  and (_10350_, _10349_, _10346_);
  or (_10351_, _10350_, _03815_);
  not (_10352_, _08189_);
  nand (_10353_, _08725_, _10352_);
  and (_10354_, _10353_, _03517_);
  nor (_10355_, _08701_, _08188_);
  and (_10356_, _10355_, _10354_);
  or (_10357_, _10356_, _10351_);
  or (_10358_, _10357_, _10345_);
  not (_10359_, _08780_);
  or (_10360_, _09880_, _04246_);
  and (_10361_, _10360_, _10359_);
  and (_10362_, _10361_, _10358_);
  or (_10363_, _10362_, _09656_);
  and (_10364_, _10363_, _03823_);
  and (_10365_, _09914_, _03453_);
  or (_10366_, _10365_, _03447_);
  or (_10367_, _10366_, _10364_);
  and (_10368_, _05831_, _05245_);
  or (_10369_, _09657_, _03514_);
  or (_10370_, _10369_, _10368_);
  and (_10371_, _10370_, _10367_);
  or (_10372_, _10371_, _43004_);
  or (_10373_, _43000_, \oc8051_golden_model_1.PSW [7]);
  and (_10374_, _10373_, _41806_);
  and (_40578_, _10374_, _10372_);
  not (_10375_, \oc8051_golden_model_1.PCON [7]);
  nor (_10376_, _05212_, _10375_);
  not (_10377_, _05212_);
  nor (_10378_, _06377_, _10377_);
  nor (_10379_, _10378_, _10376_);
  nor (_10380_, _10379_, _07793_);
  and (_10381_, _06171_, _05212_);
  nor (_10382_, _10381_, _10376_);
  and (_10383_, _10382_, _03601_);
  nor (_10384_, _10377_, _05204_);
  nor (_10385_, _10384_, _10376_);
  and (_10386_, _10385_, _07390_);
  and (_10387_, _05212_, \oc8051_golden_model_1.ACC [7]);
  nor (_10388_, _10387_, _10376_);
  nor (_10389_, _10388_, _03737_);
  nor (_10390_, _10388_, _09029_);
  nor (_10391_, _04409_, _10375_);
  or (_10392_, _10391_, _10390_);
  and (_10393_, _10392_, _04081_);
  and (_10394_, _05964_, _05212_);
  nor (_10395_, _10394_, _10376_);
  nor (_10396_, _10395_, _04081_);
  or (_10397_, _10396_, _10393_);
  and (_10398_, _10397_, _03996_);
  nor (_10399_, _10385_, _03996_);
  nor (_10400_, _10399_, _10398_);
  nor (_10401_, _10400_, _03729_);
  or (_10402_, _10401_, _07390_);
  nor (_10403_, _10402_, _10389_);
  nor (_10404_, _10403_, _10386_);
  nor (_10405_, _10404_, _04481_);
  and (_10406_, _06069_, _05212_);
  nor (_10407_, _10376_, _07400_);
  not (_10408_, _10407_);
  nor (_10409_, _10408_, _10406_);
  or (_10410_, _10409_, _03222_);
  nor (_10411_, _10410_, _10405_);
  nor (_10412_, _06363_, _10377_);
  nor (_10413_, _10412_, _10376_);
  nor (_10414_, _10413_, _03589_);
  or (_10415_, _10414_, _03601_);
  nor (_10416_, _10415_, _10411_);
  nor (_10417_, _10416_, _10383_);
  or (_10418_, _10417_, _03600_);
  and (_10419_, _05884_, _05212_);
  or (_10420_, _10419_, _10376_);
  or (_10421_, _10420_, _07766_);
  and (_10422_, _10421_, _07778_);
  and (_10423_, _10422_, _10418_);
  and (_10424_, _06378_, _05212_);
  nor (_10425_, _10424_, _10376_);
  nor (_10426_, _10425_, _07778_);
  nor (_10427_, _10426_, _10423_);
  nor (_10428_, _10427_, _03622_);
  nor (_10429_, _10376_, _05310_);
  not (_10430_, _10429_);
  nor (_10431_, _10382_, _07777_);
  and (_10432_, _10431_, _10430_);
  nor (_10433_, _10432_, _10428_);
  nor (_10434_, _10433_, _03790_);
  nor (_10435_, _10388_, _06828_);
  and (_10436_, _10435_, _10430_);
  or (_10437_, _10436_, _10434_);
  and (_10438_, _10437_, _07795_);
  nor (_10439_, _05882_, _10377_);
  nor (_10440_, _10439_, _10376_);
  nor (_10441_, _10440_, _07795_);
  or (_10442_, _10441_, _10438_);
  and (_10443_, _10442_, _07793_);
  nor (_10444_, _10443_, _10380_);
  nor (_10445_, _10444_, _03815_);
  nor (_10446_, _10395_, _04246_);
  or (_10447_, _10446_, _03447_);
  nor (_10448_, _10447_, _10445_);
  and (_10449_, _05831_, _05212_);
  or (_10450_, _10376_, _03514_);
  nor (_10451_, _10450_, _10449_);
  nor (_10452_, _10451_, _10448_);
  or (_10453_, _10452_, _43004_);
  or (_10454_, _43000_, \oc8051_golden_model_1.PCON [7]);
  and (_10455_, _10454_, _41806_);
  and (_40579_, _10455_, _10453_);
  not (_10456_, \oc8051_golden_model_1.SBUF [7]);
  nor (_10457_, _05221_, _10456_);
  not (_10458_, _05221_);
  nor (_10459_, _06377_, _10458_);
  nor (_10460_, _10459_, _10457_);
  nor (_10461_, _10460_, _07793_);
  and (_10462_, _06171_, _05221_);
  nor (_10463_, _10462_, _10457_);
  and (_10464_, _10463_, _03601_);
  and (_10465_, _05221_, \oc8051_golden_model_1.ACC [7]);
  nor (_10466_, _10465_, _10457_);
  nor (_10467_, _10466_, _03737_);
  nor (_10468_, _10466_, _09029_);
  nor (_10469_, _04409_, _10456_);
  or (_10470_, _10469_, _10468_);
  and (_10471_, _10470_, _04081_);
  and (_10472_, _05964_, _05221_);
  nor (_10473_, _10472_, _10457_);
  nor (_10474_, _10473_, _04081_);
  or (_10475_, _10474_, _10471_);
  and (_10476_, _10475_, _03996_);
  nor (_10477_, _10458_, _05204_);
  nor (_10478_, _10477_, _10457_);
  nor (_10479_, _10478_, _03996_);
  nor (_10480_, _10479_, _10476_);
  nor (_10481_, _10480_, _03729_);
  or (_10482_, _10481_, _07390_);
  nor (_10483_, _10482_, _10467_);
  and (_10484_, _10478_, _07390_);
  nor (_10485_, _10484_, _10483_);
  nor (_10486_, _10485_, _04481_);
  and (_10487_, _06069_, _05221_);
  nor (_10488_, _10457_, _07400_);
  not (_10489_, _10488_);
  nor (_10490_, _10489_, _10487_);
  or (_10491_, _10490_, _03222_);
  nor (_10492_, _10491_, _10486_);
  nor (_10493_, _06363_, _10458_);
  nor (_10494_, _10493_, _10457_);
  nor (_10495_, _10494_, _03589_);
  or (_10496_, _10495_, _03601_);
  nor (_10497_, _10496_, _10492_);
  nor (_10498_, _10497_, _10464_);
  or (_10499_, _10498_, _03600_);
  and (_10500_, _05884_, _05221_);
  or (_10501_, _10500_, _10457_);
  or (_10502_, _10501_, _07766_);
  and (_10503_, _10502_, _07778_);
  and (_10504_, _10503_, _10499_);
  and (_10505_, _06378_, _05221_);
  nor (_10506_, _10505_, _10457_);
  nor (_10507_, _10506_, _07778_);
  nor (_10508_, _10507_, _10504_);
  nor (_10509_, _10508_, _03622_);
  nor (_10510_, _10457_, _05310_);
  not (_10511_, _10510_);
  nor (_10512_, _10463_, _07777_);
  and (_10513_, _10512_, _10511_);
  nor (_10514_, _10513_, _10509_);
  nor (_10515_, _10514_, _03790_);
  nor (_10516_, _10466_, _06828_);
  and (_10517_, _10516_, _10511_);
  or (_10518_, _10517_, _10515_);
  and (_10519_, _10518_, _07795_);
  nor (_10520_, _05882_, _10458_);
  nor (_10521_, _10520_, _10457_);
  nor (_10522_, _10521_, _07795_);
  or (_10523_, _10522_, _10519_);
  and (_10524_, _10523_, _07793_);
  nor (_10525_, _10524_, _10461_);
  nor (_10526_, _10525_, _03815_);
  nor (_10527_, _10473_, _04246_);
  or (_10528_, _10527_, _03447_);
  nor (_10529_, _10528_, _10526_);
  and (_10530_, _05831_, _05221_);
  or (_10531_, _10457_, _03514_);
  nor (_10532_, _10531_, _10530_);
  nor (_10533_, _10532_, _10529_);
  or (_10534_, _10533_, _43004_);
  or (_10535_, _43000_, \oc8051_golden_model_1.SBUF [7]);
  and (_10536_, _10535_, _41806_);
  and (_40580_, _10536_, _10534_);
  not (_10537_, \oc8051_golden_model_1.SCON [7]);
  nor (_10538_, _05275_, _10537_);
  not (_10539_, _05275_);
  nor (_10540_, _10539_, _05204_);
  nor (_10541_, _10540_, _10538_);
  and (_10542_, _10541_, _07390_);
  nor (_10543_, _05922_, _10537_);
  and (_10544_, _05952_, _05922_);
  nor (_10545_, _10544_, _10543_);
  nor (_10546_, _10545_, _03736_);
  and (_10547_, _05275_, \oc8051_golden_model_1.ACC [7]);
  nor (_10548_, _10547_, _10538_);
  nor (_10549_, _10548_, _09029_);
  nor (_10550_, _04409_, _10537_);
  or (_10551_, _10550_, _10549_);
  and (_10552_, _10551_, _04081_);
  and (_10553_, _05964_, _05275_);
  nor (_10554_, _10553_, _10538_);
  nor (_10555_, _10554_, _04081_);
  or (_10556_, _10555_, _10552_);
  and (_10557_, _10556_, _04055_);
  and (_10558_, _06095_, _05922_);
  nor (_10559_, _10558_, _10543_);
  nor (_10560_, _10559_, _04055_);
  or (_10561_, _10560_, _03723_);
  or (_10562_, _10561_, _10557_);
  nand (_10563_, _10541_, _03723_);
  and (_10564_, _10563_, _10562_);
  and (_10565_, _10564_, _03737_);
  nor (_10566_, _10548_, _03737_);
  or (_10567_, _10566_, _10565_);
  and (_10568_, _10567_, _03736_);
  nor (_10569_, _10568_, _10546_);
  nor (_10570_, _10569_, _03719_);
  nor (_10571_, _10543_, _06138_);
  or (_10572_, _10559_, _06840_);
  nor (_10573_, _10572_, _10571_);
  nor (_10574_, _10573_, _10570_);
  nor (_10575_, _10574_, _03505_);
  not (_10576_, _05922_);
  nor (_10577_, _05938_, _10576_);
  nor (_10578_, _10577_, _10543_);
  nor (_10579_, _10578_, _03710_);
  nor (_10580_, _10579_, _07390_);
  not (_10581_, _10580_);
  nor (_10582_, _10581_, _10575_);
  nor (_10583_, _10582_, _10542_);
  nor (_10584_, _10583_, _04481_);
  and (_10585_, _06069_, _05275_);
  nor (_10586_, _10538_, _07400_);
  not (_10587_, _10586_);
  nor (_10588_, _10587_, _10585_);
  nor (_10589_, _10588_, _03222_);
  not (_10590_, _10589_);
  nor (_10591_, _10590_, _10584_);
  nor (_10592_, _06363_, _10539_);
  nor (_10593_, _10592_, _10538_);
  nor (_10594_, _10593_, _03589_);
  or (_10595_, _10594_, _08828_);
  or (_10596_, _10595_, _10591_);
  and (_10597_, _05884_, _05275_);
  or (_10598_, _10538_, _07766_);
  or (_10599_, _10598_, _10597_);
  and (_10600_, _06171_, _05275_);
  nor (_10601_, _10600_, _10538_);
  and (_10602_, _10601_, _03601_);
  nor (_10603_, _10602_, _03780_);
  and (_10604_, _10603_, _10599_);
  and (_10605_, _10604_, _10596_);
  and (_10606_, _06378_, _05275_);
  nor (_10607_, _10606_, _10538_);
  nor (_10608_, _10607_, _07778_);
  nor (_10609_, _10608_, _10605_);
  nor (_10610_, _10609_, _03622_);
  nor (_10611_, _10538_, _05310_);
  not (_10612_, _10611_);
  nor (_10613_, _10601_, _07777_);
  and (_10614_, _10613_, _10612_);
  nor (_10615_, _10614_, _10610_);
  nor (_10616_, _10615_, _03790_);
  nor (_10617_, _10548_, _06828_);
  and (_10618_, _10617_, _10612_);
  nor (_10619_, _10618_, _03624_);
  not (_10620_, _10619_);
  nor (_10621_, _10620_, _10616_);
  nor (_10622_, _05882_, _10539_);
  or (_10623_, _10538_, _07795_);
  nor (_10624_, _10623_, _10622_);
  or (_10625_, _10624_, _03785_);
  nor (_10626_, _10625_, _10621_);
  nor (_10627_, _06377_, _10539_);
  nor (_10628_, _10627_, _10538_);
  nor (_10629_, _10628_, _07793_);
  or (_10630_, _10629_, _10626_);
  and (_10631_, _10630_, _04246_);
  nor (_10632_, _10554_, _04246_);
  or (_10633_, _10632_, _10631_);
  and (_10634_, _10633_, _03823_);
  nor (_10635_, _10545_, _03823_);
  or (_10636_, _10635_, _10634_);
  and (_10637_, _10636_, _03514_);
  and (_10638_, _05831_, _05275_);
  nor (_10639_, _10638_, _10538_);
  nor (_10640_, _10639_, _03514_);
  or (_10641_, _10640_, _10637_);
  or (_10642_, _10641_, _43004_);
  or (_10643_, _43000_, \oc8051_golden_model_1.SCON [7]);
  and (_10644_, _10643_, _41806_);
  and (_40581_, _10644_, _10642_);
  and (_10645_, _05010_, \oc8051_golden_model_1.SP [4]);
  and (_10646_, _10645_, \oc8051_golden_model_1.SP [5]);
  and (_10647_, _10646_, \oc8051_golden_model_1.SP [6]);
  nor (_10648_, _10647_, \oc8051_golden_model_1.SP [7]);
  and (_10649_, _10647_, \oc8051_golden_model_1.SP [7]);
  nor (_10650_, _10649_, _10648_);
  nor (_10651_, _10650_, _04540_);
  not (_10652_, _03798_);
  not (_10653_, \oc8051_golden_model_1.SP [7]);
  nor (_10654_, _05300_, _10653_);
  and (_10655_, _06378_, _05300_);
  nor (_10656_, _10655_, _10654_);
  nor (_10657_, _10656_, _07778_);
  not (_10658_, _06837_);
  nor (_10659_, _10650_, _04767_);
  nor (_10660_, _04409_, _10653_);
  and (_10661_, _05300_, \oc8051_golden_model_1.ACC [7]);
  nor (_10662_, _10661_, _10654_);
  nor (_10663_, _10662_, _09029_);
  or (_10664_, _10663_, _10660_);
  and (_10665_, _10664_, _04763_);
  and (_10666_, _10650_, _03980_);
  nor (_10667_, _10666_, _10665_);
  nor (_10668_, _10667_, _03610_);
  and (_10669_, _05964_, _05300_);
  nor (_10670_, _10669_, _10654_);
  nor (_10671_, _10670_, _04081_);
  or (_10672_, _10671_, _10668_);
  and (_10673_, _10672_, _03230_);
  and (_10674_, _10650_, _04768_);
  or (_10675_, _10674_, _10673_);
  and (_10676_, _10675_, _03996_);
  not (_10677_, \oc8051_golden_model_1.SP [6]);
  not (_10678_, \oc8051_golden_model_1.SP [5]);
  not (_10679_, \oc8051_golden_model_1.SP [4]);
  and (_10680_, _05971_, _10679_);
  and (_10681_, _10680_, _10678_);
  and (_10682_, _10681_, _10677_);
  and (_10683_, _10682_, _03498_);
  nor (_10684_, _10683_, _10653_);
  and (_10685_, _10683_, _10653_);
  nor (_10686_, _10685_, _10684_);
  nor (_10687_, _10686_, _03996_);
  or (_10688_, _10687_, _10676_);
  and (_10689_, _10688_, _03737_);
  nor (_10691_, _10662_, _03737_);
  or (_10692_, _10691_, _10689_);
  and (_10693_, _10692_, _03510_);
  not (_10694_, _04767_);
  and (_10695_, _10647_, \oc8051_golden_model_1.SP [0]);
  nor (_10696_, _10695_, _10653_);
  and (_10697_, _10695_, _10653_);
  nor (_10698_, _10697_, _10696_);
  nor (_10699_, _10698_, _03510_);
  nor (_10700_, _10699_, _10694_);
  not (_10702_, _10700_);
  nor (_10703_, _10702_, _10693_);
  nor (_10704_, _10703_, _10659_);
  nor (_10705_, _10704_, _10658_);
  not (_10706_, _05300_);
  nor (_10707_, _10706_, _05204_);
  nor (_10708_, _10707_, _10654_);
  and (_10709_, _10708_, _10658_);
  nor (_10710_, _10709_, _06833_);
  not (_10711_, _10710_);
  nor (_10713_, _10711_, _10705_);
  nor (_10714_, _10708_, _06834_);
  nor (_10715_, _10714_, _04481_);
  not (_10716_, _10715_);
  nor (_10717_, _10716_, _10713_);
  and (_10718_, _06069_, _05300_);
  nor (_10719_, _10654_, _07400_);
  not (_10720_, _10719_);
  nor (_10721_, _10720_, _10718_);
  nor (_10722_, _10721_, _10717_);
  nor (_10724_, _10722_, _03222_);
  nor (_10725_, _06363_, _10706_);
  or (_10726_, _10654_, _03589_);
  nor (_10727_, _10726_, _10725_);
  or (_10728_, _10727_, _03601_);
  nor (_10729_, _10728_, _10724_);
  and (_10730_, _06171_, _05300_);
  nor (_10731_, _10730_, _10654_);
  nor (_10732_, _10731_, _05886_);
  or (_10733_, _10732_, _03178_);
  or (_10735_, _10733_, _10729_);
  not (_10736_, _03178_);
  or (_10737_, _10650_, _10736_);
  and (_10738_, _10737_, _10735_);
  nor (_10739_, _10738_, _03600_);
  and (_10740_, _05884_, _05300_);
  or (_10741_, _10654_, _07766_);
  nor (_10742_, _10741_, _10740_);
  or (_10743_, _10742_, _03780_);
  nor (_10744_, _10743_, _10739_);
  nor (_10746_, _10744_, _10657_);
  nor (_10747_, _10746_, _03622_);
  nor (_10748_, _10654_, _05310_);
  not (_10749_, _10748_);
  nor (_10750_, _10731_, _07777_);
  and (_10751_, _10750_, _10749_);
  nor (_10752_, _10751_, _10747_);
  nor (_10753_, _03790_, _03192_);
  not (_10754_, _10753_);
  nor (_10755_, _10754_, _10752_);
  and (_10757_, _10650_, _03192_);
  or (_10758_, _10748_, _06828_);
  nor (_10759_, _10758_, _10662_);
  nor (_10760_, _10759_, _10757_);
  and (_10761_, _10760_, _07795_);
  not (_10762_, _10761_);
  nor (_10763_, _10762_, _10755_);
  nor (_10764_, _05882_, _10706_);
  nor (_10765_, _10764_, _10654_);
  and (_10766_, _10765_, _03624_);
  nor (_10767_, _10766_, _10763_);
  and (_10768_, _10767_, _07793_);
  nor (_10769_, _06377_, _10706_);
  nor (_10770_, _10769_, _10654_);
  nor (_10771_, _10770_, _07793_);
  or (_10772_, _10771_, _10768_);
  and (_10773_, _10772_, _10652_);
  nor (_10774_, _03798_, _03188_);
  nor (_10775_, _10682_, \oc8051_golden_model_1.SP [7]);
  and (_10776_, _10682_, \oc8051_golden_model_1.SP [7]);
  nor (_10777_, _10776_, _10775_);
  nor (_10778_, _10777_, _03188_);
  nor (_10779_, _10778_, _10774_);
  nor (_10780_, _10779_, _10773_);
  nor (_10781_, _10650_, _06399_);
  nor (_10782_, _10781_, _10780_);
  and (_10783_, _10782_, _03516_);
  and (_10784_, _10777_, _03515_);
  or (_10785_, _10784_, _10783_);
  and (_10786_, _10785_, _04246_);
  nor (_10787_, _10670_, _04246_);
  nor (_10788_, _10787_, _05103_);
  not (_10789_, _10788_);
  nor (_10790_, _10789_, _10786_);
  nor (_10791_, _10790_, _10651_);
  and (_10792_, _10791_, _03514_);
  and (_10793_, _05831_, _05300_);
  nor (_10794_, _10793_, _10654_);
  nor (_10795_, _10794_, _03514_);
  or (_10796_, _10795_, _10792_);
  or (_10797_, _10796_, _43004_);
  or (_10798_, _43000_, \oc8051_golden_model_1.SP [7]);
  and (_10799_, _10798_, _41806_);
  and (_40583_, _10799_, _10797_);
  not (_10800_, \oc8051_golden_model_1.TCON [7]);
  nor (_10801_, _05258_, _10800_);
  not (_10802_, _05258_);
  nor (_10803_, _10802_, _05204_);
  nor (_10804_, _10803_, _10801_);
  and (_10805_, _10804_, _07390_);
  nor (_10806_, _05927_, _10800_);
  and (_10807_, _05952_, _05927_);
  nor (_10808_, _10807_, _10806_);
  nor (_10809_, _10808_, _03736_);
  and (_10810_, _05258_, \oc8051_golden_model_1.ACC [7]);
  nor (_10811_, _10810_, _10801_);
  nor (_10812_, _10811_, _09029_);
  nor (_10813_, _04409_, _10800_);
  or (_10814_, _10813_, _10812_);
  and (_10815_, _10814_, _04081_);
  and (_10816_, _05964_, _05258_);
  nor (_10817_, _10816_, _10801_);
  nor (_10818_, _10817_, _04081_);
  or (_10819_, _10818_, _10815_);
  and (_10820_, _10819_, _04055_);
  and (_10821_, _06095_, _05927_);
  nor (_10822_, _10821_, _10806_);
  nor (_10823_, _10822_, _04055_);
  or (_10824_, _10823_, _03723_);
  or (_10825_, _10824_, _10820_);
  nand (_10826_, _10804_, _03723_);
  and (_10827_, _10826_, _10825_);
  and (_10828_, _10827_, _03737_);
  nor (_10829_, _10811_, _03737_);
  or (_10830_, _10829_, _10828_);
  and (_10831_, _10830_, _03736_);
  nor (_10832_, _10831_, _10809_);
  nor (_10833_, _10832_, _03719_);
  and (_10834_, _06139_, _05927_);
  nor (_10835_, _10834_, _10806_);
  nor (_10836_, _10835_, _06840_);
  nor (_10837_, _10836_, _10833_);
  nor (_10838_, _10837_, _03505_);
  not (_10839_, _05927_);
  nor (_10840_, _05938_, _10839_);
  nor (_10841_, _10840_, _10806_);
  nor (_10842_, _10841_, _03710_);
  nor (_10843_, _10842_, _07390_);
  not (_10844_, _10843_);
  nor (_10845_, _10844_, _10838_);
  nor (_10846_, _10845_, _10805_);
  nor (_10847_, _10846_, _04481_);
  and (_10848_, _06069_, _05258_);
  nor (_10849_, _10801_, _07400_);
  not (_10850_, _10849_);
  nor (_10851_, _10850_, _10848_);
  nor (_10852_, _10851_, _03222_);
  not (_10853_, _10852_);
  nor (_10854_, _10853_, _10847_);
  nor (_10855_, _06363_, _10802_);
  nor (_10856_, _10855_, _10801_);
  nor (_10857_, _10856_, _03589_);
  or (_10858_, _10857_, _08828_);
  or (_10859_, _10858_, _10854_);
  and (_10860_, _05884_, _05258_);
  or (_10861_, _10801_, _07766_);
  or (_10862_, _10861_, _10860_);
  and (_10863_, _06171_, _05258_);
  nor (_10864_, _10863_, _10801_);
  and (_10865_, _10864_, _03601_);
  nor (_10866_, _10865_, _03780_);
  and (_10867_, _10866_, _10862_);
  and (_10868_, _10867_, _10859_);
  and (_10869_, _06378_, _05258_);
  nor (_10870_, _10869_, _10801_);
  nor (_10871_, _10870_, _07778_);
  nor (_10872_, _10871_, _10868_);
  nor (_10873_, _10872_, _03622_);
  nor (_10874_, _10801_, _05310_);
  not (_10875_, _10874_);
  nor (_10876_, _10864_, _07777_);
  and (_10877_, _10876_, _10875_);
  nor (_10878_, _10877_, _10873_);
  nor (_10879_, _10878_, _03790_);
  nor (_10880_, _10811_, _06828_);
  and (_10881_, _10880_, _10875_);
  or (_10882_, _10881_, _10879_);
  and (_10883_, _10882_, _07795_);
  nor (_10884_, _05882_, _10802_);
  nor (_10885_, _10884_, _10801_);
  nor (_10886_, _10885_, _07795_);
  or (_10887_, _10886_, _10883_);
  and (_10888_, _10887_, _07793_);
  nor (_10889_, _06377_, _10802_);
  nor (_10890_, _10889_, _10801_);
  nor (_10891_, _10890_, _07793_);
  or (_10892_, _10891_, _10888_);
  and (_10893_, _10892_, _04246_);
  nor (_10894_, _10817_, _04246_);
  or (_10895_, _10894_, _10893_);
  and (_10896_, _10895_, _03823_);
  nor (_10897_, _10808_, _03823_);
  or (_10898_, _10897_, _10896_);
  and (_10899_, _10898_, _03514_);
  and (_10900_, _05831_, _05258_);
  nor (_10901_, _10900_, _10801_);
  nor (_10902_, _10901_, _03514_);
  or (_10903_, _10902_, _10899_);
  or (_10904_, _10903_, _43004_);
  or (_10905_, _43000_, \oc8051_golden_model_1.TCON [7]);
  and (_10906_, _10905_, _41806_);
  and (_40584_, _10906_, _10904_);
  not (_10907_, \oc8051_golden_model_1.TH0 [7]);
  nor (_10908_, _05263_, _10907_);
  not (_10909_, _05263_);
  nor (_10910_, _06377_, _10909_);
  nor (_10911_, _10910_, _10908_);
  nor (_10912_, _10911_, _07793_);
  and (_10913_, _06171_, _05263_);
  nor (_10914_, _10913_, _10908_);
  and (_10915_, _10914_, _03601_);
  nor (_10916_, _10909_, _05204_);
  nor (_10917_, _10916_, _10908_);
  and (_10918_, _10917_, _07390_);
  and (_10919_, _05263_, \oc8051_golden_model_1.ACC [7]);
  nor (_10920_, _10919_, _10908_);
  nor (_10921_, _10920_, _03737_);
  nor (_10922_, _10920_, _09029_);
  nor (_10923_, _04409_, _10907_);
  or (_10924_, _10923_, _10922_);
  and (_10925_, _10924_, _04081_);
  and (_10926_, _05964_, _05263_);
  nor (_10927_, _10926_, _10908_);
  nor (_10928_, _10927_, _04081_);
  or (_10929_, _10928_, _10925_);
  and (_10930_, _10929_, _03996_);
  nor (_10931_, _10917_, _03996_);
  nor (_10932_, _10931_, _10930_);
  nor (_10933_, _10932_, _03729_);
  or (_10934_, _10933_, _07390_);
  nor (_10935_, _10934_, _10921_);
  nor (_10936_, _10935_, _10918_);
  nor (_10937_, _10936_, _04481_);
  and (_10938_, _06069_, _05263_);
  nor (_10939_, _10908_, _07400_);
  not (_10940_, _10939_);
  nor (_10941_, _10940_, _10938_);
  or (_10942_, _10941_, _03222_);
  nor (_10943_, _10942_, _10937_);
  nor (_10944_, _06363_, _10909_);
  nor (_10945_, _10944_, _10908_);
  nor (_10946_, _10945_, _03589_);
  or (_10947_, _10946_, _03601_);
  nor (_10948_, _10947_, _10943_);
  nor (_10949_, _10948_, _10915_);
  or (_10950_, _10949_, _03600_);
  and (_10951_, _05884_, _05263_);
  or (_10952_, _10951_, _10908_);
  or (_10953_, _10952_, _07766_);
  and (_10954_, _10953_, _07778_);
  and (_10955_, _10954_, _10950_);
  and (_10956_, _06378_, _05263_);
  nor (_10957_, _10956_, _10908_);
  nor (_10958_, _10957_, _07778_);
  nor (_10959_, _10958_, _10955_);
  nor (_10960_, _10959_, _03622_);
  nor (_10961_, _10908_, _05310_);
  not (_10962_, _10961_);
  nor (_10963_, _10914_, _07777_);
  and (_10964_, _10963_, _10962_);
  nor (_10965_, _10964_, _10960_);
  nor (_10966_, _10965_, _03790_);
  nor (_10967_, _10920_, _06828_);
  and (_10968_, _10967_, _10962_);
  nor (_10969_, _10968_, _03624_);
  not (_10970_, _10969_);
  nor (_10971_, _10970_, _10966_);
  nor (_10972_, _05882_, _10909_);
  or (_10973_, _10908_, _07795_);
  nor (_10974_, _10973_, _10972_);
  or (_10975_, _10974_, _03785_);
  nor (_10976_, _10975_, _10971_);
  nor (_10977_, _10976_, _10912_);
  nor (_10978_, _10977_, _03815_);
  nor (_10979_, _10927_, _04246_);
  or (_10980_, _10979_, _03447_);
  nor (_10981_, _10980_, _10978_);
  and (_10982_, _05831_, _05263_);
  or (_10983_, _10908_, _03514_);
  nor (_10984_, _10983_, _10982_);
  nor (_10985_, _10984_, _10981_);
  or (_10986_, _10985_, _43004_);
  or (_10987_, _43000_, \oc8051_golden_model_1.TH0 [7]);
  and (_10988_, _10987_, _41806_);
  and (_40585_, _10988_, _10986_);
  not (_10989_, \oc8051_golden_model_1.TH1 [7]);
  nor (_10990_, _05278_, _10989_);
  not (_10991_, _05278_);
  nor (_10992_, _06377_, _10991_);
  nor (_10993_, _10992_, _10990_);
  nor (_10994_, _10993_, _07793_);
  and (_10995_, _06171_, _05278_);
  nor (_10996_, _10995_, _10990_);
  and (_10997_, _10996_, _03601_);
  and (_10998_, _05278_, \oc8051_golden_model_1.ACC [7]);
  nor (_10999_, _10998_, _10990_);
  nor (_11000_, _10999_, _03737_);
  nor (_11001_, _10999_, _09029_);
  nor (_11002_, _04409_, _10989_);
  or (_11003_, _11002_, _11001_);
  and (_11004_, _11003_, _04081_);
  and (_11005_, _05964_, _05278_);
  nor (_11006_, _11005_, _10990_);
  nor (_11007_, _11006_, _04081_);
  or (_11008_, _11007_, _11004_);
  and (_11009_, _11008_, _03996_);
  nor (_11010_, _10991_, _05204_);
  nor (_11011_, _11010_, _10990_);
  nor (_11012_, _11011_, _03996_);
  nor (_11013_, _11012_, _11009_);
  nor (_11014_, _11013_, _03729_);
  or (_11015_, _11014_, _07390_);
  nor (_11016_, _11015_, _11000_);
  and (_11017_, _11011_, _07390_);
  nor (_11018_, _11017_, _11016_);
  nor (_11019_, _11018_, _04481_);
  and (_11020_, _06069_, _05278_);
  nor (_11021_, _10990_, _07400_);
  not (_11022_, _11021_);
  nor (_11023_, _11022_, _11020_);
  or (_11024_, _11023_, _03222_);
  nor (_11025_, _11024_, _11019_);
  nor (_11026_, _06363_, _10991_);
  nor (_11027_, _11026_, _10990_);
  nor (_11028_, _11027_, _03589_);
  or (_11029_, _11028_, _03601_);
  nor (_11030_, _11029_, _11025_);
  nor (_11031_, _11030_, _10997_);
  or (_11032_, _11031_, _03600_);
  and (_11033_, _05884_, _05278_);
  or (_11034_, _11033_, _10990_);
  or (_11035_, _11034_, _07766_);
  and (_11036_, _11035_, _07778_);
  and (_11037_, _11036_, _11032_);
  and (_11038_, _06378_, _05278_);
  nor (_11039_, _11038_, _10990_);
  nor (_11040_, _11039_, _07778_);
  nor (_11041_, _11040_, _11037_);
  nor (_11042_, _11041_, _03622_);
  nor (_11043_, _10990_, _05310_);
  not (_11044_, _11043_);
  nor (_11045_, _10996_, _07777_);
  and (_11046_, _11045_, _11044_);
  nor (_11047_, _11046_, _11042_);
  nor (_11048_, _11047_, _03790_);
  nor (_11049_, _10999_, _06828_);
  and (_11050_, _11049_, _11044_);
  or (_11051_, _11050_, _11048_);
  and (_11052_, _11051_, _07795_);
  nor (_11053_, _05882_, _10991_);
  nor (_11054_, _11053_, _10990_);
  nor (_11055_, _11054_, _07795_);
  or (_11056_, _11055_, _11052_);
  and (_11057_, _11056_, _07793_);
  nor (_11058_, _11057_, _10994_);
  nor (_11059_, _11058_, _03815_);
  nor (_11060_, _11006_, _04246_);
  or (_11061_, _11060_, _03447_);
  nor (_11062_, _11061_, _11059_);
  and (_11063_, _05831_, _05278_);
  or (_11064_, _10990_, _03514_);
  nor (_11065_, _11064_, _11063_);
  nor (_11066_, _11065_, _11062_);
  or (_11067_, _11066_, _43004_);
  or (_11068_, _43000_, \oc8051_golden_model_1.TH1 [7]);
  and (_11069_, _11068_, _41806_);
  and (_40586_, _11069_, _11067_);
  not (_11070_, \oc8051_golden_model_1.TL0 [7]);
  nor (_11071_, _05284_, _11070_);
  not (_11072_, _05284_);
  nor (_11073_, _06377_, _11072_);
  nor (_11074_, _11073_, _11071_);
  nor (_11075_, _11074_, _07793_);
  and (_11076_, _06171_, _05284_);
  nor (_11077_, _11076_, _11071_);
  and (_11078_, _11077_, _03601_);
  and (_11079_, _05284_, \oc8051_golden_model_1.ACC [7]);
  nor (_11080_, _11079_, _11071_);
  nor (_11081_, _11080_, _03737_);
  nor (_11082_, _11080_, _09029_);
  nor (_11083_, _04409_, _11070_);
  or (_11084_, _11083_, _11082_);
  and (_11085_, _11084_, _04081_);
  and (_11086_, _05964_, _05284_);
  nor (_11087_, _11086_, _11071_);
  nor (_11088_, _11087_, _04081_);
  or (_11089_, _11088_, _11085_);
  and (_11090_, _11089_, _03996_);
  nor (_11091_, _11072_, _05204_);
  nor (_11092_, _11091_, _11071_);
  nor (_11093_, _11092_, _03996_);
  nor (_11094_, _11093_, _11090_);
  nor (_11095_, _11094_, _03729_);
  or (_11096_, _11095_, _07390_);
  nor (_11097_, _11096_, _11081_);
  and (_11098_, _11092_, _07390_);
  nor (_11099_, _11098_, _11097_);
  nor (_11100_, _11099_, _04481_);
  and (_11101_, _06069_, _05284_);
  nor (_11102_, _11071_, _07400_);
  not (_11103_, _11102_);
  nor (_11104_, _11103_, _11101_);
  or (_11105_, _11104_, _03222_);
  nor (_11106_, _11105_, _11100_);
  nor (_11107_, _06363_, _11072_);
  nor (_11108_, _11107_, _11071_);
  nor (_11109_, _11108_, _03589_);
  or (_11110_, _11109_, _03601_);
  nor (_11111_, _11110_, _11106_);
  nor (_11112_, _11111_, _11078_);
  or (_11113_, _11112_, _03600_);
  and (_11114_, _05884_, _05284_);
  or (_11115_, _11114_, _11071_);
  or (_11116_, _11115_, _07766_);
  and (_11117_, _11116_, _07778_);
  and (_11118_, _11117_, _11113_);
  and (_11119_, _06378_, _05284_);
  nor (_11120_, _11119_, _11071_);
  nor (_11121_, _11120_, _07778_);
  nor (_11122_, _11121_, _11118_);
  nor (_11123_, _11122_, _03622_);
  nor (_11124_, _11071_, _05310_);
  not (_11125_, _11124_);
  nor (_11126_, _11077_, _07777_);
  and (_11127_, _11126_, _11125_);
  nor (_11128_, _11127_, _11123_);
  nor (_11129_, _11128_, _03790_);
  nor (_11130_, _11080_, _06828_);
  and (_11131_, _11130_, _11125_);
  nor (_11132_, _11131_, _03624_);
  not (_11133_, _11132_);
  nor (_11134_, _11133_, _11129_);
  nor (_11135_, _05882_, _11072_);
  or (_11136_, _11071_, _07795_);
  nor (_11137_, _11136_, _11135_);
  or (_11138_, _11137_, _03785_);
  nor (_11139_, _11138_, _11134_);
  nor (_11140_, _11139_, _11075_);
  nor (_11141_, _11140_, _03815_);
  nor (_11142_, _11087_, _04246_);
  or (_11143_, _11142_, _03447_);
  nor (_11144_, _11143_, _11141_);
  and (_11145_, _05831_, _05284_);
  nor (_11146_, _11145_, _11071_);
  and (_11147_, _11146_, _03447_);
  nor (_11148_, _11147_, _11144_);
  or (_11149_, _11148_, _43004_);
  or (_11150_, _43000_, \oc8051_golden_model_1.TL0 [7]);
  and (_11151_, _11150_, _41806_);
  and (_40587_, _11151_, _11149_);
  not (_11152_, \oc8051_golden_model_1.TL1 [7]);
  nor (_11153_, _05271_, _11152_);
  not (_11154_, _05271_);
  nor (_11155_, _06377_, _11154_);
  nor (_11156_, _11155_, _11153_);
  nor (_11157_, _11156_, _07793_);
  and (_11158_, _06171_, _05271_);
  nor (_11159_, _11158_, _11153_);
  and (_11160_, _11159_, _03601_);
  and (_11161_, _05271_, \oc8051_golden_model_1.ACC [7]);
  nor (_11162_, _11161_, _11153_);
  nor (_11163_, _11162_, _03737_);
  nor (_11164_, _11162_, _09029_);
  nor (_11165_, _04409_, _11152_);
  or (_11166_, _11165_, _11164_);
  and (_11167_, _11166_, _04081_);
  and (_11168_, _05964_, _05271_);
  nor (_11169_, _11168_, _11153_);
  nor (_11170_, _11169_, _04081_);
  or (_11171_, _11170_, _11167_);
  and (_11172_, _11171_, _03996_);
  nor (_11173_, _11154_, _05204_);
  nor (_11174_, _11173_, _11153_);
  nor (_11175_, _11174_, _03996_);
  nor (_11176_, _11175_, _11172_);
  nor (_11177_, _11176_, _03729_);
  or (_11178_, _11177_, _07390_);
  nor (_11179_, _11178_, _11163_);
  and (_11180_, _11174_, _07390_);
  nor (_11181_, _11180_, _11179_);
  nor (_11182_, _11181_, _04481_);
  and (_11183_, _06069_, _05271_);
  nor (_11184_, _11153_, _07400_);
  not (_11185_, _11184_);
  nor (_11186_, _11185_, _11183_);
  or (_11187_, _11186_, _03222_);
  nor (_11188_, _11187_, _11182_);
  nor (_11189_, _06363_, _11154_);
  nor (_11190_, _11189_, _11153_);
  nor (_11191_, _11190_, _03589_);
  or (_11192_, _11191_, _03601_);
  nor (_11193_, _11192_, _11188_);
  nor (_11194_, _11193_, _11160_);
  or (_11195_, _11194_, _03600_);
  and (_11196_, _05884_, _05271_);
  or (_11197_, _11196_, _11153_);
  or (_11198_, _11197_, _07766_);
  and (_11199_, _11198_, _07778_);
  and (_11200_, _11199_, _11195_);
  and (_11201_, _06378_, _05271_);
  nor (_11202_, _11201_, _11153_);
  nor (_11203_, _11202_, _07778_);
  nor (_11204_, _11203_, _11200_);
  nor (_11205_, _11204_, _03622_);
  nor (_11206_, _11153_, _05310_);
  not (_11207_, _11206_);
  nor (_11208_, _11159_, _07777_);
  and (_11209_, _11208_, _11207_);
  nor (_11210_, _11209_, _11205_);
  nor (_11211_, _11210_, _03790_);
  nor (_11212_, _11162_, _06828_);
  and (_11213_, _11212_, _11207_);
  nor (_11214_, _11213_, _03624_);
  not (_11215_, _11214_);
  nor (_11216_, _11215_, _11211_);
  nor (_11217_, _05882_, _11154_);
  or (_11218_, _11153_, _07795_);
  nor (_11219_, _11218_, _11217_);
  or (_11220_, _11219_, _03785_);
  nor (_11221_, _11220_, _11216_);
  nor (_11222_, _11221_, _11157_);
  nor (_11223_, _11222_, _03815_);
  nor (_11224_, _11169_, _04246_);
  or (_11225_, _11224_, _03447_);
  nor (_11226_, _11225_, _11223_);
  and (_11227_, _05831_, _05271_);
  or (_11228_, _11153_, _03514_);
  nor (_11229_, _11228_, _11227_);
  nor (_11230_, _11229_, _11226_);
  or (_11231_, _11230_, _43004_);
  or (_11232_, _43000_, \oc8051_golden_model_1.TL1 [7]);
  and (_11233_, _11232_, _41806_);
  and (_40589_, _11233_, _11231_);
  not (_11234_, \oc8051_golden_model_1.TMOD [7]);
  nor (_11235_, _05286_, _11234_);
  not (_11236_, _05286_);
  nor (_11237_, _06377_, _11236_);
  nor (_11238_, _11237_, _11235_);
  nor (_11239_, _11238_, _07793_);
  and (_11240_, _06171_, _05286_);
  nor (_11241_, _11240_, _11235_);
  and (_11242_, _11241_, _03601_);
  and (_11243_, _05286_, \oc8051_golden_model_1.ACC [7]);
  nor (_11244_, _11243_, _11235_);
  nor (_11245_, _11244_, _03737_);
  nor (_11246_, _11244_, _09029_);
  nor (_11247_, _04409_, _11234_);
  or (_11248_, _11247_, _11246_);
  and (_11249_, _11248_, _04081_);
  and (_11250_, _05964_, _05286_);
  nor (_11251_, _11250_, _11235_);
  nor (_11252_, _11251_, _04081_);
  or (_11253_, _11252_, _11249_);
  and (_11254_, _11253_, _03996_);
  nor (_11255_, _11236_, _05204_);
  nor (_11256_, _11255_, _11235_);
  nor (_11257_, _11256_, _03996_);
  nor (_11258_, _11257_, _11254_);
  nor (_11259_, _11258_, _03729_);
  or (_11260_, _11259_, _07390_);
  nor (_11261_, _11260_, _11245_);
  and (_11262_, _11256_, _07390_);
  nor (_11263_, _11262_, _11261_);
  nor (_11264_, _11263_, _04481_);
  and (_11265_, _06069_, _05286_);
  nor (_11266_, _11235_, _07400_);
  not (_11267_, _11266_);
  nor (_11268_, _11267_, _11265_);
  or (_11269_, _11268_, _03222_);
  nor (_11270_, _11269_, _11264_);
  nor (_11271_, _06363_, _11236_);
  nor (_11272_, _11271_, _11235_);
  nor (_11273_, _11272_, _03589_);
  or (_11274_, _11273_, _03601_);
  nor (_11275_, _11274_, _11270_);
  nor (_11276_, _11275_, _11242_);
  or (_11277_, _11276_, _03600_);
  and (_11278_, _05884_, _05286_);
  or (_11279_, _11278_, _11235_);
  or (_11280_, _11279_, _07766_);
  and (_11281_, _11280_, _07778_);
  and (_11282_, _11281_, _11277_);
  and (_11283_, _06378_, _05286_);
  nor (_11284_, _11283_, _11235_);
  nor (_11285_, _11284_, _07778_);
  nor (_11286_, _11285_, _11282_);
  nor (_11287_, _11286_, _03622_);
  nor (_11288_, _11235_, _05310_);
  not (_11289_, _11288_);
  nor (_11290_, _11241_, _07777_);
  and (_11291_, _11290_, _11289_);
  nor (_11292_, _11291_, _11287_);
  nor (_11293_, _11292_, _03790_);
  nor (_11294_, _11244_, _06828_);
  and (_11295_, _11294_, _11289_);
  or (_11296_, _11295_, _11293_);
  and (_11297_, _11296_, _07795_);
  nor (_11298_, _05882_, _11236_);
  nor (_11299_, _11298_, _11235_);
  nor (_11300_, _11299_, _07795_);
  or (_11301_, _11300_, _11297_);
  and (_11302_, _11301_, _07793_);
  nor (_11303_, _11302_, _11239_);
  nor (_11304_, _11303_, _03815_);
  nor (_11305_, _11251_, _04246_);
  or (_11306_, _11305_, _03447_);
  nor (_11307_, _11306_, _11304_);
  and (_11308_, _05831_, _05286_);
  or (_11309_, _11235_, _03514_);
  nor (_11310_, _11309_, _11308_);
  nor (_11311_, _11310_, _11307_);
  or (_11312_, _11311_, _43004_);
  or (_11313_, _43000_, \oc8051_golden_model_1.TMOD [7]);
  and (_11314_, _11313_, _41806_);
  and (_40590_, _11314_, _11312_);
  not (_11315_, _02892_);
  and (_11316_, _06078_, _11315_);
  and (_11317_, _11316_, \oc8051_golden_model_1.PC [7]);
  and (_11318_, _11317_, \oc8051_golden_model_1.PC [8]);
  and (_11319_, _11318_, \oc8051_golden_model_1.PC [9]);
  and (_11320_, _11319_, \oc8051_golden_model_1.PC [10]);
  and (_11321_, _11320_, \oc8051_golden_model_1.PC [11]);
  and (_11322_, _11321_, \oc8051_golden_model_1.PC [12]);
  and (_11323_, _11322_, \oc8051_golden_model_1.PC [13]);
  and (_11324_, _11323_, \oc8051_golden_model_1.PC [14]);
  or (_11325_, _11324_, \oc8051_golden_model_1.PC [15]);
  nand (_11326_, _11324_, \oc8051_golden_model_1.PC [15]);
  and (_11327_, _11326_, _11325_);
  nor (_11328_, _08620_, _08618_);
  or (_11329_, _11328_, _11327_);
  and (_11330_, _08477_, _07898_);
  or (_11331_, _11330_, _11327_);
  nor (_11332_, _08441_, _04306_);
  and (_11333_, _03494_, _03200_);
  nor (_11334_, _08450_, _11333_);
  and (_11335_, _11334_, _11332_);
  or (_11336_, _11335_, _11327_);
  and (_11337_, _03191_, _03452_);
  not (_11338_, _11337_);
  or (_11339_, _10753_, _06813_);
  and (_11340_, _11339_, _11338_);
  nor (_11341_, _07904_, _03778_);
  not (_11342_, _11341_);
  nand (_11343_, _03181_, _02962_);
  not (_11344_, _11343_);
  nor (_11345_, _11344_, _08392_);
  or (_11346_, _11345_, _11327_);
  and (_11347_, _03599_, _03176_);
  not (_11348_, _11347_);
  and (_11349_, _06821_, _03222_);
  and (_11350_, _08059_, _10201_);
  or (_11351_, _11350_, _11327_);
  and (_11352_, _03751_, _03221_);
  not (_11353_, _11352_);
  nor (_11354_, _08847_, _06869_);
  and (_11355_, _11354_, _11353_);
  not (_11356_, _11355_);
  and (_11357_, _11356_, _11327_);
  not (_11358_, _10025_);
  and (_11359_, _06813_, _03729_);
  and (_11360_, _03730_, _03230_);
  or (_11361_, _11360_, _06813_);
  nor (_11362_, _09895_, _08089_);
  and (_11363_, _05666_, _05617_);
  and (_11364_, _05958_, _11363_);
  and (_11365_, _05411_, _05309_);
  and (_11366_, _11365_, _05955_);
  nand (_11367_, _11366_, _11364_);
  or (_11368_, _11367_, _06821_);
  and (_11369_, _11366_, _11364_);
  and (_11370_, _06746_, \oc8051_golden_model_1.PC [8]);
  and (_11371_, _11370_, \oc8051_golden_model_1.PC [9]);
  and (_11372_, _11371_, \oc8051_golden_model_1.PC [10]);
  and (_11373_, _11372_, \oc8051_golden_model_1.PC [11]);
  and (_11374_, _11373_, \oc8051_golden_model_1.PC [12]);
  and (_11375_, _11374_, \oc8051_golden_model_1.PC [13]);
  and (_11376_, _11375_, \oc8051_golden_model_1.PC [14]);
  nor (_11377_, _11375_, \oc8051_golden_model_1.PC [14]);
  nor (_11378_, _11377_, _11376_);
  not (_11379_, _11378_);
  nor (_11380_, _11379_, _05881_);
  and (_11381_, _11379_, _05881_);
  nor (_11382_, _11381_, _11380_);
  not (_11383_, _11382_);
  nor (_11384_, _11374_, \oc8051_golden_model_1.PC [13]);
  nor (_11385_, _11384_, _11375_);
  not (_11386_, _11385_);
  nor (_11387_, _11386_, _05881_);
  and (_11388_, _11386_, _05881_);
  nor (_11389_, _11373_, \oc8051_golden_model_1.PC [12]);
  nor (_11390_, _11389_, _11374_);
  not (_11391_, _11390_);
  nor (_11392_, _11391_, _05881_);
  nor (_11393_, _11371_, \oc8051_golden_model_1.PC [10]);
  nor (_11394_, _11393_, _11372_);
  not (_11395_, _11394_);
  nor (_11396_, _11395_, _05881_);
  not (_11397_, _11396_);
  nor (_11398_, _11372_, \oc8051_golden_model_1.PC [11]);
  nor (_11399_, _11398_, _11373_);
  not (_11400_, _11399_);
  nor (_11401_, _11400_, _05881_);
  and (_11402_, _11400_, _05881_);
  nor (_11403_, _11402_, _11401_);
  and (_11404_, _11395_, _05881_);
  nor (_11405_, _11404_, _11396_);
  and (_11406_, _11405_, _11403_);
  nor (_11407_, _11370_, \oc8051_golden_model_1.PC [9]);
  nor (_11408_, _11407_, _11371_);
  not (_11409_, _11408_);
  nor (_11410_, _11409_, _05881_);
  and (_11411_, _11409_, _05881_);
  nor (_11412_, _11411_, _11410_);
  nor (_11413_, _06749_, _05881_);
  and (_11414_, _06749_, _05881_);
  and (_11415_, _06744_, _06077_);
  nor (_11416_, _11415_, \oc8051_golden_model_1.PC [6]);
  nor (_11417_, _11416_, _06745_);
  not (_11418_, _11417_);
  nor (_11419_, _11418_, _06204_);
  and (_11420_, _11418_, _06204_);
  nor (_11421_, _11420_, _11419_);
  not (_11422_, _11421_);
  and (_11423_, _06744_, \oc8051_golden_model_1.PC [4]);
  nor (_11424_, _11423_, \oc8051_golden_model_1.PC [5]);
  nor (_11425_, _11424_, _11415_);
  not (_11426_, _11425_);
  nor (_11427_, _11426_, _06267_);
  and (_11428_, _11426_, _06267_);
  nor (_11429_, _06744_, \oc8051_golden_model_1.PC [4]);
  nor (_11430_, _11429_, _11423_);
  not (_11431_, _11430_);
  nor (_11432_, _11431_, _06236_);
  nor (_11433_, _06743_, \oc8051_golden_model_1.PC [3]);
  nor (_11434_, _11433_, _06744_);
  not (_11435_, _11434_);
  nor (_11436_, _11435_, _03708_);
  and (_11437_, _11435_, _03708_);
  nor (_11438_, _02909_, \oc8051_golden_model_1.PC [2]);
  nor (_11439_, _11438_, _06743_);
  not (_11440_, _11439_);
  nor (_11441_, _11440_, _03946_);
  not (_11442_, _03275_);
  nor (_11443_, _04303_, _11442_);
  nor (_11444_, _04163_, \oc8051_golden_model_1.PC [0]);
  and (_11445_, _04303_, _11442_);
  nor (_11446_, _11445_, _11443_);
  and (_11447_, _11446_, _11444_);
  nor (_11448_, _11447_, _11443_);
  and (_11449_, _11440_, _03946_);
  nor (_11450_, _11449_, _11441_);
  not (_11451_, _11450_);
  nor (_11452_, _11451_, _11448_);
  nor (_11453_, _11452_, _11441_);
  nor (_11454_, _11453_, _11437_);
  nor (_11455_, _11454_, _11436_);
  and (_11456_, _11431_, _06236_);
  nor (_11457_, _11456_, _11432_);
  not (_11458_, _11457_);
  nor (_11459_, _11458_, _11455_);
  nor (_11460_, _11459_, _11432_);
  nor (_11461_, _11460_, _11428_);
  nor (_11462_, _11461_, _11427_);
  nor (_11463_, _11462_, _11422_);
  nor (_11464_, _11463_, _11419_);
  nor (_11465_, _11464_, _11414_);
  or (_11466_, _11465_, _11413_);
  nor (_11467_, _06746_, \oc8051_golden_model_1.PC [8]);
  nor (_11468_, _11467_, _11370_);
  not (_11469_, _11468_);
  nor (_11470_, _11469_, _05881_);
  and (_11471_, _11469_, _05881_);
  nor (_11472_, _11471_, _11470_);
  and (_11473_, _11472_, _11466_);
  and (_11474_, _11473_, _11412_);
  and (_11475_, _11474_, _11406_);
  nor (_11476_, _11470_, _11410_);
  not (_11477_, _11476_);
  and (_11478_, _11477_, _11406_);
  or (_11479_, _11478_, _11401_);
  nor (_11480_, _11479_, _11475_);
  and (_11481_, _11480_, _11397_);
  and (_11482_, _11391_, _05881_);
  nor (_11483_, _11482_, _11392_);
  not (_11484_, _11483_);
  nor (_11485_, _11484_, _11481_);
  nor (_11486_, _11485_, _11392_);
  nor (_11487_, _11486_, _11388_);
  nor (_11488_, _11487_, _11387_);
  nor (_11489_, _11488_, _11383_);
  nor (_11490_, _11489_, _11380_);
  not (_11491_, _06821_);
  and (_11492_, _11491_, _05881_);
  nor (_11493_, _11491_, _05881_);
  nor (_11494_, _11493_, _11492_);
  and (_11495_, _11494_, _11490_);
  nor (_11496_, _11494_, _11490_);
  or (_11497_, _11496_, _11495_);
  or (_11498_, _11497_, _11369_);
  and (_11499_, _11498_, _03610_);
  and (_11500_, _11499_, _11368_);
  and (_11501_, _05836_, _05834_);
  and (_11502_, _04406_, _04620_);
  and (_11503_, _06770_, _11502_);
  and (_11504_, _11503_, _11501_);
  and (_11505_, _11504_, _06813_);
  and (_11506_, _06080_, \oc8051_golden_model_1.PC [8]);
  and (_11507_, _11506_, \oc8051_golden_model_1.PC [9]);
  and (_11508_, _11507_, \oc8051_golden_model_1.PC [10]);
  and (_11509_, _11508_, \oc8051_golden_model_1.PC [11]);
  and (_11510_, _11509_, \oc8051_golden_model_1.PC [12]);
  and (_11511_, _11510_, \oc8051_golden_model_1.PC [13]);
  and (_11512_, _11511_, \oc8051_golden_model_1.PC [14]);
  nor (_11513_, _11511_, \oc8051_golden_model_1.PC [14]);
  nor (_11514_, _11513_, _11512_);
  not (_11515_, _11514_);
  nor (_11516_, _11515_, _03446_);
  and (_11517_, _11515_, _03446_);
  nor (_11518_, _11517_, _11516_);
  not (_11519_, _11518_);
  nor (_11520_, _11510_, \oc8051_golden_model_1.PC [13]);
  nor (_11521_, _11520_, _11511_);
  and (_11522_, _11521_, _03454_);
  nor (_11523_, _11521_, _03454_);
  nor (_11524_, _11509_, \oc8051_golden_model_1.PC [12]);
  nor (_11525_, _11524_, _11510_);
  not (_11526_, _11525_);
  nor (_11527_, _11526_, _03446_);
  nor (_11528_, _11507_, \oc8051_golden_model_1.PC [10]);
  nor (_11529_, _11528_, _11508_);
  and (_11530_, _11529_, _03454_);
  not (_11531_, _11530_);
  nor (_11532_, _11508_, \oc8051_golden_model_1.PC [11]);
  nor (_11533_, _11532_, _11509_);
  not (_11534_, _11533_);
  nor (_11535_, _11534_, _03446_);
  and (_11536_, _11534_, _03446_);
  nor (_11537_, _11536_, _11535_);
  nor (_11538_, _11529_, _03454_);
  nor (_11539_, _11538_, _11530_);
  and (_11540_, _11539_, _11537_);
  nor (_11541_, _11506_, \oc8051_golden_model_1.PC [9]);
  nor (_11542_, _11541_, _11507_);
  not (_11543_, _11542_);
  nor (_11544_, _11543_, _03446_);
  and (_11545_, _11543_, _03446_);
  nor (_11546_, _11545_, _11544_);
  nor (_11547_, _06143_, _03446_);
  and (_11548_, _06143_, _03446_);
  and (_11549_, _06077_, _03295_);
  nor (_11550_, _11549_, \oc8051_golden_model_1.PC [6]);
  nor (_11551_, _11550_, _06079_);
  not (_11552_, _11551_);
  nor (_11553_, _11552_, _03549_);
  and (_11554_, _11552_, _03549_);
  nor (_11555_, _11554_, _11553_);
  not (_11556_, _11555_);
  and (_11557_, _03295_, \oc8051_golden_model_1.PC [4]);
  nor (_11558_, _11557_, \oc8051_golden_model_1.PC [5]);
  nor (_11559_, _11558_, _11549_);
  not (_11560_, _11559_);
  nor (_11561_, _11560_, _03860_);
  and (_11562_, _11560_, _03860_);
  nor (_11563_, _03295_, \oc8051_golden_model_1.PC [4]);
  nor (_11564_, _11563_, _11557_);
  not (_11565_, _11564_);
  nor (_11566_, _11565_, _03486_);
  nor (_11567_, _03581_, _03648_);
  and (_11568_, _03581_, _03648_);
  nor (_11569_, _03904_, _03245_);
  nor (_11570_, _03414_, \oc8051_golden_model_1.PC [1]);
  nor (_11571_, _04048_, _02905_);
  and (_11572_, _03414_, \oc8051_golden_model_1.PC [1]);
  nor (_11573_, _11572_, _11570_);
  and (_11574_, _11573_, _11571_);
  nor (_11575_, _11574_, _11570_);
  and (_11576_, _03904_, _03245_);
  nor (_11577_, _11576_, _11569_);
  not (_11578_, _11577_);
  nor (_11579_, _11578_, _11575_);
  nor (_11580_, _11579_, _11569_);
  nor (_11581_, _11580_, _11568_);
  nor (_11582_, _11581_, _11567_);
  and (_11583_, _11565_, _03486_);
  nor (_11584_, _11583_, _11566_);
  not (_11585_, _11584_);
  nor (_11586_, _11585_, _11582_);
  nor (_11587_, _11586_, _11566_);
  nor (_11588_, _11587_, _11562_);
  nor (_11589_, _11588_, _11561_);
  nor (_11590_, _11589_, _11556_);
  nor (_11591_, _11590_, _11553_);
  nor (_11592_, _11591_, _11548_);
  or (_11593_, _11592_, _11547_);
  nor (_11594_, _06080_, \oc8051_golden_model_1.PC [8]);
  nor (_11595_, _11594_, _11506_);
  not (_11596_, _11595_);
  nor (_11597_, _11596_, _03446_);
  and (_11598_, _11596_, _03446_);
  nor (_11599_, _11598_, _11597_);
  and (_11600_, _11599_, _11593_);
  and (_11601_, _11600_, _11546_);
  and (_11602_, _11601_, _11540_);
  nor (_11603_, _11597_, _11544_);
  not (_11604_, _11603_);
  and (_11605_, _11604_, _11540_);
  or (_11606_, _11605_, _11535_);
  nor (_11607_, _11606_, _11602_);
  and (_11608_, _11607_, _11531_);
  and (_11609_, _11526_, _03446_);
  nor (_11610_, _11609_, _11527_);
  not (_11611_, _11610_);
  nor (_11612_, _11611_, _11608_);
  nor (_11613_, _11612_, _11527_);
  nor (_11614_, _11613_, _11523_);
  nor (_11615_, _11614_, _11522_);
  nor (_11616_, _11615_, _11519_);
  nor (_11617_, _11616_, _11516_);
  and (_11618_, _06814_, _03446_);
  nor (_11619_, _06814_, _03446_);
  nor (_11620_, _11619_, _11618_);
  and (_11621_, _11620_, _11617_);
  nor (_11622_, _11620_, _11617_);
  or (_11623_, _11622_, _11621_);
  nand (_11624_, _11503_, _11501_);
  and (_11625_, _11624_, _11623_);
  or (_11626_, _11625_, _06072_);
  or (_11627_, _11626_, _11505_);
  nor (_11628_, _04622_, _03234_);
  not (_11629_, _11628_);
  and (_11630_, _11629_, _08078_);
  not (_11631_, _11630_);
  and (_11632_, _03979_, _02994_);
  nand (_11633_, _06814_, _03979_);
  nor (_11634_, _04729_, _03980_);
  nor (_11635_, _04409_, \oc8051_golden_model_1.PC [15]);
  nand (_11636_, _11635_, _11634_);
  and (_11637_, _11636_, _11633_);
  or (_11638_, _11637_, _11632_);
  nand (_11639_, _06814_, _03980_);
  and (_11640_, _11639_, _11638_);
  or (_11641_, _11640_, _11631_);
  nor (_11642_, _04729_, _11632_);
  and (_11643_, _11642_, _11630_);
  or (_11644_, _11643_, _11327_);
  and (_11645_, _11644_, _11641_);
  or (_11646_, _11645_, _06073_);
  nor (_11647_, _04422_, _03610_);
  and (_11648_, _11647_, _11646_);
  and (_11649_, _11648_, _11627_);
  or (_11650_, _11649_, _11500_);
  and (_11651_, _11650_, _11362_);
  not (_11652_, _11360_);
  and (_11653_, _11362_, _05966_);
  not (_11654_, _11653_);
  and (_11655_, _11654_, _11327_);
  or (_11656_, _11655_, _11652_);
  or (_11657_, _11656_, _11651_);
  and (_11658_, _11657_, _11361_);
  and (_11659_, _08063_, _08128_);
  not (_11660_, _11659_);
  or (_11661_, _11660_, _11658_);
  or (_11662_, _11659_, _11327_);
  and (_11663_, _11662_, _03737_);
  and (_11664_, _11663_, _11661_);
  or (_11665_, _11664_, _11359_);
  nor (_11666_, _09909_, _08132_);
  and (_11667_, _11666_, _11665_);
  not (_11668_, _11666_);
  and (_11669_, _11668_, _11327_);
  not (_11670_, _03233_);
  nor (_11671_, _03508_, _11670_);
  and (_11672_, _11671_, _03736_);
  not (_11673_, _11672_);
  or (_11674_, _11673_, _11669_);
  or (_11675_, _11674_, _11667_);
  or (_11676_, _11672_, _06813_);
  and (_11677_, _11676_, _09921_);
  and (_11678_, _11677_, _11675_);
  or (_11679_, _11497_, _09969_);
  nand (_11680_, _09969_, _11491_);
  and (_11681_, _11680_, _09917_);
  and (_11682_, _11681_, _11679_);
  or (_11683_, _11682_, _09919_);
  or (_11684_, _11683_, _11678_);
  and (_11685_, _10017_, _10006_);
  and (_11686_, _11685_, _06821_);
  and (_11687_, _11497_, _10018_);
  or (_11688_, _11687_, _11686_);
  or (_11689_, _11688_, _09920_);
  and (_11690_, _11689_, _11684_);
  or (_11691_, _11690_, _03615_);
  and (_11692_, _09876_, _06821_);
  not (_11693_, _09876_);
  and (_11694_, _11497_, _11693_);
  or (_11695_, _11694_, _04107_);
  or (_11696_, _11695_, _11692_);
  and (_11697_, _11696_, _09856_);
  and (_11698_, _11697_, _11691_);
  or (_11699_, _11497_, _10061_);
  nand (_11700_, _10061_, _11491_);
  and (_11701_, _11700_, _03604_);
  and (_11702_, _11701_, _11699_);
  or (_11703_, _11702_, _11698_);
  and (_11704_, _11703_, _11358_);
  nand (_11705_, _11327_, _10025_);
  nor (_11706_, _04746_, _03718_);
  and (_11707_, _11706_, _03227_);
  and (_11708_, _03593_, _03751_);
  not (_11709_, _11708_);
  and (_11710_, _11709_, _11707_);
  nor (_11711_, _08070_, _03237_);
  not (_11712_, _11711_);
  nor (_11713_, _03616_, _03494_);
  nor (_11714_, _11713_, _03237_);
  and (_11715_, _04066_, _03751_);
  or (_11716_, _04115_, _03719_);
  or (_11717_, _11716_, _11715_);
  nor (_11718_, _11717_, _11714_);
  and (_11719_, _11718_, _11712_);
  and (_11720_, _11719_, _11710_);
  nand (_11721_, _11720_, _11705_);
  or (_11722_, _11721_, _11704_);
  or (_11723_, _11720_, _06813_);
  and (_11724_, _11723_, _11355_);
  and (_11725_, _11724_, _11722_);
  or (_11726_, _11725_, _11357_);
  not (_11727_, _03238_);
  nor (_11728_, _03752_, _11727_);
  and (_11729_, _11728_, _09669_);
  and (_11730_, _11729_, _11726_);
  or (_11731_, _11729_, _06814_);
  nand (_11732_, _11731_, _11350_);
  or (_11733_, _11732_, _11730_);
  and (_11734_, _11733_, _11351_);
  or (_11735_, _11734_, _08187_);
  or (_11736_, _08186_, _06813_);
  and (_11737_, _11736_, _03248_);
  and (_11738_, _11737_, _11735_);
  and (_11739_, _11327_, _07912_);
  nor (_11740_, _03505_, _03224_);
  not (_11741_, _11740_);
  or (_11742_, _11741_, _11739_);
  or (_11743_, _11742_, _11738_);
  or (_11744_, _11740_, _06813_);
  and (_11745_, _11744_, _08832_);
  and (_11746_, _11745_, _11743_);
  nand (_11747_, _06821_, _03625_);
  nor (_11748_, _04481_, _06833_);
  and (_11749_, _11748_, _06837_);
  nand (_11750_, _11749_, _11747_);
  or (_11751_, _11750_, _11746_);
  or (_11752_, _11749_, _06813_);
  and (_11753_, _11752_, _03589_);
  and (_11754_, _11753_, _11751_);
  or (_11755_, _11754_, _11349_);
  nor (_11756_, _07405_, _03216_);
  and (_11757_, _11756_, _11755_);
  not (_11758_, _11756_);
  and (_11759_, _11758_, _11327_);
  nor (_11760_, _03585_, _03169_);
  not (_11761_, _11760_);
  or (_11762_, _11761_, _11759_);
  or (_11763_, _11762_, _11757_);
  and (_11764_, _03168_, _03452_);
  not (_11765_, _11764_);
  or (_11766_, _11760_, _06813_);
  and (_11767_, _11766_, _11765_);
  and (_11768_, _11767_, _11763_);
  and (_11769_, _11764_, _11623_);
  or (_11770_, _11769_, _06168_);
  or (_11771_, _11770_, _11768_);
  or (_11772_, _06813_, _05894_);
  and (_11773_, _11772_, _11771_);
  or (_11774_, _11773_, _03601_);
  nand (_11775_, _11491_, _03601_);
  and (_11776_, _11775_, _08364_);
  and (_11777_, _11776_, _11774_);
  and (_11778_, _08363_, _06813_);
  or (_11779_, _11778_, _11777_);
  and (_11780_, _11779_, _11348_);
  and (_11781_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_11782_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_11783_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_11784_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_11785_, _11784_, _11783_);
  not (_11786_, _11785_);
  and (_11787_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_11788_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_11789_, _11788_, _11787_);
  not (_11790_, _11789_);
  and (_11791_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_11792_, _03305_, _03301_);
  nor (_11793_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_11794_, _11793_, _11791_);
  not (_11795_, _11794_);
  nor (_11796_, _11795_, _11792_);
  nor (_11797_, _11796_, _11791_);
  nor (_11798_, _11797_, _11790_);
  nor (_11799_, _11798_, _11787_);
  nor (_11800_, _11799_, _11786_);
  nor (_11801_, _11800_, _11783_);
  nor (_11802_, _11801_, _11782_);
  or (_11803_, _11802_, _11781_);
  and (_11804_, _11803_, \oc8051_golden_model_1.DPH [0]);
  and (_11805_, _11804_, \oc8051_golden_model_1.DPH [1]);
  and (_11806_, _11805_, \oc8051_golden_model_1.DPH [2]);
  and (_11807_, _11806_, \oc8051_golden_model_1.DPH [3]);
  and (_11808_, _11807_, \oc8051_golden_model_1.DPH [4]);
  and (_11809_, _11808_, \oc8051_golden_model_1.DPH [5]);
  and (_11810_, _11809_, \oc8051_golden_model_1.DPH [6]);
  nand (_11811_, _11810_, \oc8051_golden_model_1.DPH [7]);
  or (_11812_, _11810_, \oc8051_golden_model_1.DPH [7]);
  and (_11813_, _11812_, _11347_);
  and (_11814_, _11813_, _11811_);
  nor (_11815_, _03584_, _03178_);
  not (_11816_, _11815_);
  or (_11817_, _11816_, _11814_);
  or (_11818_, _11817_, _11780_);
  and (_11819_, _03176_, _03452_);
  not (_11820_, _11819_);
  or (_11821_, _11815_, _06813_);
  and (_11822_, _11821_, _11820_);
  and (_11823_, _11822_, _11818_);
  not (_11824_, _11345_);
  or (_11825_, _11623_, _08786_);
  not (_11826_, _08786_);
  or (_11827_, _11826_, _06813_);
  and (_11828_, _11827_, _11819_);
  and (_11829_, _11828_, _11825_);
  or (_11830_, _11829_, _11824_);
  or (_11831_, _11830_, _11823_);
  and (_11832_, _11831_, _11346_);
  or (_11833_, _11832_, _11342_);
  or (_11834_, _11341_, _06813_);
  and (_11835_, _11834_, _07766_);
  and (_11836_, _11835_, _11833_);
  nand (_11837_, _06821_, _03600_);
  nor (_11838_, _03780_, _03182_);
  nand (_11839_, _11838_, _11837_);
  or (_11840_, _11839_, _11836_);
  and (_11841_, _03181_, _03452_);
  not (_11842_, _11841_);
  or (_11843_, _11838_, _06813_);
  and (_11844_, _11843_, _11842_);
  and (_11845_, _11844_, _11840_);
  or (_11846_, _11623_, _11826_);
  or (_11847_, _08786_, _06813_);
  and (_11848_, _11847_, _11841_);
  and (_11849_, _11848_, _11846_);
  or (_11850_, _11849_, _11845_);
  and (_11851_, _08425_, _08417_);
  and (_11852_, _11851_, _11850_);
  not (_11853_, _11851_);
  and (_11854_, _11853_, _11327_);
  or (_11855_, _11854_, _08431_);
  or (_11856_, _11855_, _11852_);
  or (_11857_, _08430_, _06813_);
  and (_11858_, _11857_, _07777_);
  and (_11859_, _11858_, _11856_);
  nand (_11860_, _06821_, _03622_);
  nand (_11861_, _11860_, _10753_);
  or (_11862_, _11861_, _11859_);
  and (_11863_, _11862_, _11340_);
  not (_11864_, _11335_);
  or (_11865_, _11623_, \oc8051_golden_model_1.PSW [7]);
  or (_11866_, _06813_, _07871_);
  and (_11867_, _11866_, _11337_);
  and (_11868_, _11867_, _11865_);
  or (_11869_, _11868_, _11864_);
  or (_11870_, _11869_, _11863_);
  and (_11871_, _11870_, _11336_);
  or (_11872_, _11871_, _08460_);
  or (_11873_, _08459_, _06813_);
  and (_11874_, _11873_, _07795_);
  and (_11875_, _11874_, _11872_);
  nand (_11876_, _06821_, _03624_);
  nor (_11877_, _03785_, _03201_);
  nand (_11878_, _11877_, _11876_);
  or (_11879_, _11878_, _11875_);
  and (_11880_, _03200_, _03452_);
  not (_11881_, _11880_);
  or (_11882_, _11877_, _06813_);
  and (_11883_, _11882_, _11881_);
  and (_11884_, _11883_, _11879_);
  not (_11885_, _11330_);
  or (_11886_, _11623_, _07871_);
  or (_11887_, _06813_, \oc8051_golden_model_1.PSW [7]);
  and (_11888_, _11887_, _11880_);
  and (_11889_, _11888_, _11886_);
  or (_11890_, _11889_, _11885_);
  or (_11891_, _11890_, _11884_);
  and (_11892_, _11891_, _11331_);
  or (_11893_, _11892_, _08508_);
  or (_11894_, _08507_, _06813_);
  and (_11895_, _11894_, _08588_);
  and (_11896_, _11895_, _11893_);
  and (_11897_, _11327_, _08587_);
  or (_11898_, _11897_, _03798_);
  or (_11899_, _11898_, _11896_);
  nand (_11900_, _05204_, _03798_);
  and (_11901_, _11900_, _11899_);
  or (_11902_, _11901_, _03188_);
  not (_11903_, _03621_);
  nand (_11904_, _06814_, _03188_);
  and (_11905_, _11904_, _11903_);
  and (_11906_, _11905_, _11902_);
  not (_11907_, _11328_);
  not (_11908_, _09854_);
  or (_11909_, _11497_, _11908_);
  or (_11910_, _09854_, _06821_);
  and (_11911_, _11910_, _03621_);
  and (_11912_, _11911_, _11909_);
  or (_11913_, _11912_, _11907_);
  or (_11914_, _11913_, _11906_);
  and (_11915_, _11914_, _11329_);
  or (_11916_, _11915_, _08703_);
  or (_11917_, _08702_, _06813_);
  and (_11918_, _11917_, _08733_);
  and (_11919_, _11918_, _11916_);
  and (_11920_, _11327_, _08732_);
  or (_11921_, _11920_, _03515_);
  or (_11922_, _11921_, _11919_);
  nand (_11923_, _05204_, _03515_);
  and (_11924_, _11923_, _11922_);
  or (_11925_, _11924_, _03203_);
  nand (_11926_, _06814_, _03203_);
  and (_11927_, _11926_, _03816_);
  and (_11928_, _11927_, _11925_);
  or (_11929_, _11497_, _09854_);
  nand (_11930_, _09854_, _11491_);
  and (_11931_, _11930_, _11929_);
  and (_11932_, _11931_, _03628_);
  and (_11933_, _05848_, _06409_);
  not (_11934_, _11933_);
  or (_11935_, _11934_, _11932_);
  or (_11936_, _11935_, _11928_);
  or (_11937_, _11933_, _11327_);
  and (_11938_, _11937_, _04246_);
  and (_11939_, _11938_, _11936_);
  nor (_11940_, _08780_, _08775_);
  nand (_11941_, _06813_, _03815_);
  nand (_11942_, _11941_, _11940_);
  or (_11943_, _11942_, _11939_);
  not (_11944_, _03629_);
  or (_11945_, _11327_, _11940_);
  and (_11946_, _11945_, _11944_);
  and (_11947_, _11946_, _11943_);
  nor (_11948_, _11944_, _03446_);
  or (_11949_, _11948_, _03198_);
  or (_11950_, _11949_, _11947_);
  nand (_11951_, _06814_, _03198_);
  and (_11952_, _11951_, _03823_);
  and (_11953_, _11952_, _11950_);
  and (_11954_, _11931_, _03453_);
  nand (_11955_, _03195_, _02962_);
  not (_11956_, _11955_);
  nor (_11957_, _11956_, _04552_);
  not (_11958_, _11957_);
  or (_11959_, _11958_, _11954_);
  or (_11960_, _11959_, _11953_);
  or (_11961_, _11957_, _11327_);
  and (_11962_, _11961_, _03514_);
  and (_11963_, _11962_, _11960_);
  nor (_11964_, _08805_, _08798_);
  nand (_11965_, _06813_, _03447_);
  nand (_11966_, _11965_, _11964_);
  or (_11967_, _11966_, _11963_);
  not (_11968_, _03631_);
  or (_11969_, _11327_, _11964_);
  and (_11970_, _11969_, _11968_);
  and (_11971_, _11970_, _11967_);
  nor (_11972_, _11968_, _03446_);
  or (_11973_, _11972_, _03196_);
  or (_11974_, _11973_, _11971_);
  and (_11975_, _03195_, _03452_);
  not (_11976_, _11975_);
  nand (_11977_, _06814_, _03196_);
  and (_11978_, _11977_, _11976_);
  and (_11979_, _11978_, _11974_);
  and (_11980_, _11975_, _11327_);
  or (_11981_, _11980_, _11979_);
  or (_11982_, _11981_, _43004_);
  or (_11983_, _43000_, \oc8051_golden_model_1.PC [15]);
  and (_11984_, _11983_, _41806_);
  and (_40591_, _11984_, _11982_);
  and (_11985_, _43004_, \oc8051_golden_model_1.P0INREG [7]);
  or (_11986_, _11985_, _01195_);
  and (_40592_, _11986_, _41806_);
  and (_11987_, _43004_, \oc8051_golden_model_1.P1INREG [7]);
  or (_11988_, _11987_, _01092_);
  and (_40593_, _11988_, _41806_);
  and (_11989_, _43004_, \oc8051_golden_model_1.P2INREG [7]);
  or (_11990_, _11989_, _00908_);
  and (_40595_, _11990_, _41806_);
  and (_11991_, _43004_, \oc8051_golden_model_1.P3INREG [7]);
  or (_11992_, _11991_, _01028_);
  and (_40596_, _11992_, _41806_);
  nor (_11993_, _04797_, _04556_);
  nor (_11994_, _11993_, _04798_);
  nor (_11995_, _04797_, _04951_);
  nor (_11996_, _11995_, _05123_);
  and (_11997_, _11996_, _04796_);
  and (_11998_, _11997_, _11994_);
  not (_11999_, _11998_);
  nand (_12000_, _03198_, _02905_);
  or (_12001_, _04533_, _04634_);
  and (_12002_, _12001_, _11934_);
  nor (_12003_, _05666_, \oc8051_golden_model_1.ACC [0]);
  nand (_12004_, _12003_, _06394_);
  and (_12005_, _05666_, \oc8051_golden_model_1.ACC [0]);
  or (_12006_, _12005_, _06382_);
  or (_12007_, _04480_, _04620_);
  nand (_12008_, _08285_, _03745_);
  nor (_12009_, _10122_, _05224_);
  or (_12010_, _12009_, _05940_);
  or (_12011_, _06072_, _04634_);
  nand (_12012_, _03980_, _02905_);
  or (_12013_, _03980_, \oc8051_golden_model_1.ACC [0]);
  and (_12014_, _12013_, _12012_);
  nor (_12015_, _12014_, _06073_);
  nor (_12016_, _12015_, _04421_);
  and (_12017_, _12016_, _12011_);
  nor (_12018_, _05666_, _06071_);
  or (_12019_, _12018_, _12017_);
  and (_12020_, _12019_, _05954_);
  nand (_12021_, _10122_, _09750_);
  and (_12022_, _12021_, _04428_);
  or (_12023_, _12022_, _04768_);
  or (_12024_, _12023_, _12020_);
  nor (_12025_, _03230_, \oc8051_golden_model_1.PC [0]);
  nor (_12026_, _12025_, _04431_);
  and (_12027_, _12026_, _12024_);
  and (_12028_, _04431_, _04620_);
  or (_12029_, _12028_, _04449_);
  or (_12030_, _12029_, _12027_);
  and (_12031_, _12030_, _12010_);
  or (_12032_, _12031_, _03508_);
  nand (_12033_, _08285_, _03508_);
  and (_12034_, _12033_, _04562_);
  and (_12035_, _12034_, _12032_);
  nor (_12036_, _10123_, _04562_);
  and (_12037_, _12036_, _12021_);
  or (_12038_, _12037_, _12035_);
  and (_12039_, _12038_, _03227_);
  nor (_12040_, _03227_, _02905_);
  or (_12041_, _03745_, _12040_);
  or (_12042_, _12041_, _12039_);
  and (_12043_, _12042_, _12008_);
  or (_12044_, _12043_, _04463_);
  and (_12045_, _06546_, _03446_);
  nand (_12046_, _08284_, _04463_);
  or (_12047_, _12046_, _12045_);
  and (_12048_, _12047_, _12044_);
  or (_12049_, _12048_, _04462_);
  nor (_12050_, _09773_, _05224_);
  and (_12051_, _05224_, \oc8051_golden_model_1.PSW [7]);
  nor (_12052_, _12051_, _12050_);
  nand (_12053_, _12052_, _04462_);
  and (_12054_, _12053_, _05897_);
  and (_12055_, _12054_, _12049_);
  nand (_12056_, _03224_, \oc8051_golden_model_1.PC [0]);
  nand (_12057_, _04480_, _12056_);
  or (_12058_, _12057_, _12055_);
  and (_12059_, _12058_, _12007_);
  or (_12060_, _12059_, _04482_);
  or (_12061_, _06546_, _06164_);
  and (_12062_, _12061_, _06163_);
  and (_12063_, _12062_, _12060_);
  and (_12064_, _05881_, _04620_);
  and (_12065_, _06340_, \oc8051_golden_model_1.P1INREG [0]);
  not (_12066_, _12065_);
  and (_12067_, _06343_, \oc8051_golden_model_1.P0INREG [0]);
  not (_12068_, _12067_);
  and (_12069_, _06346_, \oc8051_golden_model_1.P2INREG [0]);
  and (_12070_, _06348_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_12071_, _12070_, _12069_);
  and (_12072_, _12071_, _12068_);
  and (_12073_, _12072_, _12066_);
  and (_12074_, _06354_, \oc8051_golden_model_1.SP [0]);
  and (_12075_, _06284_, \oc8051_golden_model_1.TL0 [0]);
  nor (_12076_, _12075_, _12074_);
  and (_12077_, _12076_, _12073_);
  and (_12078_, _06315_, \oc8051_golden_model_1.IE [0]);
  and (_12079_, _06319_, \oc8051_golden_model_1.SBUF [0]);
  and (_12080_, _06321_, \oc8051_golden_model_1.SCON [0]);
  or (_12081_, _12080_, _12079_);
  nor (_12082_, _12081_, _12078_);
  and (_12083_, _06296_, \oc8051_golden_model_1.IP [0]);
  and (_12084_, _06310_, \oc8051_golden_model_1.B [0]);
  nor (_12085_, _12084_, _12083_);
  and (_12086_, _06303_, \oc8051_golden_model_1.PSW [0]);
  and (_12087_, _06308_, \oc8051_golden_model_1.ACC [0]);
  nor (_12088_, _12087_, _12086_);
  and (_12089_, _12088_, _12085_);
  and (_12090_, _12089_, _12082_);
  and (_12091_, _12090_, _12077_);
  and (_12092_, _06327_, \oc8051_golden_model_1.TH0 [0]);
  and (_12093_, _06329_, \oc8051_golden_model_1.TL1 [0]);
  nor (_12094_, _12093_, _12092_);
  and (_12095_, _06334_, \oc8051_golden_model_1.PCON [0]);
  and (_12096_, _06336_, \oc8051_golden_model_1.TCON [0]);
  nor (_12097_, _12096_, _12095_);
  and (_12098_, _12097_, _12094_);
  and (_12099_, _06272_, \oc8051_golden_model_1.DPH [0]);
  and (_12100_, _06279_, \oc8051_golden_model_1.TMOD [0]);
  nor (_12101_, _12100_, _12099_);
  and (_12102_, _06356_, \oc8051_golden_model_1.DPL [0]);
  and (_12103_, _06288_, \oc8051_golden_model_1.TH1 [0]);
  nor (_12104_, _12103_, _12102_);
  and (_12105_, _12104_, _12101_);
  and (_12106_, _12105_, _12098_);
  and (_12107_, _12106_, _12091_);
  not (_12108_, _12107_);
  nor (_12109_, _12108_, _12064_);
  nor (_12110_, _12109_, _06170_);
  or (_12111_, _12110_, _06168_);
  or (_12112_, _12111_, _12063_);
  and (_12113_, _06168_, _04048_);
  nor (_12114_, _12113_, _04500_);
  and (_12115_, _12114_, _12112_);
  and (_12116_, _04500_, _06274_);
  or (_12117_, _12116_, _03178_);
  or (_12118_, _12117_, _12115_);
  and (_12119_, _03178_, _02905_);
  nor (_12120_, _12119_, _04512_);
  and (_12121_, _12120_, _12118_);
  nor (_12122_, _05666_, _06274_);
  and (_12123_, _05666_, _06274_);
  nor (_12124_, _12123_, _12122_);
  nor (_12125_, _12124_, _04511_);
  nor (_12126_, _12125_, _04513_);
  or (_12127_, _12126_, _12121_);
  nor (_12128_, _12005_, _12003_);
  or (_12129_, _12128_, _05850_);
  and (_12130_, _12129_, _06383_);
  and (_12131_, _12130_, _12127_);
  and (_12132_, _12123_, _04515_);
  or (_12133_, _12132_, _04514_);
  or (_12134_, _12133_, _12131_);
  and (_12135_, _12134_, _12006_);
  or (_12136_, _12135_, _03192_);
  and (_12137_, _03192_, _02905_);
  nor (_12138_, _12137_, _06390_);
  and (_12139_, _12138_, _12136_);
  nor (_12140_, _12122_, _06395_);
  or (_12141_, _12140_, _06394_);
  or (_12142_, _12141_, _12139_);
  and (_12143_, _12142_, _12004_);
  or (_12144_, _12143_, _03188_);
  nand (_12145_, _03188_, _02905_);
  and (_12146_, _12145_, _05848_);
  and (_12147_, _12146_, _12144_);
  or (_12148_, _12147_, _12002_);
  nand (_12149_, _06546_, _04533_);
  and (_12150_, _12149_, _12148_);
  or (_12151_, _12150_, _04531_);
  nand (_12152_, _05666_, _04531_);
  and (_12153_, _12152_, _11944_);
  and (_12154_, _12153_, _12151_);
  and (_12155_, _03629_, _02905_);
  or (_12156_, _12155_, _03198_);
  or (_12157_, _12156_, _12154_);
  and (_12158_, _12157_, _12000_);
  or (_12159_, _12158_, _04539_);
  or (_12160_, _12050_, _04558_);
  and (_12161_, _12160_, _11955_);
  and (_12162_, _12161_, _12159_);
  or (_12163_, _04552_, _04634_);
  and (_12164_, _12163_, _11958_);
  or (_12165_, _12164_, _12162_);
  nand (_12166_, _06546_, _04552_);
  and (_12167_, _12166_, _12165_);
  or (_12168_, _12167_, _03448_);
  nand (_12169_, _05666_, _03448_);
  and (_12170_, _12169_, _04796_);
  and (_12171_, _12170_, _12168_);
  or (_12172_, _12171_, _11999_);
  not (_12173_, _00000_);
  nor (_12174_, _04793_, _12173_);
  not (_12175_, _12174_);
  nor (_12176_, _04951_, _12175_);
  nor (_12177_, _05122_, _12175_);
  nor (_12178_, _12177_, _12176_);
  nor (_12179_, _12175_, _04556_);
  nor (_12180_, _12175_, _04711_);
  nor (_12181_, _12180_, _12179_);
  and (_12182_, _12181_, _12174_);
  and (_12183_, _12182_, _12178_);
  or (_12184_, _12183_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_12185_, _05137_, _05129_);
  nor (_12186_, _12185_, _05138_);
  and (_12187_, _12186_, _05137_);
  nand (_12188_, _12187_, _03499_);
  and (_12189_, _12188_, _12184_);
  and (_12190_, _12189_, _12172_);
  nor (_12191_, _05136_, _12173_);
  not (_12192_, _05129_);
  and (_12193_, _12192_, _05132_);
  and (_12194_, _12193_, _12191_);
  and (_12195_, _12194_, _03499_);
  and (_12196_, _11468_, _03629_);
  nor (_12197_, _11596_, _03629_);
  or (_12198_, _12197_, _12196_);
  and (_12199_, _12198_, _12195_);
  or (_40634_, _12199_, _12190_);
  not (_12200_, _12195_);
  or (_12201_, _12183_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_12202_, _12201_, _12200_);
  nor (_12203_, _06786_, _06547_);
  or (_12204_, _12203_, _06785_);
  nor (_12205_, _06765_, _05835_);
  nand (_12206_, _12205_, _03972_);
  nor (_12207_, _05617_, _04303_);
  and (_12208_, _12207_, _04515_);
  or (_12209_, _06764_, _04480_);
  nand (_12210_, _08271_, _03745_);
  nor (_12211_, _10095_, _05216_);
  or (_12212_, _12211_, _05940_);
  nor (_12213_, _05957_, _05667_);
  nor (_12214_, _12213_, _06071_);
  nand (_12215_, _12205_, _06073_);
  and (_12216_, _03980_, _02878_);
  nor (_12217_, _03980_, _03274_);
  or (_12218_, _12217_, _12216_);
  nor (_12219_, _12218_, _06073_);
  nor (_12220_, _12219_, _04421_);
  and (_12221_, _12220_, _12215_);
  or (_12222_, _12221_, _04428_);
  or (_12223_, _12222_, _12214_);
  nand (_12224_, _10095_, _09695_);
  or (_12225_, _12224_, _05954_);
  and (_12226_, _12225_, _12223_);
  or (_12227_, _12226_, _04768_);
  nor (_12228_, _03230_, _02878_);
  nor (_12229_, _12228_, _04431_);
  and (_12230_, _12229_, _12227_);
  and (_12231_, _06764_, _04431_);
  or (_12232_, _12231_, _04449_);
  or (_12233_, _12232_, _12230_);
  and (_12234_, _12233_, _12212_);
  or (_12235_, _12234_, _03508_);
  nand (_12236_, _08271_, _03508_);
  and (_12237_, _12236_, _04562_);
  and (_12238_, _12237_, _12235_);
  not (_12239_, _10096_);
  and (_12240_, _12224_, _12239_);
  and (_12241_, _12240_, _04454_);
  or (_12242_, _12241_, _12238_);
  and (_12243_, _12242_, _03227_);
  nor (_12244_, _03227_, \oc8051_golden_model_1.PC [1]);
  or (_12245_, _03745_, _12244_);
  or (_12246_, _12245_, _12243_);
  and (_12247_, _12246_, _12210_);
  or (_12248_, _12247_, _04463_);
  and (_12249_, _06501_, _03446_);
  nand (_12250_, _08270_, _04463_);
  or (_12251_, _12250_, _12249_);
  and (_12252_, _12251_, _12248_);
  or (_12253_, _12252_, _04462_);
  nor (_12254_, _09718_, _05216_);
  and (_12255_, _05216_, \oc8051_golden_model_1.PSW [7]);
  nor (_12256_, _12255_, _12254_);
  nand (_12257_, _12256_, _04462_);
  and (_12258_, _12257_, _05897_);
  and (_12259_, _12258_, _12253_);
  nand (_12260_, _03224_, _02878_);
  nand (_12261_, _04480_, _12260_);
  or (_12262_, _12261_, _12259_);
  and (_12263_, _12262_, _12209_);
  or (_12264_, _12263_, _04482_);
  or (_12265_, _06501_, _06164_);
  and (_12266_, _12265_, _06163_);
  and (_12267_, _12266_, _12264_);
  and (_12268_, _05881_, _06764_);
  and (_12269_, _06340_, \oc8051_golden_model_1.P1INREG [1]);
  not (_12270_, _12269_);
  and (_12271_, _06343_, \oc8051_golden_model_1.P0INREG [1]);
  not (_12272_, _12271_);
  and (_12273_, _06346_, \oc8051_golden_model_1.P2INREG [1]);
  and (_12274_, _06348_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_12275_, _12274_, _12273_);
  and (_12276_, _12275_, _12272_);
  and (_12277_, _12276_, _12270_);
  and (_12278_, _06354_, \oc8051_golden_model_1.SP [1]);
  and (_12279_, _06284_, \oc8051_golden_model_1.TL0 [1]);
  nor (_12280_, _12279_, _12278_);
  and (_12281_, _12280_, _12277_);
  and (_12282_, _06315_, \oc8051_golden_model_1.IE [1]);
  and (_12283_, _06319_, \oc8051_golden_model_1.SBUF [1]);
  and (_12284_, _06321_, \oc8051_golden_model_1.SCON [1]);
  or (_12285_, _12284_, _12283_);
  nor (_12286_, _12285_, _12282_);
  and (_12287_, _06296_, \oc8051_golden_model_1.IP [1]);
  and (_12288_, _06310_, \oc8051_golden_model_1.B [1]);
  nor (_12289_, _12288_, _12287_);
  and (_12290_, _06303_, \oc8051_golden_model_1.PSW [1]);
  and (_12291_, _06308_, \oc8051_golden_model_1.ACC [1]);
  nor (_12292_, _12291_, _12290_);
  and (_12293_, _12292_, _12289_);
  and (_12294_, _12293_, _12286_);
  and (_12295_, _12294_, _12281_);
  and (_12296_, _06327_, \oc8051_golden_model_1.TH0 [1]);
  and (_12297_, _06329_, \oc8051_golden_model_1.TL1 [1]);
  nor (_12298_, _12297_, _12296_);
  and (_12299_, _06334_, \oc8051_golden_model_1.PCON [1]);
  and (_12300_, _06336_, \oc8051_golden_model_1.TCON [1]);
  nor (_12301_, _12300_, _12299_);
  and (_12302_, _12301_, _12298_);
  and (_12303_, _06272_, \oc8051_golden_model_1.DPH [1]);
  and (_12304_, _06279_, \oc8051_golden_model_1.TMOD [1]);
  nor (_12305_, _12304_, _12303_);
  and (_12306_, _06356_, \oc8051_golden_model_1.DPL [1]);
  and (_12307_, _06288_, \oc8051_golden_model_1.TH1 [1]);
  nor (_12308_, _12307_, _12306_);
  and (_12309_, _12308_, _12305_);
  and (_12310_, _12309_, _12302_);
  and (_12311_, _12310_, _12295_);
  not (_12312_, _12311_);
  nor (_12313_, _12312_, _12268_);
  nor (_12314_, _12313_, _06170_);
  or (_12315_, _12314_, _06168_);
  or (_12316_, _12315_, _12267_);
  and (_12317_, _06168_, _03414_);
  nor (_12318_, _12317_, _04500_);
  and (_12319_, _12318_, _12316_);
  and (_12320_, _04500_, _06282_);
  or (_12321_, _12320_, _03178_);
  or (_12322_, _12321_, _12319_);
  and (_12323_, _03178_, \oc8051_golden_model_1.PC [1]);
  nor (_12324_, _12323_, _04512_);
  and (_12325_, _12324_, _12322_);
  and (_12326_, _05617_, _04303_);
  nor (_12327_, _12326_, _12207_);
  nor (_12328_, _12327_, _04511_);
  nor (_12329_, _12328_, _04513_);
  or (_12330_, _12329_, _12325_);
  nor (_12331_, _05617_, _03274_);
  and (_12332_, _05617_, _03274_);
  nor (_12333_, _12332_, _12331_);
  or (_12334_, _12333_, _05850_);
  and (_12335_, _12334_, _06383_);
  and (_12336_, _12335_, _12330_);
  or (_12337_, _12336_, _12208_);
  and (_12338_, _12337_, _06382_);
  and (_12339_, _12331_, _04514_);
  or (_12340_, _12339_, _03192_);
  or (_12341_, _12340_, _12338_);
  and (_12342_, _03192_, \oc8051_golden_model_1.PC [1]);
  nor (_12343_, _12342_, _06390_);
  and (_12344_, _12343_, _12341_);
  nor (_12345_, _12326_, _06395_);
  or (_12346_, _12345_, _06394_);
  or (_12347_, _12346_, _12344_);
  nand (_12348_, _12332_, _06394_);
  and (_12349_, _12348_, _06399_);
  and (_12350_, _12349_, _12347_);
  and (_12351_, _03188_, _02878_);
  or (_12352_, _03972_, _12351_);
  or (_12353_, _12352_, _12350_);
  and (_12354_, _12353_, _12206_);
  or (_12355_, _12354_, _03491_);
  and (_12356_, _12205_, _03491_);
  nor (_12357_, _12356_, _04322_);
  and (_12358_, _12357_, _12355_);
  nand (_12359_, _12205_, _03027_);
  and (_12360_, _12359_, _04803_);
  or (_12361_, _12360_, _12358_);
  nand (_12362_, _12205_, _03495_);
  and (_12363_, _12362_, _06409_);
  and (_12364_, _12363_, _12361_);
  nor (_12365_, _12203_, _06409_);
  or (_12366_, _12365_, _04531_);
  or (_12367_, _12366_, _12364_);
  nand (_12368_, _12213_, _04531_);
  and (_12369_, _12368_, _12367_);
  or (_12370_, _12369_, _03629_);
  not (_12371_, _03198_);
  nand (_12372_, _03629_, _11442_);
  and (_12373_, _12372_, _12371_);
  and (_12374_, _12373_, _12370_);
  and (_12375_, _03198_, _02878_);
  or (_12376_, _04539_, _12375_);
  or (_12377_, _12376_, _12374_);
  or (_12378_, _12254_, _04558_);
  and (_12379_, _12378_, _11955_);
  and (_12380_, _12379_, _12377_);
  and (_12381_, _12205_, _11956_);
  or (_12382_, _12381_, _04552_);
  or (_12383_, _12382_, _12380_);
  and (_12384_, _12383_, _12204_);
  or (_12385_, _12384_, _03448_);
  or (_12386_, _12213_, _04713_);
  and (_12387_, _12386_, _04796_);
  and (_12388_, _12387_, _12385_);
  or (_12389_, _12388_, _11999_);
  and (_12390_, _12389_, _12202_);
  nor (_12391_, _11543_, _03629_);
  and (_12392_, _11408_, _03629_);
  or (_12393_, _12392_, _12391_);
  and (_12394_, _12393_, _12195_);
  or (_40635_, _12394_, _12390_);
  or (_12395_, _12183_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_12396_, _12395_, _12200_);
  not (_12397_, _12183_);
  nor (_12398_, _06765_, _07849_);
  nor (_12399_, _12398_, _07850_);
  and (_12400_, _12399_, _11956_);
  not (_12401_, _06637_);
  and (_12402_, _06547_, _12401_);
  nor (_12403_, _06547_, _12401_);
  or (_12404_, _12403_, _12402_);
  and (_12405_, _12404_, _04242_);
  and (_12406_, _03210_, _03188_);
  nor (_12407_, _05717_, _03946_);
  and (_12408_, _12407_, _04515_);
  nor (_12409_, _10083_, _05302_);
  or (_12410_, _12409_, _05940_);
  nand (_12411_, _10083_, _09670_);
  or (_12412_, _12411_, _05954_);
  and (_12413_, _05717_, _05617_);
  and (_12414_, _12413_, _05956_);
  nor (_12415_, _05957_, _05717_);
  nor (_12416_, _12415_, _12414_);
  nor (_12417_, _12416_, _06071_);
  and (_12418_, _05835_, _04875_);
  nor (_12419_, _05835_, _04875_);
  or (_12420_, _12419_, _12418_);
  or (_12421_, _12420_, _06072_);
  and (_12422_, _03980_, _03210_);
  nor (_12423_, _03980_, _07584_);
  or (_12424_, _12423_, _12422_);
  nor (_12425_, _12424_, _06073_);
  nor (_12426_, _12425_, _04421_);
  and (_12427_, _12426_, _12421_);
  or (_12428_, _12427_, _04428_);
  or (_12429_, _12428_, _12417_);
  and (_12430_, _12429_, _12412_);
  or (_12431_, _12430_, _04768_);
  nor (_12432_, _03210_, _03230_);
  nor (_12433_, _12432_, _04431_);
  and (_12434_, _12433_, _12431_);
  and (_12435_, _07849_, _04431_);
  or (_12436_, _12435_, _04449_);
  or (_12437_, _12436_, _12434_);
  and (_12438_, _12437_, _12410_);
  or (_12439_, _12438_, _03508_);
  nand (_12440_, _08260_, _03508_);
  and (_12441_, _12440_, _04562_);
  and (_12442_, _12441_, _12439_);
  not (_12443_, _10084_);
  and (_12444_, _12411_, _12443_);
  and (_12445_, _12444_, _04454_);
  or (_12446_, _12445_, _12442_);
  and (_12447_, _12446_, _03227_);
  nor (_12448_, _03245_, _03227_);
  or (_12449_, _03745_, _12448_);
  or (_12450_, _12449_, _12447_);
  nand (_12451_, _08260_, _03745_);
  and (_12452_, _12451_, _12450_);
  or (_12453_, _12452_, _04463_);
  and (_12454_, _06637_, _03446_);
  nand (_12455_, _08259_, _04463_);
  or (_12456_, _12455_, _12454_);
  and (_12457_, _12456_, _12453_);
  or (_12458_, _12457_, _04462_);
  nor (_12459_, _09693_, _05302_);
  and (_12460_, _05302_, \oc8051_golden_model_1.PSW [7]);
  nor (_12461_, _12460_, _12459_);
  nand (_12462_, _12461_, _04462_);
  and (_12463_, _12462_, _05897_);
  and (_12464_, _12463_, _12458_);
  nand (_12465_, _03210_, _03224_);
  nand (_12466_, _04480_, _12465_);
  or (_12467_, _12466_, _12464_);
  or (_12468_, _07849_, _04480_);
  and (_12469_, _12468_, _12467_);
  or (_12470_, _12469_, _04482_);
  or (_12471_, _06637_, _06164_);
  and (_12472_, _12471_, _06163_);
  and (_12473_, _12472_, _12470_);
  nor (_12474_, _06171_, _04875_);
  and (_12475_, _06340_, \oc8051_golden_model_1.P1INREG [2]);
  not (_12476_, _12475_);
  and (_12477_, _06343_, \oc8051_golden_model_1.P0INREG [2]);
  not (_12478_, _12477_);
  and (_12479_, _06346_, \oc8051_golden_model_1.P2INREG [2]);
  and (_12480_, _06348_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_12481_, _12480_, _12479_);
  and (_12482_, _12481_, _12478_);
  and (_12483_, _12482_, _12476_);
  and (_12484_, _06284_, \oc8051_golden_model_1.TL0 [2]);
  and (_12485_, _06279_, \oc8051_golden_model_1.TMOD [2]);
  nor (_12486_, _12485_, _12484_);
  and (_12487_, _12486_, _12483_);
  and (_12488_, _06315_, \oc8051_golden_model_1.IE [2]);
  and (_12489_, _06319_, \oc8051_golden_model_1.SBUF [2]);
  and (_12490_, _06321_, \oc8051_golden_model_1.SCON [2]);
  or (_12491_, _12490_, _12489_);
  nor (_12492_, _12491_, _12488_);
  and (_12493_, _06272_, \oc8051_golden_model_1.DPH [2]);
  and (_12494_, _06288_, \oc8051_golden_model_1.TH1 [2]);
  nor (_12495_, _12494_, _12493_);
  and (_12496_, _12495_, _12492_);
  and (_12497_, _12496_, _12487_);
  and (_12498_, _06327_, \oc8051_golden_model_1.TH0 [2]);
  and (_12499_, _06329_, \oc8051_golden_model_1.TL1 [2]);
  nor (_12500_, _12499_, _12498_);
  and (_12501_, _06334_, \oc8051_golden_model_1.PCON [2]);
  and (_12502_, _06336_, \oc8051_golden_model_1.TCON [2]);
  nor (_12503_, _12502_, _12501_);
  and (_12504_, _12503_, _12500_);
  and (_12505_, _06296_, \oc8051_golden_model_1.IP [2]);
  and (_12506_, _06303_, \oc8051_golden_model_1.PSW [2]);
  nor (_12507_, _12506_, _12505_);
  and (_12508_, _06308_, \oc8051_golden_model_1.ACC [2]);
  and (_12509_, _06310_, \oc8051_golden_model_1.B [2]);
  nor (_12510_, _12509_, _12508_);
  and (_12511_, _12510_, _12507_);
  and (_12512_, _06354_, \oc8051_golden_model_1.SP [2]);
  and (_12513_, _06356_, \oc8051_golden_model_1.DPL [2]);
  nor (_12514_, _12513_, _12512_);
  and (_12515_, _12514_, _12511_);
  and (_12516_, _12515_, _12504_);
  and (_12517_, _12516_, _12497_);
  not (_12518_, _12517_);
  nor (_12519_, _12518_, _12474_);
  nor (_12520_, _12519_, _06170_);
  or (_12521_, _12520_, _06168_);
  or (_12522_, _12521_, _12473_);
  and (_12523_, _06168_, _03904_);
  nor (_12524_, _12523_, _04500_);
  and (_12525_, _12524_, _12522_);
  and (_12526_, _04500_, _06332_);
  or (_12527_, _12526_, _03178_);
  or (_12528_, _12527_, _12525_);
  and (_12529_, _03245_, _03178_);
  nor (_12530_, _12529_, _04512_);
  and (_12531_, _12530_, _12528_);
  and (_12532_, _05717_, _03946_);
  nor (_12533_, _12532_, _12407_);
  nor (_12534_, _12533_, _04511_);
  nor (_12535_, _12534_, _04513_);
  or (_12536_, _12535_, _12531_);
  nor (_12537_, _05717_, _07584_);
  and (_12538_, _05717_, _07584_);
  nor (_12539_, _12538_, _12537_);
  or (_12540_, _12539_, _05850_);
  and (_12541_, _12540_, _06383_);
  and (_12542_, _12541_, _12536_);
  or (_12543_, _12542_, _12408_);
  and (_12544_, _12543_, _06382_);
  and (_12545_, _12537_, _04514_);
  or (_12546_, _12545_, _03192_);
  or (_12547_, _12546_, _12544_);
  and (_12548_, _03245_, _03192_);
  nor (_12549_, _12548_, _06390_);
  and (_12550_, _12549_, _12547_);
  nor (_12551_, _12532_, _06395_);
  or (_12552_, _12551_, _06394_);
  or (_12553_, _12552_, _12550_);
  nand (_12554_, _12538_, _06394_);
  and (_12555_, _12554_, _06399_);
  and (_12556_, _12555_, _12553_);
  or (_12557_, _12556_, _12406_);
  and (_12558_, _12557_, _05848_);
  not (_12559_, _02994_);
  and (_12560_, _04533_, _12559_);
  not (_12561_, _05848_);
  and (_12562_, _12420_, _12561_);
  or (_12563_, _12562_, _12560_);
  or (_12564_, _12563_, _12558_);
  not (_12565_, _04242_);
  nand (_12566_, _04533_, _12559_);
  or (_12567_, _12566_, _12404_);
  and (_12568_, _12567_, _12565_);
  and (_12569_, _12568_, _12564_);
  or (_12570_, _12569_, _12405_);
  and (_12571_, _12570_, _06408_);
  nor (_12572_, _12416_, _06408_);
  or (_12573_, _12572_, _03629_);
  or (_12574_, _12573_, _12571_);
  nand (_12575_, _11440_, _03629_);
  and (_12576_, _12575_, _12371_);
  and (_12577_, _12576_, _12574_);
  and (_12578_, _03210_, _03198_);
  or (_12579_, _04539_, _12578_);
  or (_12580_, _12579_, _12577_);
  or (_12581_, _12459_, _04558_);
  and (_12582_, _12581_, _11955_);
  and (_12583_, _12582_, _12580_);
  or (_12584_, _12583_, _12400_);
  and (_12585_, _12584_, _06785_);
  or (_12586_, _06786_, _06637_);
  nor (_12587_, _08016_, _06785_);
  and (_12588_, _12587_, _12586_);
  or (_12589_, _12588_, _03448_);
  or (_12590_, _12589_, _12585_);
  nor (_12591_, _05718_, _05667_);
  nor (_12592_, _12591_, _05719_);
  or (_12593_, _12592_, _04713_);
  and (_12594_, _12593_, _12174_);
  and (_12595_, _12594_, _12590_);
  or (_12596_, _12595_, _12397_);
  and (_12597_, _12596_, _12396_);
  and (_12598_, _11394_, _03629_);
  and (_12599_, _11529_, _11944_);
  or (_12600_, _12599_, _12598_);
  and (_12601_, _12600_, _12195_);
  or (_40637_, _12601_, _12597_);
  or (_12602_, _12183_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_12603_, _12602_, _12200_);
  nor (_12604_, _12402_, _08636_);
  or (_12605_, _12604_, _06639_);
  and (_12606_, _12605_, _04533_);
  and (_12607_, _03297_, _03188_);
  nor (_12608_, _05566_, _03708_);
  and (_12609_, _12608_, _04515_);
  and (_12610_, _05296_, \oc8051_golden_model_1.PSW [7]);
  nor (_12611_, _09825_, _05296_);
  nor (_12612_, _12611_, _12610_);
  nor (_12613_, _12612_, _05063_);
  or (_12614_, _08636_, _03454_);
  nand (_12615_, _12614_, _08247_);
  and (_12616_, _12615_, _04463_);
  nor (_12617_, _12418_, _05005_);
  or (_12618_, _12617_, _05837_);
  or (_12619_, _12618_, _06072_);
  and (_12620_, _03980_, _03297_);
  nor (_12621_, _03980_, _07578_);
  or (_12622_, _12621_, _06073_);
  or (_12623_, _12622_, _12620_);
  and (_12624_, _12623_, _12619_);
  and (_12625_, _12624_, _06071_);
  nor (_12626_, _12414_, _05566_);
  nor (_12627_, _12626_, _05959_);
  nor (_12628_, _12627_, _06071_);
  or (_12629_, _12628_, _12625_);
  or (_12630_, _12629_, _04428_);
  nand (_12631_, _10146_, _09802_);
  or (_12632_, _12631_, _05954_);
  and (_12633_, _12632_, _12630_);
  or (_12634_, _12633_, _04768_);
  nor (_12635_, _03297_, _03230_);
  nor (_12636_, _12635_, _04431_);
  and (_12637_, _12636_, _12634_);
  and (_12638_, _07848_, _04431_);
  or (_12639_, _12638_, _04449_);
  or (_12640_, _12639_, _12637_);
  nor (_12641_, _10146_, _05296_);
  or (_12642_, _12641_, _05940_);
  and (_12643_, _12642_, _12640_);
  or (_12644_, _12643_, _03508_);
  nand (_12645_, _08248_, _03508_);
  and (_12646_, _12645_, _04562_);
  and (_12647_, _12646_, _12644_);
  not (_12648_, _10147_);
  and (_12649_, _12631_, _12648_);
  and (_12650_, _12649_, _04454_);
  or (_12651_, _12650_, _12647_);
  and (_12652_, _12651_, _03227_);
  nor (_12653_, _03648_, _03227_);
  or (_12654_, _03745_, _12653_);
  or (_12655_, _12654_, _12652_);
  nand (_12656_, _08248_, _03745_);
  and (_12657_, _12656_, _05976_);
  and (_12658_, _12657_, _12655_);
  or (_12659_, _12658_, _12616_);
  and (_12660_, _12659_, _05063_);
  or (_12661_, _12660_, _12613_);
  and (_12662_, _12661_, _05897_);
  nand (_12663_, _03297_, _03224_);
  nand (_12664_, _04480_, _12663_);
  or (_12665_, _12664_, _12662_);
  or (_12666_, _07848_, _04480_);
  and (_12667_, _12666_, _12665_);
  or (_12668_, _12667_, _04482_);
  or (_12669_, _06592_, _06164_);
  and (_12670_, _12669_, _06163_);
  and (_12671_, _12670_, _12668_);
  nor (_12672_, _06171_, _05005_);
  and (_12673_, _06356_, \oc8051_golden_model_1.DPL [3]);
  and (_12674_, _06284_, \oc8051_golden_model_1.TL0 [3]);
  nor (_12675_, _12674_, _12673_);
  and (_12676_, _06272_, \oc8051_golden_model_1.DPH [3]);
  and (_12677_, _06288_, \oc8051_golden_model_1.TH1 [3]);
  nor (_12678_, _12677_, _12676_);
  and (_12679_, _12678_, _12675_);
  and (_12680_, _06315_, \oc8051_golden_model_1.IE [3]);
  and (_12681_, _06319_, \oc8051_golden_model_1.SBUF [3]);
  and (_12682_, _06321_, \oc8051_golden_model_1.SCON [3]);
  or (_12683_, _12682_, _12681_);
  nor (_12684_, _12683_, _12680_);
  and (_12685_, _06296_, \oc8051_golden_model_1.IP [3]);
  and (_12686_, _06303_, \oc8051_golden_model_1.PSW [3]);
  nor (_12687_, _12686_, _12685_);
  and (_12688_, _06308_, \oc8051_golden_model_1.ACC [3]);
  and (_12689_, _06310_, \oc8051_golden_model_1.B [3]);
  nor (_12690_, _12689_, _12688_);
  and (_12691_, _12690_, _12687_);
  and (_12692_, _12691_, _12684_);
  and (_12693_, _12692_, _12679_);
  and (_12694_, _06327_, \oc8051_golden_model_1.TH0 [3]);
  and (_12695_, _06329_, \oc8051_golden_model_1.TL1 [3]);
  nor (_12696_, _12695_, _12694_);
  and (_12697_, _06334_, \oc8051_golden_model_1.PCON [3]);
  and (_12698_, _06336_, \oc8051_golden_model_1.TCON [3]);
  nor (_12699_, _12698_, _12697_);
  and (_12700_, _12699_, _12696_);
  and (_12701_, _06340_, \oc8051_golden_model_1.P1INREG [3]);
  not (_12703_, _12701_);
  and (_12704_, _06343_, \oc8051_golden_model_1.P0INREG [3]);
  not (_12705_, _12704_);
  and (_12706_, _06346_, \oc8051_golden_model_1.P2INREG [3]);
  and (_12707_, _06348_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_12708_, _12707_, _12706_);
  and (_12709_, _12708_, _12705_);
  and (_12710_, _12709_, _12703_);
  and (_12711_, _06354_, \oc8051_golden_model_1.SP [3]);
  and (_12712_, _06279_, \oc8051_golden_model_1.TMOD [3]);
  nor (_12713_, _12712_, _12711_);
  and (_12714_, _12713_, _12710_);
  and (_12715_, _12714_, _12700_);
  and (_12716_, _12715_, _12693_);
  not (_12717_, _12716_);
  nor (_12718_, _12717_, _12672_);
  nor (_12719_, _12718_, _06170_);
  or (_12720_, _12719_, _06168_);
  or (_12721_, _12720_, _12671_);
  and (_12722_, _06168_, _03581_);
  nor (_12724_, _12722_, _04500_);
  and (_12725_, _12724_, _12721_);
  and (_12726_, _04500_, _06276_);
  or (_12727_, _12726_, _03178_);
  or (_12728_, _12727_, _12725_);
  and (_12729_, _03648_, _03178_);
  nor (_12730_, _12729_, _04512_);
  and (_12731_, _12730_, _12728_);
  and (_12732_, _05566_, _03708_);
  nor (_12733_, _12732_, _12608_);
  nor (_12734_, _12733_, _04511_);
  nor (_12735_, _12734_, _04513_);
  or (_12736_, _12735_, _12731_);
  nor (_12737_, _05566_, _07578_);
  and (_12738_, _05566_, _07578_);
  nor (_12739_, _12738_, _12737_);
  or (_12740_, _12739_, _05850_);
  and (_12741_, _12740_, _06383_);
  and (_12742_, _12741_, _12736_);
  or (_12743_, _12742_, _12609_);
  and (_12744_, _12743_, _06382_);
  and (_12745_, _12737_, _04514_);
  or (_12746_, _12745_, _03192_);
  or (_12747_, _12746_, _12744_);
  and (_12748_, _03648_, _03192_);
  nor (_12749_, _12748_, _06390_);
  and (_12750_, _12749_, _12747_);
  nor (_12751_, _12732_, _06395_);
  or (_12752_, _12751_, _06394_);
  or (_12753_, _12752_, _12750_);
  nand (_12754_, _12738_, _06394_);
  and (_12755_, _12754_, _06399_);
  and (_12756_, _12755_, _12753_);
  or (_12757_, _12756_, _12607_);
  and (_12758_, _12757_, _05847_);
  not (_12759_, _05847_);
  and (_12760_, _12618_, _12759_);
  or (_12761_, _12760_, _03495_);
  or (_12762_, _12761_, _12758_);
  or (_12763_, _12618_, _04745_);
  and (_12764_, _12763_, _06409_);
  and (_12765_, _12764_, _12762_);
  or (_12766_, _12765_, _12606_);
  and (_12767_, _12766_, _06408_);
  nor (_12768_, _12627_, _06408_);
  or (_12769_, _12768_, _03629_);
  or (_12770_, _12769_, _12767_);
  nand (_12771_, _11435_, _03629_);
  and (_12772_, _12771_, _12371_);
  and (_12773_, _12772_, _12770_);
  and (_12774_, _03297_, _03198_);
  or (_12775_, _04539_, _12774_);
  or (_12776_, _12775_, _12773_);
  or (_12777_, _12611_, _04558_);
  and (_12778_, _12777_, _06757_);
  and (_12779_, _12778_, _12776_);
  nor (_12780_, _07850_, _07848_);
  nor (_12781_, _12780_, _06767_);
  and (_12782_, _12781_, _06758_);
  or (_12783_, _12782_, _04547_);
  or (_12784_, _12783_, _12779_);
  or (_12785_, _12781_, _06780_);
  and (_12786_, _12785_, _06785_);
  and (_12787_, _12786_, _12784_);
  or (_12788_, _08016_, _06592_);
  nor (_12789_, _06788_, _06785_);
  and (_12790_, _12789_, _12788_);
  or (_12791_, _12790_, _03448_);
  or (_12792_, _12791_, _12787_);
  nor (_12793_, _05719_, _05567_);
  nor (_12794_, _12793_, _05720_);
  or (_12795_, _12794_, _04713_);
  and (_12796_, _12795_, _12174_);
  and (_12797_, _12796_, _12792_);
  or (_12798_, _12797_, _12397_);
  and (_12799_, _12798_, _12603_);
  nor (_12800_, _11534_, _03629_);
  and (_12801_, _11399_, _03629_);
  or (_12802_, _12801_, _12800_);
  and (_12803_, _12802_, _12195_);
  or (_40638_, _12803_, _12799_);
  or (_12804_, _12183_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_12805_, _12804_, _12200_);
  not (_12806_, _06730_);
  and (_12807_, _06639_, _12806_);
  nor (_12808_, _06639_, _12806_);
  or (_12809_, _12808_, _12807_);
  and (_12810_, _12809_, _04533_);
  nor (_12811_, _05837_, _05777_);
  and (_12812_, _05837_, _05777_);
  or (_12813_, _12812_, _12811_);
  or (_12814_, _12813_, _05847_);
  nor (_12815_, _05824_, _07484_);
  and (_12816_, _05824_, _07484_);
  nor (_12817_, _12816_, _12815_);
  and (_12818_, _12817_, _04511_);
  and (_12819_, _06236_, _05824_);
  nor (_12820_, _06236_, _05824_);
  nor (_12821_, _12820_, _12819_);
  and (_12822_, _12821_, _04512_);
  nor (_12823_, _09745_, _09721_);
  and (_12824_, _09721_, \oc8051_golden_model_1.PSW [7]);
  nor (_12825_, _12824_, _12823_);
  nor (_12826_, _12825_, _05063_);
  nor (_12827_, _09721_, _10109_);
  or (_12828_, _12827_, _05940_);
  and (_12829_, _11564_, _03980_);
  nor (_12830_, _03980_, _07484_);
  or (_12831_, _12830_, _12829_);
  and (_12832_, _12831_, _06072_);
  and (_12833_, _12813_, _06073_);
  or (_12834_, _12833_, _12832_);
  and (_12835_, _12834_, _05966_);
  and (_12836_, _06730_, _04422_);
  or (_12837_, _12836_, _12835_);
  and (_12838_, _12837_, _06071_);
  and (_12839_, _05959_, _05824_);
  nor (_12840_, _05959_, _05824_);
  nor (_12841_, _12840_, _12839_);
  nor (_12842_, _12841_, _06071_);
  or (_12843_, _12842_, _12838_);
  and (_12844_, _12843_, _05954_);
  nand (_12845_, _09722_, _10109_);
  and (_12846_, _12845_, _04428_);
  or (_12847_, _12846_, _04768_);
  or (_12848_, _12847_, _12844_);
  nor (_12849_, _11564_, _03230_);
  nor (_12850_, _12849_, _04431_);
  and (_12851_, _12850_, _12848_);
  and (_12852_, _06763_, _04431_);
  or (_12853_, _12852_, _04449_);
  or (_12854_, _12853_, _12851_);
  and (_12855_, _12854_, _12828_);
  or (_12856_, _12855_, _03508_);
  nand (_12857_, _08235_, _03508_);
  and (_12858_, _12857_, _04562_);
  and (_12859_, _12858_, _12856_);
  not (_12860_, _10110_);
  and (_12861_, _12845_, _12860_);
  and (_12862_, _12861_, _04454_);
  or (_12863_, _12862_, _12859_);
  and (_12864_, _12863_, _03227_);
  nor (_12865_, _11565_, _03227_);
  or (_12866_, _12865_, _03745_);
  or (_12867_, _12866_, _12864_);
  nand (_12868_, _08235_, _03745_);
  and (_12869_, _12868_, _12867_);
  or (_12870_, _12869_, _04463_);
  and (_12871_, _06730_, _03446_);
  nand (_12872_, _08234_, _04463_);
  or (_12873_, _12872_, _12871_);
  and (_12874_, _12873_, _05063_);
  and (_12875_, _12874_, _12870_);
  or (_12876_, _12875_, _12826_);
  and (_12877_, _12876_, _05897_);
  nand (_12878_, _11564_, _03224_);
  nand (_12879_, _12878_, _04480_);
  or (_12880_, _12879_, _12877_);
  or (_12881_, _06763_, _04480_);
  and (_12882_, _12881_, _12880_);
  or (_12883_, _12882_, _04482_);
  or (_12884_, _06730_, _06164_);
  and (_12885_, _12884_, _06163_);
  and (_12886_, _12885_, _12883_);
  nor (_12887_, _06171_, _05777_);
  and (_12888_, _06340_, \oc8051_golden_model_1.P1INREG [4]);
  not (_12889_, _12888_);
  and (_12890_, _06343_, \oc8051_golden_model_1.P0INREG [4]);
  not (_12891_, _12890_);
  and (_12892_, _06346_, \oc8051_golden_model_1.P2INREG [4]);
  and (_12893_, _06348_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_12894_, _12893_, _12892_);
  and (_12895_, _12894_, _12891_);
  and (_12896_, _12895_, _12889_);
  and (_12897_, _06354_, \oc8051_golden_model_1.SP [4]);
  and (_12898_, _06284_, \oc8051_golden_model_1.TL0 [4]);
  nor (_12899_, _12898_, _12897_);
  and (_12900_, _12899_, _12896_);
  and (_12901_, _06315_, \oc8051_golden_model_1.IE [4]);
  and (_12902_, _06319_, \oc8051_golden_model_1.SBUF [4]);
  and (_12903_, _06321_, \oc8051_golden_model_1.SCON [4]);
  or (_12904_, _12903_, _12902_);
  nor (_12905_, _12904_, _12901_);
  and (_12906_, _06296_, \oc8051_golden_model_1.IP [4]);
  and (_12907_, _06310_, \oc8051_golden_model_1.B [4]);
  nor (_12908_, _12907_, _12906_);
  and (_12909_, _06303_, \oc8051_golden_model_1.PSW [4]);
  and (_12910_, _06308_, \oc8051_golden_model_1.ACC [4]);
  nor (_12911_, _12910_, _12909_);
  and (_12912_, _12911_, _12908_);
  and (_12913_, _12912_, _12905_);
  and (_12914_, _12913_, _12900_);
  and (_12915_, _06272_, \oc8051_golden_model_1.DPH [4]);
  and (_12916_, _06279_, \oc8051_golden_model_1.TMOD [4]);
  nor (_12917_, _12916_, _12915_);
  and (_12918_, _06356_, \oc8051_golden_model_1.DPL [4]);
  and (_12919_, _06288_, \oc8051_golden_model_1.TH1 [4]);
  nor (_12920_, _12919_, _12918_);
  and (_12921_, _12920_, _12917_);
  and (_12922_, _06293_, _06269_);
  and (_12923_, _12922_, \oc8051_golden_model_1.TCON [4]);
  and (_12924_, _06327_, \oc8051_golden_model_1.TH0 [4]);
  nor (_12925_, _12924_, _12923_);
  and (_12926_, _06334_, \oc8051_golden_model_1.PCON [4]);
  and (_12927_, _06329_, \oc8051_golden_model_1.TL1 [4]);
  nor (_12928_, _12927_, _12926_);
  and (_12929_, _12928_, _12925_);
  and (_12930_, _12929_, _12921_);
  and (_12931_, _12930_, _12914_);
  not (_12932_, _12931_);
  nor (_12933_, _12932_, _12887_);
  nor (_12934_, _12933_, _06170_);
  or (_12935_, _12934_, _06168_);
  or (_12936_, _12935_, _12886_);
  and (_12937_, _06168_, _03486_);
  nor (_12938_, _12937_, _04500_);
  and (_12939_, _12938_, _12936_);
  and (_12940_, _06298_, _04500_);
  or (_12941_, _12940_, _03178_);
  or (_12942_, _12941_, _12939_);
  and (_12943_, _11565_, _03178_);
  nor (_12944_, _12943_, _04512_);
  and (_12945_, _12944_, _12942_);
  or (_12946_, _12945_, _12822_);
  and (_12947_, _12946_, _05850_);
  or (_12948_, _12947_, _12818_);
  and (_12949_, _12948_, _06383_);
  and (_12950_, _12820_, _04515_);
  or (_12951_, _12950_, _12949_);
  and (_12952_, _12951_, _06382_);
  and (_12953_, _12815_, _04514_);
  or (_12954_, _12953_, _03192_);
  or (_12955_, _12954_, _12952_);
  and (_12956_, _11565_, _03192_);
  nor (_12957_, _12956_, _06390_);
  and (_12958_, _12957_, _12955_);
  nor (_12959_, _12819_, _06395_);
  or (_12960_, _12959_, _06394_);
  or (_12961_, _12960_, _12958_);
  nand (_12962_, _12816_, _06394_);
  and (_12963_, _12962_, _06399_);
  and (_12964_, _12963_, _12961_);
  nand (_12965_, _11564_, _03188_);
  nand (_12966_, _12965_, _05847_);
  or (_12967_, _12966_, _12964_);
  and (_12968_, _12967_, _12814_);
  or (_12969_, _12968_, _03495_);
  or (_12970_, _12813_, _04745_);
  and (_12971_, _12970_, _06409_);
  and (_12972_, _12971_, _12969_);
  or (_12973_, _12972_, _12810_);
  and (_12974_, _12973_, _06408_);
  nor (_12975_, _12841_, _06408_);
  or (_12976_, _12975_, _03629_);
  or (_12977_, _12976_, _12974_);
  nand (_12978_, _11431_, _03629_);
  and (_12979_, _12978_, _12371_);
  and (_12980_, _12979_, _12977_);
  and (_12981_, _11564_, _03198_);
  or (_12982_, _12981_, _04539_);
  or (_12983_, _12982_, _12980_);
  or (_12984_, _12823_, _04558_);
  and (_12985_, _12984_, _11955_);
  and (_12986_, _12985_, _12983_);
  and (_12987_, _03616_, _03195_);
  or (_12988_, _06767_, _06763_);
  nor (_12989_, _11955_, _06768_);
  and (_12990_, _12989_, _12988_);
  or (_12991_, _12990_, _12987_);
  or (_12992_, _12991_, _12986_);
  not (_12993_, _12987_);
  nor (_12994_, _06788_, _06730_);
  nor (_12995_, _12994_, _07999_);
  nor (_12996_, _12995_, _12993_);
  nor (_12997_, _12996_, _04256_);
  and (_12998_, _12997_, _12992_);
  and (_12999_, _12995_, _04256_);
  or (_13000_, _12999_, _03448_);
  or (_13001_, _13000_, _12998_);
  nor (_13002_, _05825_, _05720_);
  nor (_13003_, _13002_, _05826_);
  or (_13004_, _13003_, _04713_);
  and (_13005_, _13004_, _12174_);
  and (_13006_, _13005_, _13001_);
  or (_13007_, _13006_, _12397_);
  and (_13008_, _13007_, _12805_);
  and (_13009_, _11390_, _03629_);
  nor (_13010_, _11526_, _03629_);
  or (_13011_, _13010_, _13009_);
  and (_13012_, _13011_, _12195_);
  or (_40640_, _13012_, _13008_);
  nor (_13013_, _12839_, _05517_);
  nor (_13014_, _13013_, _05960_);
  nand (_13015_, _13014_, _04531_);
  nor (_13016_, _06267_, _05517_);
  and (_13017_, _13016_, _04515_);
  nor (_13018_, _09850_, _09827_);
  and (_13019_, _09827_, \oc8051_golden_model_1.PSW [7]);
  nor (_13020_, _13019_, _13018_);
  nor (_13021_, _13020_, _05063_);
  nor (_13022_, _12812_, _05469_);
  or (_13023_, _13022_, _05838_);
  and (_13024_, _13023_, _06073_);
  nor (_13025_, _03980_, _07478_);
  and (_13026_, _11559_, _03980_);
  or (_13027_, _13026_, _13025_);
  and (_13028_, _13027_, _06072_);
  or (_13029_, _13028_, _13024_);
  and (_13030_, _13029_, _05966_);
  and (_13031_, _06684_, _04422_);
  or (_13032_, _13031_, _13030_);
  and (_13033_, _13032_, _06071_);
  nor (_13034_, _13014_, _06071_);
  or (_13035_, _13034_, _13033_);
  and (_13036_, _13035_, _05954_);
  nand (_13037_, _09828_, _10158_);
  and (_13038_, _13037_, _04428_);
  or (_13039_, _13038_, _04768_);
  or (_13040_, _13039_, _13036_);
  nor (_13041_, _11559_, _03230_);
  nor (_13042_, _13041_, _04431_);
  and (_13043_, _13042_, _13040_);
  and (_13044_, _06762_, _04431_);
  or (_13045_, _13044_, _04449_);
  or (_13046_, _13045_, _13043_);
  nor (_13047_, _09827_, _10158_);
  or (_13048_, _13047_, _05940_);
  and (_13049_, _13048_, _13046_);
  or (_13050_, _13049_, _03508_);
  nand (_13051_, _08218_, _03508_);
  and (_13052_, _13051_, _04562_);
  and (_13053_, _13052_, _13050_);
  not (_13054_, _10159_);
  and (_13055_, _13037_, _13054_);
  and (_13056_, _13055_, _04454_);
  or (_13057_, _13056_, _13053_);
  and (_13058_, _13057_, _03227_);
  nor (_13059_, _11560_, _03227_);
  or (_13060_, _13059_, _03745_);
  or (_13061_, _13060_, _13058_);
  nand (_13062_, _08218_, _03745_);
  and (_13063_, _13062_, _13061_);
  or (_13064_, _13063_, _04463_);
  and (_13065_, _06684_, _03446_);
  nand (_13066_, _08217_, _04463_);
  or (_13067_, _13066_, _13065_);
  and (_13068_, _13067_, _05063_);
  and (_13069_, _13068_, _13064_);
  or (_13070_, _13069_, _13021_);
  and (_13071_, _13070_, _05897_);
  nand (_13072_, _11559_, _03224_);
  nand (_13073_, _13072_, _04480_);
  or (_13074_, _13073_, _13071_);
  or (_13075_, _06762_, _04480_);
  and (_13076_, _13075_, _13074_);
  or (_13077_, _13076_, _04482_);
  or (_13078_, _06684_, _06164_);
  and (_13079_, _13078_, _06163_);
  and (_13080_, _13079_, _13077_);
  nor (_13081_, _06171_, _05469_);
  and (_13082_, _06296_, \oc8051_golden_model_1.IP [5]);
  and (_13083_, _06310_, \oc8051_golden_model_1.B [5]);
  nor (_13084_, _13083_, _13082_);
  and (_13085_, _06303_, \oc8051_golden_model_1.PSW [5]);
  and (_13086_, _06308_, \oc8051_golden_model_1.ACC [5]);
  nor (_13087_, _13086_, _13085_);
  and (_13088_, _13087_, _13084_);
  and (_13089_, _06288_, \oc8051_golden_model_1.TH1 [5]);
  not (_13090_, _13089_);
  and (_13091_, _06354_, \oc8051_golden_model_1.SP [5]);
  and (_13092_, _06284_, \oc8051_golden_model_1.TL0 [5]);
  nor (_13093_, _13092_, _13091_);
  and (_13094_, _13093_, _13090_);
  and (_13095_, _13094_, _13088_);
  and (_13096_, _06327_, \oc8051_golden_model_1.TH0 [5]);
  and (_13097_, _06329_, \oc8051_golden_model_1.TL1 [5]);
  nor (_13098_, _13097_, _13096_);
  and (_13099_, _06334_, \oc8051_golden_model_1.PCON [5]);
  and (_13100_, _06336_, \oc8051_golden_model_1.TCON [5]);
  nor (_13101_, _13100_, _13099_);
  and (_13102_, _13101_, _13098_);
  and (_13103_, _06356_, \oc8051_golden_model_1.DPL [5]);
  not (_13104_, _13103_);
  and (_13105_, _06343_, \oc8051_golden_model_1.P0INREG [5]);
  not (_13106_, _13105_);
  and (_13107_, _06348_, \oc8051_golden_model_1.P3INREG [5]);
  and (_13108_, _06340_, \oc8051_golden_model_1.P1INREG [5]);
  and (_13109_, _06346_, \oc8051_golden_model_1.P2INREG [5]);
  or (_13110_, _13109_, _13108_);
  nor (_13111_, _13110_, _13107_);
  and (_13112_, _13111_, _13106_);
  and (_13113_, _13112_, _13104_);
  and (_13114_, _06315_, \oc8051_golden_model_1.IE [5]);
  and (_13115_, _06319_, \oc8051_golden_model_1.SBUF [5]);
  and (_13116_, _06321_, \oc8051_golden_model_1.SCON [5]);
  or (_13117_, _13116_, _13115_);
  nor (_13118_, _13117_, _13114_);
  and (_13119_, _06272_, \oc8051_golden_model_1.DPH [5]);
  and (_13120_, _06279_, \oc8051_golden_model_1.TMOD [5]);
  nor (_13121_, _13120_, _13119_);
  and (_13122_, _13121_, _13118_);
  and (_13123_, _13122_, _13113_);
  and (_13124_, _13123_, _13102_);
  and (_13125_, _13124_, _13095_);
  not (_13126_, _13125_);
  nor (_13127_, _13126_, _13081_);
  nor (_13128_, _13127_, _06170_);
  or (_13129_, _13128_, _06168_);
  or (_13130_, _13129_, _13080_);
  and (_13131_, _06168_, _03860_);
  nor (_13132_, _13131_, _04500_);
  and (_13133_, _13132_, _13130_);
  and (_13134_, _06306_, _04500_);
  or (_13135_, _13134_, _03178_);
  or (_13136_, _13135_, _13133_);
  and (_13137_, _11560_, _03178_);
  nor (_13138_, _13137_, _04512_);
  and (_13139_, _13138_, _13136_);
  and (_13140_, _06267_, _05517_);
  nor (_13141_, _13140_, _13016_);
  nor (_13142_, _13141_, _04511_);
  nor (_13143_, _13142_, _04513_);
  or (_13144_, _13143_, _13139_);
  nor (_13145_, _05517_, _07478_);
  and (_13146_, _05517_, _07478_);
  nor (_13147_, _13146_, _13145_);
  or (_13148_, _13147_, _05850_);
  and (_13149_, _13148_, _06383_);
  and (_13150_, _13149_, _13144_);
  or (_13151_, _13150_, _13017_);
  and (_13152_, _13151_, _06382_);
  and (_13153_, _13145_, _04514_);
  or (_13154_, _13153_, _03192_);
  or (_13155_, _13154_, _13152_);
  and (_13156_, _11560_, _03192_);
  nor (_13157_, _13156_, _06390_);
  and (_13158_, _13157_, _13155_);
  nor (_13159_, _13140_, _06395_);
  or (_13160_, _13159_, _06394_);
  or (_13161_, _13160_, _13158_);
  nand (_13162_, _13146_, _06394_);
  and (_13163_, _13162_, _06399_);
  and (_13164_, _13163_, _13161_);
  nand (_13165_, _11559_, _03188_);
  nand (_13166_, _13165_, _05848_);
  or (_13167_, _13166_, _13164_);
  and (_13168_, _13023_, _06409_);
  or (_13169_, _13168_, _11933_);
  and (_13170_, _13169_, _13167_);
  not (_13171_, _06684_);
  nor (_13172_, _12807_, _13171_);
  or (_13173_, _13172_, _06732_);
  and (_13174_, _13173_, _04533_);
  or (_13175_, _13174_, _04531_);
  or (_13176_, _13175_, _13170_);
  and (_13177_, _13176_, _13015_);
  or (_13178_, _13177_, _03629_);
  nand (_13179_, _11426_, _03629_);
  and (_13180_, _13179_, _12371_);
  and (_13181_, _13180_, _13178_);
  and (_13182_, _11559_, _03198_);
  or (_13183_, _13182_, _04539_);
  or (_13184_, _13183_, _13181_);
  or (_13185_, _13018_, _04558_);
  and (_13186_, _13185_, _11955_);
  and (_13187_, _13186_, _13184_);
  nor (_13188_, _06768_, _06762_);
  or (_13189_, _13188_, _06769_);
  nor (_13190_, _13189_, _11955_);
  or (_13191_, _13190_, _04552_);
  or (_13192_, _13191_, _13187_);
  nor (_13193_, _07999_, _06684_);
  nor (_13194_, _13193_, _06790_);
  or (_13195_, _13194_, _06785_);
  and (_13196_, _13195_, _13192_);
  or (_13197_, _13196_, _03448_);
  nor (_13198_, _05826_, _05518_);
  nor (_13199_, _13198_, _05827_);
  or (_13200_, _13199_, _04713_);
  and (_13201_, _13200_, _04796_);
  and (_13202_, _13201_, _13197_);
  or (_13203_, _13202_, _11999_);
  or (_13204_, _11998_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_13205_, _13204_, _12188_);
  and (_13206_, _13205_, _13203_);
  and (_13207_, _11385_, _03629_);
  and (_13208_, _11521_, _11944_);
  or (_13209_, _13208_, _13207_);
  and (_13210_, _13209_, _12195_);
  or (_40641_, _13210_, _13206_);
  or (_13211_, _12183_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_13212_, _13211_, _12200_);
  nor (_13213_, _06790_, _06455_);
  nor (_13214_, _13213_, _06791_);
  or (_13215_, _13214_, _06785_);
  nor (_13216_, _06732_, _06456_);
  or (_13217_, _13216_, _06733_);
  and (_13218_, _13217_, _04533_);
  nor (_13219_, _05838_, _05363_);
  or (_13220_, _13219_, _05839_);
  or (_13221_, _13220_, _05847_);
  nor (_13222_, _06204_, _05411_);
  and (_13223_, _13222_, _04515_);
  nor (_13224_, _09799_, _09775_);
  and (_13225_, _09775_, \oc8051_golden_model_1.PSW [7]);
  nor (_13226_, _13225_, _13224_);
  nor (_13227_, _13226_, _05063_);
  and (_13228_, _07818_, _04431_);
  nand (_13229_, _09776_, _10133_);
  or (_13230_, _13229_, _05954_);
  or (_13231_, _13220_, _06072_);
  and (_13232_, _11551_, _03980_);
  nor (_13233_, _03980_, _07433_);
  or (_13234_, _13233_, _06073_);
  or (_13235_, _13234_, _13232_);
  and (_13236_, _13235_, _13231_);
  or (_13237_, _13236_, _04422_);
  or (_13238_, _06455_, _05966_);
  and (_13239_, _13238_, _13237_);
  or (_13240_, _13239_, _04421_);
  nor (_13241_, _05960_, _05411_);
  nor (_13242_, _13241_, _05961_);
  nand (_13243_, _13242_, _04421_);
  and (_13244_, _13243_, _13240_);
  or (_13245_, _13244_, _04428_);
  and (_13246_, _13245_, _13230_);
  or (_13247_, _13246_, _04768_);
  nor (_13248_, _11551_, _03230_);
  nor (_13249_, _13248_, _04431_);
  and (_13250_, _13249_, _13247_);
  or (_13251_, _13250_, _13228_);
  and (_13252_, _13251_, _05940_);
  nor (_13253_, _09775_, _10133_);
  and (_13254_, _13253_, _04449_);
  or (_13255_, _13254_, _03508_);
  or (_13256_, _13255_, _13252_);
  nand (_13257_, _08203_, _03508_);
  and (_13258_, _13257_, _04562_);
  and (_13259_, _13258_, _13256_);
  not (_13260_, _10134_);
  and (_13261_, _13229_, _13260_);
  and (_13262_, _13261_, _04454_);
  or (_13263_, _13262_, _13259_);
  and (_13264_, _13263_, _03227_);
  nor (_13265_, _11552_, _03227_);
  or (_13266_, _13265_, _03745_);
  or (_13267_, _13266_, _13264_);
  nand (_13268_, _08203_, _03745_);
  and (_13269_, _13268_, _13267_);
  or (_13270_, _13269_, _04463_);
  and (_13271_, _06455_, _03446_);
  nand (_13272_, _08202_, _04463_);
  or (_13273_, _13272_, _13271_);
  and (_13274_, _13273_, _05063_);
  and (_13275_, _13274_, _13270_);
  or (_13276_, _13275_, _13227_);
  and (_13277_, _13276_, _05897_);
  nand (_13278_, _11551_, _03224_);
  nand (_13279_, _13278_, _04480_);
  or (_13280_, _13279_, _13277_);
  or (_13281_, _07818_, _04480_);
  and (_13282_, _13281_, _13280_);
  or (_13283_, _13282_, _04482_);
  or (_13284_, _06455_, _06164_);
  and (_13285_, _13284_, _06163_);
  and (_13286_, _13285_, _13283_);
  nor (_13287_, _06171_, _05363_);
  and (_13288_, _06272_, \oc8051_golden_model_1.DPH [6]);
  and (_13289_, _06288_, \oc8051_golden_model_1.TH1 [6]);
  nor (_13290_, _13289_, _13288_);
  and (_13291_, _06340_, \oc8051_golden_model_1.P1INREG [6]);
  not (_13292_, _13291_);
  and (_13293_, _06343_, \oc8051_golden_model_1.P0INREG [6]);
  not (_13294_, _13293_);
  and (_13295_, _06346_, \oc8051_golden_model_1.P2INREG [6]);
  and (_13296_, _06348_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_13297_, _13296_, _13295_);
  and (_13298_, _13297_, _13294_);
  and (_13299_, _13298_, _13292_);
  and (_13300_, _13299_, _13290_);
  and (_13301_, _06315_, \oc8051_golden_model_1.IE [6]);
  and (_13302_, _06319_, \oc8051_golden_model_1.SBUF [6]);
  and (_13303_, _06321_, \oc8051_golden_model_1.SCON [6]);
  or (_13304_, _13303_, _13302_);
  nor (_13305_, _13304_, _13301_);
  and (_13306_, _06296_, \oc8051_golden_model_1.IP [6]);
  and (_13307_, _06310_, \oc8051_golden_model_1.B [6]);
  nor (_13308_, _13307_, _13306_);
  and (_13309_, _06303_, \oc8051_golden_model_1.PSW [6]);
  and (_13310_, _06308_, \oc8051_golden_model_1.ACC [6]);
  nor (_13311_, _13310_, _13309_);
  and (_13312_, _13311_, _13308_);
  and (_13313_, _13312_, _13305_);
  and (_13314_, _13313_, _13300_);
  and (_13315_, _06327_, \oc8051_golden_model_1.TH0 [6]);
  and (_13316_, _06329_, \oc8051_golden_model_1.TL1 [6]);
  nor (_13317_, _13316_, _13315_);
  and (_13318_, _06334_, \oc8051_golden_model_1.PCON [6]);
  and (_13319_, _06336_, \oc8051_golden_model_1.TCON [6]);
  nor (_13320_, _13319_, _13318_);
  and (_13321_, _13320_, _13317_);
  and (_13322_, _06354_, \oc8051_golden_model_1.SP [6]);
  and (_13323_, _06356_, \oc8051_golden_model_1.DPL [6]);
  nor (_13324_, _13323_, _13322_);
  and (_13325_, _06284_, \oc8051_golden_model_1.TL0 [6]);
  and (_13326_, _06279_, \oc8051_golden_model_1.TMOD [6]);
  nor (_13327_, _13326_, _13325_);
  and (_13328_, _13327_, _13324_);
  and (_13329_, _13328_, _13321_);
  and (_13330_, _13329_, _13314_);
  not (_13331_, _13330_);
  nor (_13332_, _13331_, _13287_);
  nor (_13333_, _13332_, _06170_);
  or (_13334_, _13333_, _06168_);
  or (_13335_, _13334_, _13286_);
  and (_13336_, _06168_, _03549_);
  nor (_13337_, _13336_, _04500_);
  and (_13338_, _13337_, _13335_);
  not (_13339_, _06204_);
  and (_13340_, _13339_, _04500_);
  or (_13341_, _13340_, _03178_);
  or (_13342_, _13341_, _13338_);
  and (_13343_, _11552_, _03178_);
  nor (_13344_, _13343_, _04512_);
  and (_13345_, _13344_, _13342_);
  and (_13346_, _06204_, _05411_);
  nor (_13347_, _13346_, _13222_);
  nor (_13348_, _13347_, _04511_);
  nor (_13349_, _13348_, _04513_);
  or (_13350_, _13349_, _13345_);
  nor (_13351_, _05411_, _07433_);
  and (_13352_, _05411_, _07433_);
  nor (_13353_, _13352_, _13351_);
  or (_13354_, _13353_, _05850_);
  and (_13355_, _13354_, _06383_);
  and (_13356_, _13355_, _13350_);
  or (_13357_, _13356_, _13223_);
  and (_13358_, _13357_, _06382_);
  and (_13359_, _13351_, _04514_);
  or (_13360_, _13359_, _03192_);
  or (_13361_, _13360_, _13358_);
  and (_13362_, _11552_, _03192_);
  nor (_13363_, _13362_, _06390_);
  and (_13364_, _13363_, _13361_);
  nor (_13365_, _13346_, _06395_);
  or (_13366_, _13365_, _06394_);
  or (_13367_, _13366_, _13364_);
  nand (_13368_, _13352_, _06394_);
  and (_13369_, _13368_, _06399_);
  and (_13370_, _13369_, _13367_);
  nand (_13371_, _11551_, _03188_);
  nand (_13372_, _13371_, _05847_);
  or (_13373_, _13372_, _13370_);
  and (_13374_, _13373_, _13221_);
  or (_13375_, _13374_, _03495_);
  or (_13376_, _13220_, _04745_);
  and (_13377_, _13376_, _06409_);
  and (_13378_, _13377_, _13375_);
  or (_13379_, _13378_, _13218_);
  and (_13380_, _13379_, _06408_);
  nor (_13381_, _13242_, _06408_);
  or (_13382_, _13381_, _03629_);
  or (_13383_, _13382_, _13380_);
  nand (_13384_, _11418_, _03629_);
  and (_13385_, _13384_, _12371_);
  and (_13386_, _13385_, _13383_);
  and (_13387_, _11551_, _03198_);
  or (_13388_, _13387_, _04539_);
  or (_13389_, _13388_, _13386_);
  or (_13390_, _13224_, _04558_);
  and (_13391_, _13390_, _11955_);
  and (_13392_, _13391_, _13389_);
  nand (_13393_, _06769_, _07818_);
  or (_13394_, _06769_, _07818_);
  and (_13395_, _13394_, _11956_);
  and (_13396_, _13395_, _13393_);
  or (_13397_, _13396_, _04552_);
  or (_13398_, _13397_, _13392_);
  and (_13399_, _13398_, _13215_);
  or (_13400_, _13399_, _03448_);
  nor (_13401_, _05827_, _05412_);
  nor (_13402_, _13401_, _05828_);
  or (_13403_, _13402_, _04713_);
  and (_13404_, _13403_, _12174_);
  and (_13405_, _13404_, _13400_);
  or (_13406_, _13405_, _12397_);
  and (_13407_, _13406_, _13212_);
  and (_13408_, _11514_, _11944_);
  and (_13409_, _11378_, _03629_);
  or (_13410_, _13409_, _13408_);
  and (_13411_, _13410_, _12195_);
  or (_40642_, _13411_, _13407_);
  nor (_13412_, _12183_, _05144_);
  nor (_13413_, _12397_, _06799_);
  or (_13414_, _13413_, _13412_);
  and (_13415_, _13414_, _12200_);
  and (_13416_, _12195_, _06823_);
  or (_40644_, _13416_, _13415_);
  and (_13417_, _04798_, _04556_);
  and (_13418_, _13417_, _11996_);
  not (_13419_, _13418_);
  or (_13420_, _13419_, _12171_);
  or (_13421_, _13418_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand (_13422_, _12187_, _04804_);
  and (_13423_, _13422_, _13421_);
  and (_13424_, _13423_, _13420_);
  and (_13425_, _12194_, _04804_);
  and (_13426_, _13425_, _12198_);
  or (_40648_, _13426_, _13424_);
  not (_13427_, _13425_);
  or (_13428_, _13418_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_13429_, _13428_, _13427_);
  or (_13430_, _13419_, _12388_);
  and (_13431_, _13430_, _13429_);
  and (_13432_, _13425_, _12393_);
  or (_40649_, _13432_, _13431_);
  or (_13433_, _13418_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_13434_, _13433_, _13427_);
  and (_13435_, _12593_, _04796_);
  and (_13436_, _13435_, _12590_);
  or (_13437_, _13419_, _13436_);
  and (_13438_, _13437_, _13434_);
  and (_13439_, _13425_, _12600_);
  or (_40650_, _13439_, _13438_);
  or (_13440_, _13418_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_13441_, _13440_, _13427_);
  and (_13442_, _12795_, _04796_);
  and (_13443_, _13442_, _12792_);
  or (_13444_, _13419_, _13443_);
  and (_13445_, _13444_, _13441_);
  and (_13446_, _13425_, _12802_);
  or (_40651_, _13446_, _13445_);
  or (_13447_, _13418_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_13448_, _13447_, _13427_);
  and (_13449_, _13004_, _04796_);
  and (_13450_, _13449_, _13001_);
  or (_13451_, _13419_, _13450_);
  and (_13452_, _13451_, _13448_);
  and (_13453_, _13425_, _13011_);
  or (_40653_, _13453_, _13452_);
  or (_13454_, _13418_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_13455_, _13454_, _13427_);
  or (_13456_, _13419_, _13202_);
  and (_13457_, _13456_, _13455_);
  and (_13458_, _13425_, _13209_);
  or (_40654_, _13458_, _13457_);
  or (_13459_, _13418_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_13460_, _13459_, _13427_);
  and (_13461_, _13403_, _04796_);
  and (_13462_, _13461_, _13400_);
  or (_13463_, _13419_, _13462_);
  and (_13464_, _13463_, _13460_);
  and (_13465_, _13425_, _13410_);
  or (_40655_, _13465_, _13464_);
  or (_13466_, _13418_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_13467_, _13466_, _13427_);
  or (_13468_, _13419_, _06800_);
  and (_13469_, _13468_, _13467_);
  and (_13470_, _13425_, _06823_);
  or (_40656_, _13470_, _13469_);
  and (_13471_, _11993_, _04711_);
  and (_13472_, _13471_, _11996_);
  not (_13473_, _13472_);
  or (_13474_, _13473_, _12171_);
  and (_13475_, _12187_, _05967_);
  not (_13476_, _13475_);
  or (_13477_, _13472_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_13478_, _13477_, _13476_);
  and (_13479_, _13478_, _13474_);
  and (_13480_, _12198_, _05137_);
  and (_13481_, _13480_, _13475_);
  or (_40661_, _13481_, _13479_);
  or (_13482_, _13473_, _12388_);
  or (_13483_, _13472_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_13484_, _13483_, _13476_);
  and (_13485_, _13484_, _13482_);
  and (_13486_, _12393_, _05137_);
  and (_13487_, _13486_, _13475_);
  or (_40662_, _13487_, _13485_);
  and (_13488_, _12194_, _05967_);
  not (_13489_, _13488_);
  and (_13490_, _12179_, _04711_);
  and (_13491_, _13490_, _12178_);
  or (_13492_, _13491_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_13493_, _13492_, _13489_);
  not (_13494_, _13491_);
  or (_13495_, _13494_, _12595_);
  and (_13496_, _13495_, _13493_);
  and (_13497_, _12600_, _12191_);
  and (_13498_, _13497_, _13488_);
  or (_40663_, _13498_, _13496_);
  or (_13499_, _13491_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_13500_, _13499_, _13489_);
  or (_13501_, _13494_, _12797_);
  and (_13502_, _13501_, _13500_);
  and (_13503_, _12802_, _12191_);
  and (_13504_, _13503_, _13488_);
  or (_40664_, _13504_, _13502_);
  or (_13505_, _13491_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_13506_, _13505_, _13489_);
  or (_13507_, _13494_, _13006_);
  and (_13508_, _13507_, _13506_);
  and (_13509_, _13011_, _12191_);
  and (_13510_, _13509_, _13488_);
  or (_40665_, _13510_, _13508_);
  or (_13511_, _13491_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_13512_, _13511_, _13489_);
  and (_13513_, _13200_, _12174_);
  and (_13514_, _13513_, _13197_);
  or (_13515_, _13494_, _13514_);
  and (_13516_, _13515_, _13512_);
  and (_13517_, _13209_, _12191_);
  and (_13518_, _13517_, _13488_);
  or (_40667_, _13518_, _13516_);
  or (_13519_, _13491_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_13520_, _13519_, _13489_);
  or (_13521_, _13494_, _13405_);
  and (_13522_, _13521_, _13520_);
  and (_13523_, _13410_, _12191_);
  and (_13524_, _13523_, _13488_);
  or (_40668_, _13524_, _13522_);
  or (_13525_, _13491_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_13526_, _13525_, _13489_);
  nor (_13527_, _06799_, _12175_);
  or (_13528_, _13494_, _13527_);
  and (_13529_, _13528_, _13526_);
  and (_13530_, _06823_, _12191_);
  and (_13531_, _13488_, _13530_);
  or (_40669_, _13531_, _13529_);
  and (_13532_, _11996_, _04799_);
  not (_13533_, _13532_);
  or (_13534_, _13533_, _12171_);
  and (_13535_, _12187_, _03497_);
  not (_13536_, _13535_);
  or (_13537_, _13532_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_13538_, _13537_, _13536_);
  and (_13539_, _13538_, _13534_);
  and (_13540_, _13535_, _13480_);
  or (_40673_, _13540_, _13539_);
  or (_13541_, _13533_, _12388_);
  or (_13542_, _13532_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_13543_, _13542_, _13536_);
  and (_13544_, _13543_, _13541_);
  and (_13545_, _13535_, _13486_);
  or (_40674_, _13545_, _13544_);
  and (_13546_, _12194_, _03497_);
  not (_13547_, _13546_);
  not (_13548_, _12179_);
  nor (_13549_, _13548_, _04711_);
  and (_13550_, _12178_, _13549_);
  or (_13551_, _13550_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_13552_, _13551_, _13547_);
  not (_13553_, _13550_);
  or (_13554_, _13553_, _12595_);
  and (_13555_, _13554_, _13552_);
  and (_13556_, _13546_, _13497_);
  or (_40675_, _13556_, _13555_);
  or (_13557_, _13550_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_13558_, _13557_, _13547_);
  or (_13559_, _13553_, _12797_);
  and (_13560_, _13559_, _13558_);
  and (_13561_, _13546_, _13503_);
  or (_40676_, _13561_, _13560_);
  or (_13562_, _13550_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_13563_, _13562_, _13547_);
  or (_13564_, _13553_, _13006_);
  and (_13565_, _13564_, _13563_);
  and (_13566_, _13546_, _13509_);
  or (_40678_, _13566_, _13565_);
  or (_13567_, _13550_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_13568_, _13567_, _13547_);
  or (_13569_, _13553_, _13514_);
  and (_13570_, _13569_, _13568_);
  and (_13571_, _13546_, _13517_);
  or (_40679_, _13571_, _13570_);
  or (_13572_, _13550_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_13573_, _13572_, _13547_);
  or (_13574_, _13553_, _13405_);
  and (_13575_, _13574_, _13573_);
  and (_13576_, _13546_, _13523_);
  or (_40680_, _13576_, _13575_);
  or (_13577_, _13550_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_13578_, _13577_, _13547_);
  or (_13579_, _13553_, _13527_);
  and (_13580_, _13579_, _13578_);
  and (_13581_, _13546_, _13530_);
  or (_40681_, _13581_, _13580_);
  and (_13582_, _11995_, _05122_);
  and (_13583_, _13582_, _11994_);
  not (_13584_, _13583_);
  or (_13585_, _13584_, _12171_);
  and (_13586_, _12185_, _05132_);
  and (_13587_, _13586_, _03499_);
  not (_13588_, _13587_);
  or (_13589_, _13583_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_13590_, _13589_, _13588_);
  and (_13591_, _13590_, _13585_);
  and (_13592_, _13587_, _13480_);
  or (_40686_, _13592_, _13591_);
  or (_13593_, _13584_, _12388_);
  or (_13594_, _13583_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_13595_, _13594_, _13588_);
  and (_13596_, _13595_, _13593_);
  and (_13597_, _13587_, _13486_);
  or (_40687_, _13597_, _13596_);
  and (_13598_, _12191_, _05129_);
  and (_13599_, _13598_, _05132_);
  and (_13600_, _13599_, _03499_);
  not (_13601_, _13600_);
  and (_13602_, _12176_, _05122_);
  and (_13603_, _13602_, _12181_);
  or (_13604_, _13603_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_13605_, _13604_, _13601_);
  not (_13606_, _13603_);
  or (_13607_, _13606_, _12595_);
  and (_13608_, _13607_, _13605_);
  and (_13609_, _13600_, _13497_);
  or (_40688_, _13609_, _13608_);
  or (_13610_, _13603_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_13611_, _13610_, _13601_);
  or (_13613_, _13606_, _12797_);
  and (_13614_, _13613_, _13611_);
  and (_13615_, _13600_, _13503_);
  or (_40689_, _13615_, _13614_);
  or (_13616_, _13603_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_13617_, _13616_, _13601_);
  or (_13618_, _13606_, _13006_);
  and (_13619_, _13618_, _13617_);
  and (_13620_, _13600_, _13509_);
  or (_40690_, _13620_, _13619_);
  or (_13622_, _13603_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_13623_, _13622_, _13601_);
  or (_13624_, _13606_, _13514_);
  and (_13625_, _13624_, _13623_);
  and (_13626_, _13600_, _13517_);
  or (_40692_, _13626_, _13625_);
  or (_13627_, _13603_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_13628_, _13627_, _13601_);
  or (_13629_, _13606_, _13405_);
  and (_13630_, _13629_, _13628_);
  and (_13632_, _13600_, _13523_);
  or (_40693_, _13632_, _13630_);
  or (_13633_, _13603_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_13634_, _13633_, _13601_);
  or (_13635_, _13606_, _13527_);
  and (_13636_, _13635_, _13634_);
  and (_13637_, _13600_, _13530_);
  or (_40694_, _13637_, _13636_);
  and (_13638_, _13582_, _13417_);
  not (_13639_, _13638_);
  or (_13641_, _13639_, _12171_);
  and (_13642_, _12180_, _04556_);
  and (_13643_, _13602_, _13642_);
  or (_13644_, _13643_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_13645_, _13586_, _04804_);
  not (_13646_, _13645_);
  and (_13647_, _13646_, _13644_);
  and (_13648_, _13647_, _13641_);
  and (_13649_, _13645_, _13480_);
  or (_40698_, _13649_, _13648_);
  or (_13651_, _13639_, _12388_);
  or (_13652_, _13638_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_13653_, _13652_, _13646_);
  and (_13654_, _13653_, _13651_);
  and (_13655_, _13645_, _13486_);
  or (_40699_, _13655_, _13654_);
  and (_13656_, _13599_, _04804_);
  not (_13657_, _13656_);
  or (_13658_, _13643_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_13659_, _13658_, _13657_);
  not (_13661_, _13643_);
  or (_13662_, _13661_, _12595_);
  and (_13663_, _13662_, _13659_);
  and (_13664_, _13656_, _13497_);
  or (_40700_, _13664_, _13663_);
  or (_13665_, _13643_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_13666_, _13665_, _13657_);
  or (_13667_, _13661_, _12797_);
  and (_13668_, _13667_, _13666_);
  and (_13669_, _13656_, _13503_);
  or (_40701_, _13669_, _13668_);
  or (_13671_, _13643_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_13672_, _13671_, _13657_);
  or (_13673_, _13661_, _13006_);
  and (_13674_, _13673_, _13672_);
  and (_13675_, _13656_, _13509_);
  or (_40702_, _13675_, _13674_);
  or (_13676_, _13643_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_13677_, _13676_, _13657_);
  or (_13678_, _13661_, _13514_);
  and (_13680_, _13678_, _13677_);
  and (_13681_, _13656_, _13517_);
  or (_40704_, _13681_, _13680_);
  or (_13682_, _13643_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_13683_, _13682_, _13657_);
  or (_13684_, _13661_, _13405_);
  and (_13685_, _13684_, _13683_);
  and (_13686_, _13656_, _13523_);
  or (_40705_, _13686_, _13685_);
  and (_13687_, _13643_, _13527_);
  nor (_13689_, _13643_, _05166_);
  or (_13690_, _13689_, _13656_);
  or (_13691_, _13690_, _13687_);
  or (_13692_, _13657_, _13530_);
  and (_40706_, _13692_, _13691_);
  and (_13693_, _13582_, _13471_);
  not (_13694_, _13693_);
  or (_13695_, _13694_, _12171_);
  and (_13696_, _13586_, _05967_);
  not (_13697_, _13696_);
  or (_13699_, _13693_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_13700_, _13699_, _13697_);
  and (_13701_, _13700_, _13695_);
  and (_13702_, _13696_, _13480_);
  or (_40710_, _13702_, _13701_);
  or (_13703_, _13694_, _12388_);
  or (_13704_, _13693_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_13705_, _13704_, _13697_);
  and (_13706_, _13705_, _13703_);
  and (_13707_, _13696_, _13486_);
  or (_40711_, _13707_, _13706_);
  and (_13709_, _13599_, _05967_);
  not (_13710_, _13709_);
  and (_13711_, _13602_, _13490_);
  or (_13712_, _13711_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_13713_, _13712_, _13710_);
  not (_13714_, _13711_);
  or (_13715_, _13714_, _12595_);
  and (_13716_, _13715_, _13713_);
  and (_13717_, _13709_, _13497_);
  or (_40712_, _13717_, _13716_);
  or (_13719_, _13711_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_13720_, _13719_, _13710_);
  or (_13721_, _13714_, _12797_);
  and (_13722_, _13721_, _13720_);
  and (_13723_, _13709_, _13503_);
  or (_40713_, _13723_, _13722_);
  or (_13724_, _13711_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_13725_, _13724_, _13710_);
  or (_13726_, _13714_, _13006_);
  and (_13728_, _13726_, _13725_);
  and (_13729_, _13709_, _13509_);
  or (_40715_, _13729_, _13728_);
  or (_13730_, _13711_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_13731_, _13730_, _13710_);
  or (_13732_, _13714_, _13514_);
  and (_13733_, _13732_, _13731_);
  and (_13734_, _13709_, _13517_);
  or (_40716_, _13734_, _13733_);
  or (_13735_, _13711_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_13737_, _13735_, _13710_);
  or (_13738_, _13714_, _13405_);
  and (_13739_, _13738_, _13737_);
  and (_13740_, _13709_, _13523_);
  or (_40717_, _13740_, _13739_);
  or (_13741_, _13711_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_13742_, _13741_, _13710_);
  or (_13743_, _13714_, _13527_);
  and (_13744_, _13743_, _13742_);
  and (_13745_, _13709_, _13530_);
  or (_40718_, _13745_, _13744_);
  and (_13746_, _13582_, _04799_);
  not (_13747_, _13746_);
  or (_13748_, _13747_, _12171_);
  and (_13749_, _13586_, _03497_);
  not (_13750_, _13749_);
  or (_13751_, _13746_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_13752_, _13751_, _13750_);
  and (_13753_, _13752_, _13748_);
  and (_13754_, _13749_, _13480_);
  or (_40722_, _13754_, _13753_);
  or (_13755_, _13747_, _12388_);
  or (_13756_, _13746_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_13757_, _13756_, _13750_);
  and (_13758_, _13757_, _13755_);
  and (_13759_, _13749_, _13486_);
  or (_40723_, _13759_, _13758_);
  and (_13760_, _13599_, _03497_);
  not (_13761_, _13760_);
  and (_13762_, _13602_, _13549_);
  or (_13763_, _13762_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_13764_, _13763_, _13761_);
  not (_13765_, _13762_);
  or (_13766_, _13765_, _12595_);
  and (_13767_, _13766_, _13764_);
  and (_13768_, _13760_, _13497_);
  or (_40724_, _13768_, _13767_);
  or (_13769_, _13762_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_13770_, _13769_, _13761_);
  or (_13771_, _13765_, _12797_);
  and (_13772_, _13771_, _13770_);
  and (_13773_, _13760_, _13503_);
  or (_40725_, _13773_, _13772_);
  or (_13774_, _13762_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_13775_, _13774_, _13761_);
  or (_13776_, _13765_, _13006_);
  and (_13777_, _13776_, _13775_);
  and (_13778_, _13760_, _13509_);
  or (_40727_, _13778_, _13777_);
  or (_13779_, _13762_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_13780_, _13779_, _13761_);
  or (_13781_, _13765_, _13514_);
  and (_13782_, _13781_, _13780_);
  and (_13783_, _13760_, _13517_);
  or (_40728_, _13783_, _13782_);
  or (_13784_, _13762_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_13785_, _13784_, _13761_);
  or (_13786_, _13765_, _13405_);
  and (_13787_, _13786_, _13785_);
  and (_13788_, _13760_, _13523_);
  or (_40729_, _13788_, _13787_);
  or (_13789_, _13762_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_13790_, _13789_, _13761_);
  or (_13791_, _13765_, _13527_);
  and (_13792_, _13791_, _13790_);
  and (_13793_, _13760_, _13530_);
  or (_40730_, _13793_, _13792_);
  and (_13794_, _05123_, _04951_);
  and (_13795_, _13794_, _11994_);
  not (_13796_, _13795_);
  or (_13797_, _13796_, _12171_);
  and (_13798_, _05138_, _12192_);
  and (_13799_, _13798_, _03499_);
  not (_13800_, _13799_);
  or (_13801_, _13795_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_13802_, _13801_, _13800_);
  and (_13803_, _13802_, _13797_);
  and (_13804_, _13799_, _13480_);
  or (_40735_, _13804_, _13803_);
  or (_13805_, _13796_, _12388_);
  or (_13806_, _13795_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_13807_, _13806_, _13800_);
  and (_13808_, _13807_, _13805_);
  and (_13809_, _13799_, _13486_);
  or (_40736_, _13809_, _13808_);
  or (_13810_, _13795_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_13811_, _13810_, _13800_);
  or (_13812_, _13796_, _13436_);
  and (_13813_, _13812_, _13811_);
  and (_13814_, _12600_, _05137_);
  and (_13815_, _13799_, _13814_);
  or (_40737_, _13815_, _13813_);
  or (_13816_, _13795_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_13817_, _13816_, _13800_);
  or (_13818_, _13796_, _13443_);
  and (_13819_, _13818_, _13817_);
  and (_13820_, _12802_, _05137_);
  and (_13821_, _13799_, _13820_);
  or (_40738_, _13821_, _13819_);
  or (_13822_, _13795_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_13823_, _13822_, _13800_);
  or (_13824_, _13796_, _13450_);
  and (_13825_, _13824_, _13823_);
  and (_13826_, _13011_, _05137_);
  and (_13827_, _13799_, _13826_);
  or (_40739_, _13827_, _13825_);
  or (_13828_, _13795_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_13829_, _13828_, _13800_);
  or (_13830_, _13796_, _13202_);
  and (_13831_, _13830_, _13829_);
  and (_13832_, _13209_, _05137_);
  and (_13833_, _13799_, _13832_);
  or (_40741_, _13833_, _13831_);
  or (_13834_, _13795_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_13835_, _13834_, _13800_);
  or (_13836_, _13796_, _13462_);
  and (_13837_, _13836_, _13835_);
  and (_13838_, _13410_, _05137_);
  and (_13839_, _13799_, _13838_);
  or (_40742_, _13839_, _13837_);
  nor (_13840_, _13795_, \oc8051_golden_model_1.IRAM[8] [7]);
  nor (_13841_, _13796_, _06800_);
  or (_13842_, _13841_, _13840_);
  nor (_13843_, _13842_, _13799_);
  and (_13844_, _13799_, _06824_);
  or (_40743_, _13844_, _13843_);
  and (_13845_, _13794_, _13417_);
  not (_13846_, _13845_);
  or (_13847_, _13846_, _12171_);
  or (_13848_, _13845_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_13849_, _13798_, _04804_);
  not (_13850_, _13849_);
  and (_13851_, _13850_, _13848_);
  and (_13852_, _13851_, _13847_);
  and (_13853_, _13849_, _13480_);
  or (_40747_, _13853_, _13852_);
  or (_13854_, _13846_, _12388_);
  or (_13855_, _13845_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_13856_, _13855_, _13850_);
  and (_13857_, _13856_, _13854_);
  and (_13858_, _13849_, _13486_);
  or (_40748_, _13858_, _13857_);
  or (_13859_, _13845_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_13860_, _13859_, _13850_);
  or (_13861_, _13846_, _13436_);
  and (_13862_, _13861_, _13860_);
  and (_13863_, _13849_, _13814_);
  or (_40749_, _13863_, _13862_);
  or (_13864_, _13845_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_13865_, _13864_, _13850_);
  or (_13866_, _13846_, _13443_);
  and (_13867_, _13866_, _13865_);
  and (_13868_, _13849_, _13820_);
  or (_40750_, _13868_, _13867_);
  or (_13869_, _13846_, _13450_);
  or (_13870_, _13845_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_13871_, _13870_, _13850_);
  and (_13872_, _13871_, _13869_);
  and (_13873_, _13849_, _13826_);
  or (_40751_, _13873_, _13872_);
  or (_13874_, _13845_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_13875_, _13874_, _13850_);
  or (_13876_, _13846_, _13202_);
  and (_13877_, _13876_, _13875_);
  and (_13878_, _13849_, _13832_);
  or (_40753_, _13878_, _13877_);
  or (_13879_, _13845_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_13880_, _13879_, _13850_);
  or (_13881_, _13846_, _13462_);
  and (_13882_, _13881_, _13880_);
  and (_13883_, _13849_, _13838_);
  or (_40754_, _13883_, _13882_);
  or (_13884_, _13845_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_13885_, _13884_, _13850_);
  or (_13886_, _13846_, _06800_);
  and (_13887_, _13886_, _13885_);
  and (_13888_, _13849_, _06824_);
  or (_40755_, _13888_, _13887_);
  and (_13889_, _13794_, _13471_);
  not (_13890_, _13889_);
  or (_13891_, _13890_, _12171_);
  or (_13892_, _13889_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_13893_, _13798_, _05967_);
  not (_13894_, _13893_);
  and (_13895_, _13894_, _13892_);
  and (_13896_, _13895_, _13891_);
  and (_13897_, _13893_, _13480_);
  or (_40759_, _13897_, _13896_);
  or (_13898_, _13889_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_13899_, _13898_, _13894_);
  or (_13900_, _13890_, _12388_);
  and (_13901_, _13900_, _13899_);
  and (_13902_, _13893_, _13486_);
  or (_40760_, _13902_, _13901_);
  or (_13903_, _13889_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_13904_, _13903_, _13894_);
  or (_13905_, _13890_, _13436_);
  and (_13906_, _13905_, _13904_);
  and (_13907_, _13893_, _13814_);
  or (_40761_, _13907_, _13906_);
  or (_13908_, _13889_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_13909_, _13908_, _13894_);
  or (_13910_, _13890_, _13443_);
  and (_13911_, _13910_, _13909_);
  and (_13912_, _13893_, _13820_);
  or (_40762_, _13912_, _13911_);
  or (_13913_, _13889_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_13914_, _13913_, _13894_);
  or (_13915_, _13890_, _13450_);
  and (_13916_, _13915_, _13914_);
  and (_13917_, _13893_, _13826_);
  or (_40764_, _13917_, _13916_);
  or (_13918_, _13889_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_13919_, _13918_, _13894_);
  or (_13920_, _13890_, _13202_);
  and (_13921_, _13920_, _13919_);
  and (_13922_, _13893_, _13832_);
  or (_40765_, _13922_, _13921_);
  or (_13923_, _13889_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_13924_, _13923_, _13894_);
  or (_13925_, _13890_, _13462_);
  and (_13926_, _13925_, _13924_);
  and (_13927_, _13893_, _13838_);
  or (_40766_, _13927_, _13926_);
  or (_13928_, _13889_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_13929_, _13928_, _13894_);
  or (_13930_, _13890_, _06800_);
  and (_13931_, _13930_, _13929_);
  and (_13932_, _13893_, _06824_);
  or (_40767_, _13932_, _13931_);
  and (_13933_, _13794_, _04799_);
  not (_13934_, _13933_);
  or (_13935_, _13934_, _12171_);
  and (_13936_, _13798_, _03497_);
  not (_13937_, _13936_);
  or (_13938_, _13933_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_13939_, _13938_, _13937_);
  and (_13940_, _13939_, _13935_);
  and (_13941_, _13936_, _13480_);
  or (_40771_, _13941_, _13940_);
  or (_13942_, _13934_, _12388_);
  or (_13943_, _13933_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_13944_, _13943_, _13937_);
  and (_13945_, _13944_, _13942_);
  and (_13946_, _13936_, _13486_);
  or (_40772_, _13946_, _13945_);
  or (_13947_, _13933_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_13948_, _13947_, _13937_);
  or (_13949_, _13934_, _13436_);
  and (_13950_, _13949_, _13948_);
  and (_13951_, _13936_, _13814_);
  or (_40773_, _13951_, _13950_);
  or (_13952_, _13934_, _13443_);
  or (_13953_, _13933_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_13954_, _13953_, _13937_);
  and (_13955_, _13954_, _13952_);
  and (_13956_, _13936_, _13820_);
  or (_40774_, _13956_, _13955_);
  or (_13957_, _13934_, _13450_);
  or (_13958_, _13933_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_13959_, _13958_, _13937_);
  and (_13960_, _13959_, _13957_);
  and (_13961_, _13936_, _13826_);
  or (_40776_, _13961_, _13960_);
  or (_13962_, _13934_, _13202_);
  or (_13963_, _13933_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_13964_, _13963_, _13937_);
  and (_13965_, _13964_, _13962_);
  and (_13966_, _13936_, _13832_);
  or (_40777_, _13966_, _13965_);
  or (_13967_, _13934_, _13462_);
  or (_13968_, _13933_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_13969_, _13968_, _13937_);
  and (_13970_, _13969_, _13967_);
  and (_13971_, _13936_, _13838_);
  or (_40778_, _13971_, _13970_);
  or (_13972_, _13934_, _06800_);
  or (_13973_, _13933_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_13974_, _13973_, _13937_);
  and (_13975_, _13974_, _13972_);
  and (_13976_, _13936_, _06824_);
  or (_40779_, _13976_, _13975_);
  and (_13977_, _11994_, _05124_);
  not (_13978_, _13977_);
  or (_13979_, _13978_, _12171_);
  and (_13980_, _05139_, _03499_);
  not (_13981_, _13980_);
  or (_13982_, _13977_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_13983_, _13982_, _13981_);
  and (_13984_, _13983_, _13979_);
  and (_13985_, _13980_, _13480_);
  or (_40783_, _13985_, _13984_);
  or (_13986_, _13977_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_13987_, _13986_, _13981_);
  or (_13988_, _13978_, _12388_);
  and (_13989_, _13988_, _13987_);
  and (_13990_, _13980_, _13486_);
  or (_40784_, _13990_, _13989_);
  or (_13991_, _13977_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_13992_, _13991_, _13981_);
  or (_13993_, _13978_, _13436_);
  and (_13994_, _13993_, _13992_);
  and (_13995_, _13980_, _13814_);
  or (_40786_, _13995_, _13994_);
  or (_13996_, _13977_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_13997_, _13996_, _13981_);
  or (_13998_, _13978_, _13443_);
  and (_13999_, _13998_, _13997_);
  and (_14000_, _13980_, _13820_);
  or (_40787_, _14000_, _13999_);
  or (_14001_, _13977_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_14002_, _14001_, _13981_);
  or (_14003_, _13978_, _13450_);
  and (_14004_, _14003_, _14002_);
  and (_14005_, _13980_, _13826_);
  or (_40788_, _14005_, _14004_);
  or (_14006_, _13977_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_14007_, _14006_, _13981_);
  or (_14008_, _13978_, _13202_);
  and (_14009_, _14008_, _14007_);
  and (_14010_, _13980_, _13832_);
  or (_40789_, _14010_, _14009_);
  or (_14011_, _13977_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_14012_, _14011_, _13981_);
  or (_14013_, _13978_, _13462_);
  and (_14014_, _14013_, _14012_);
  and (_14015_, _13980_, _13838_);
  or (_40790_, _14015_, _14014_);
  or (_14016_, _13977_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_14017_, _14016_, _13981_);
  or (_14018_, _13978_, _06800_);
  and (_14019_, _14018_, _14017_);
  and (_14020_, _13980_, _06824_);
  or (_40792_, _14020_, _14019_);
  and (_14021_, _13417_, _05124_);
  not (_14022_, _14021_);
  or (_14023_, _14022_, _12171_);
  or (_14024_, _14021_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_14025_, _05139_, _04804_);
  not (_14026_, _14025_);
  and (_14027_, _14026_, _14024_);
  and (_14028_, _14027_, _14023_);
  and (_14029_, _14025_, _13480_);
  or (_40795_, _14029_, _14028_);
  or (_14030_, _14021_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_14031_, _14030_, _14026_);
  or (_14032_, _14022_, _12388_);
  and (_14033_, _14032_, _14031_);
  and (_14034_, _14025_, _13486_);
  or (_40796_, _14034_, _14033_);
  or (_14035_, _14021_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_14036_, _14035_, _14026_);
  or (_14037_, _14022_, _13436_);
  and (_14038_, _14037_, _14036_);
  and (_14039_, _14025_, _13814_);
  or (_40798_, _14039_, _14038_);
  or (_14040_, _14021_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_14041_, _14040_, _14026_);
  or (_14042_, _14022_, _13443_);
  and (_14043_, _14042_, _14041_);
  and (_14044_, _14025_, _13820_);
  or (_40799_, _14044_, _14043_);
  or (_14045_, _14021_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_14046_, _14045_, _14026_);
  or (_14047_, _14022_, _13450_);
  and (_14048_, _14047_, _14046_);
  and (_14049_, _14025_, _13826_);
  or (_40800_, _14049_, _14048_);
  or (_14050_, _14021_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_14051_, _14050_, _14026_);
  or (_14052_, _14022_, _13202_);
  and (_14053_, _14052_, _14051_);
  and (_14054_, _14025_, _13832_);
  or (_40801_, _14054_, _14053_);
  or (_14055_, _14021_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_14056_, _14055_, _14026_);
  or (_14057_, _14022_, _13462_);
  and (_14058_, _14057_, _14056_);
  and (_14059_, _14025_, _13838_);
  or (_40802_, _14059_, _14058_);
  nor (_14060_, _14021_, \oc8051_golden_model_1.IRAM[13] [7]);
  nor (_14061_, _14022_, _06800_);
  or (_14062_, _14061_, _14060_);
  nand (_14063_, _14062_, _14026_);
  or (_14064_, _14026_, _06824_);
  and (_40804_, _14064_, _14063_);
  and (_14065_, _13471_, _05124_);
  not (_14066_, _14065_);
  or (_14067_, _14066_, _12171_);
  or (_14068_, _14065_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_14069_, _05967_, _05139_);
  not (_14070_, _14069_);
  and (_14071_, _14070_, _14068_);
  and (_14072_, _14071_, _14067_);
  and (_14073_, _14069_, _13480_);
  or (_40807_, _14073_, _14072_);
  or (_14074_, _14066_, _12388_);
  or (_14075_, _14065_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_14076_, _14075_, _14070_);
  and (_14077_, _14076_, _14074_);
  and (_14078_, _14069_, _13486_);
  or (_40809_, _14078_, _14077_);
  or (_14079_, _14065_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_14080_, _14079_, _14070_);
  or (_14081_, _14066_, _13436_);
  and (_14082_, _14081_, _14080_);
  and (_14083_, _14069_, _13814_);
  or (_40810_, _14083_, _14082_);
  or (_14084_, _14065_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_14085_, _14084_, _14070_);
  or (_14086_, _14066_, _13443_);
  and (_14087_, _14086_, _14085_);
  and (_14088_, _14069_, _13820_);
  or (_40811_, _14088_, _14087_);
  or (_14089_, _14065_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_14090_, _14089_, _14070_);
  or (_14091_, _14066_, _13450_);
  and (_14092_, _14091_, _14090_);
  and (_14093_, _14069_, _13826_);
  or (_40812_, _14093_, _14092_);
  or (_14094_, _14065_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_14095_, _14094_, _14070_);
  or (_14096_, _14066_, _13202_);
  and (_14097_, _14096_, _14095_);
  and (_14098_, _14069_, _13832_);
  or (_40813_, _14098_, _14097_);
  or (_14099_, _14065_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_14100_, _14099_, _14070_);
  or (_14101_, _14066_, _13462_);
  and (_14102_, _14101_, _14100_);
  and (_14103_, _14069_, _13838_);
  or (_40815_, _14103_, _14102_);
  or (_14104_, _14065_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_14105_, _14104_, _14070_);
  or (_14106_, _14066_, _06800_);
  and (_14107_, _14106_, _14105_);
  and (_14108_, _14069_, _06824_);
  or (_40816_, _14108_, _14107_);
  or (_14109_, _12171_, _05143_);
  or (_14110_, _05125_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_14111_, _14110_, _05141_);
  and (_14112_, _14111_, _14109_);
  and (_14113_, _13480_, _05140_);
  or (_40819_, _14113_, _14112_);
  or (_14114_, _05125_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_14115_, _14114_, _05141_);
  or (_14116_, _12388_, _05143_);
  and (_14117_, _14116_, _14115_);
  and (_14118_, _13486_, _05140_);
  or (_40821_, _14118_, _14117_);
  or (_14119_, _05125_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_14120_, _14119_, _05141_);
  or (_14121_, _13436_, _05143_);
  and (_14122_, _14121_, _14120_);
  and (_14123_, _13814_, _05140_);
  or (_40822_, _14123_, _14122_);
  or (_14124_, _05125_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_14125_, _14124_, _05141_);
  or (_14126_, _13443_, _05143_);
  and (_14127_, _14126_, _14125_);
  and (_14128_, _13820_, _05140_);
  or (_40823_, _14128_, _14127_);
  or (_14129_, _05125_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_14130_, _14129_, _05141_);
  or (_14131_, _13450_, _05143_);
  and (_14132_, _14131_, _14130_);
  and (_14133_, _13826_, _05140_);
  or (_40824_, _14133_, _14132_);
  or (_14134_, _05125_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_14135_, _14134_, _05141_);
  or (_14136_, _13202_, _05143_);
  and (_14137_, _14136_, _14135_);
  and (_14138_, _13832_, _05140_);
  or (_40825_, _14138_, _14137_);
  or (_14139_, _05125_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_14140_, _14139_, _05141_);
  or (_14141_, _13462_, _05143_);
  and (_14142_, _14141_, _14140_);
  and (_14143_, _13838_, _05140_);
  or (_40827_, _14143_, _14142_);
  nor (_14144_, _43000_, _07418_);
  nor (_14145_, _05248_, _07418_);
  and (_14146_, _12128_, _05248_);
  or (_14147_, _14146_, _14145_);
  and (_14148_, _14147_, _03780_);
  nor (_14149_, _05666_, _06830_);
  or (_14150_, _14149_, _14145_);
  or (_14151_, _14150_, _04081_);
  and (_14152_, _05248_, \oc8051_golden_model_1.ACC [0]);
  or (_14153_, _14152_, _14145_);
  and (_14154_, _14153_, _04409_);
  nor (_14155_, _04409_, _07418_);
  or (_14156_, _14155_, _03610_);
  or (_14157_, _14156_, _14154_);
  and (_14158_, _14157_, _04055_);
  and (_14159_, _14158_, _14151_);
  and (_14160_, _12021_, _05910_);
  nor (_14161_, _05910_, _07418_);
  or (_14162_, _14161_, _14160_);
  and (_14163_, _14162_, _03715_);
  or (_14164_, _14163_, _14159_);
  and (_14165_, _14164_, _03996_);
  and (_14166_, _05248_, _04620_);
  or (_14167_, _14166_, _14145_);
  and (_14168_, _14167_, _03723_);
  or (_14169_, _14168_, _03729_);
  or (_14170_, _14169_, _14165_);
  or (_14171_, _14153_, _03737_);
  and (_14172_, _14171_, _03736_);
  and (_14173_, _14172_, _14170_);
  and (_14174_, _14145_, _03714_);
  or (_14175_, _14174_, _03719_);
  or (_14176_, _14175_, _14173_);
  or (_14177_, _14150_, _06840_);
  and (_14178_, _14177_, _14176_);
  or (_14179_, _14178_, _06869_);
  nor (_14180_, _07351_, _07349_);
  nor (_14181_, _14180_, _07352_);
  or (_14182_, _14181_, _06875_);
  and (_14183_, _14182_, _03710_);
  and (_14184_, _14183_, _14179_);
  nor (_14185_, _12052_, _07391_);
  or (_14186_, _14185_, _14161_);
  and (_14187_, _14186_, _03505_);
  or (_14188_, _14187_, _07390_);
  or (_14189_, _14188_, _14184_);
  or (_14190_, _14167_, _06838_);
  and (_14191_, _14190_, _07400_);
  and (_14192_, _14191_, _14189_);
  and (_14193_, _06546_, _05248_);
  or (_14194_, _14193_, _14145_);
  and (_14195_, _14194_, _04481_);
  or (_14196_, _14195_, _03222_);
  or (_14197_, _14196_, _14192_);
  nor (_14198_, _12109_, _06830_);
  or (_14199_, _14145_, _03589_);
  or (_14200_, _14199_, _14198_);
  and (_14201_, _14200_, _07411_);
  and (_14202_, _14201_, _14197_);
  nor (_14203_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_14204_, _14203_, _07330_);
  or (_14205_, _07760_, _14204_);
  nand (_14206_, _07760_, _03335_);
  and (_14207_, _14206_, _07405_);
  and (_14208_, _14207_, _14205_);
  or (_14209_, _14208_, _08828_);
  or (_14210_, _14209_, _14202_);
  and (_14211_, _12124_, _05248_);
  or (_14212_, _14145_, _07766_);
  or (_14213_, _14212_, _14211_);
  and (_14214_, _05248_, _06274_);
  or (_14215_, _14214_, _14145_);
  or (_14216_, _14215_, _05886_);
  and (_14217_, _14216_, _07778_);
  and (_14218_, _14217_, _14213_);
  and (_14219_, _14218_, _14210_);
  or (_14220_, _14219_, _14148_);
  and (_14221_, _14220_, _07777_);
  nand (_14222_, _14215_, _03622_);
  nor (_14223_, _14222_, _14149_);
  or (_14224_, _14223_, _14221_);
  and (_14225_, _14224_, _06828_);
  or (_14226_, _14145_, _05666_);
  and (_14227_, _14153_, _03790_);
  and (_14228_, _14227_, _14226_);
  or (_14229_, _14228_, _03624_);
  or (_14230_, _14229_, _14225_);
  nor (_14231_, _12122_, _06830_);
  or (_14232_, _14145_, _07795_);
  or (_14233_, _14232_, _14231_);
  and (_14234_, _14233_, _07793_);
  and (_14235_, _14234_, _14230_);
  nor (_14236_, _12003_, _06830_);
  or (_14237_, _14236_, _14145_);
  and (_14238_, _14237_, _03785_);
  or (_14239_, _14238_, _03815_);
  or (_14240_, _14239_, _14235_);
  or (_14241_, _14150_, _04246_);
  and (_14242_, _14241_, _03823_);
  and (_14243_, _14242_, _14240_);
  and (_14244_, _14145_, _03453_);
  or (_14245_, _14244_, _03447_);
  or (_14246_, _14245_, _14243_);
  or (_14247_, _14150_, _03514_);
  and (_14248_, _14247_, _43000_);
  and (_14249_, _14248_, _14246_);
  or (_14250_, _14249_, _14144_);
  and (_43480_, _14250_, _41806_);
  nor (_14251_, _43000_, _07412_);
  or (_14252_, _05248_, \oc8051_golden_model_1.B [1]);
  and (_14253_, _12213_, _05248_);
  not (_14254_, _14253_);
  and (_14255_, _14254_, _14252_);
  or (_14256_, _14255_, _04081_);
  nand (_14257_, _05248_, _03274_);
  and (_14258_, _14257_, _14252_);
  and (_14259_, _14258_, _04409_);
  nor (_14260_, _04409_, _07412_);
  or (_14261_, _14260_, _03610_);
  or (_14262_, _14261_, _14259_);
  and (_14263_, _14262_, _04055_);
  and (_14264_, _14263_, _14256_);
  not (_14265_, _03730_);
  and (_14266_, _12224_, _05910_);
  nor (_14267_, _05910_, _07412_);
  or (_14268_, _14267_, _03723_);
  or (_14269_, _14268_, _14266_);
  and (_14270_, _14269_, _14265_);
  or (_14271_, _14270_, _14264_);
  nor (_14272_, _05248_, _07412_);
  and (_14273_, _05248_, _06764_);
  or (_14274_, _14273_, _14272_);
  or (_14275_, _14274_, _03996_);
  and (_14276_, _14275_, _14271_);
  or (_14277_, _14276_, _03729_);
  or (_14278_, _14258_, _03737_);
  and (_14279_, _14278_, _03736_);
  and (_14280_, _14279_, _14277_);
  and (_14281_, _12211_, _05910_);
  or (_14282_, _14281_, _14267_);
  and (_14283_, _14282_, _03714_);
  or (_14284_, _14283_, _14280_);
  and (_14285_, _14284_, _06840_);
  and (_14286_, _14266_, _12239_);
  or (_14287_, _14286_, _14267_);
  and (_14288_, _14287_, _03719_);
  or (_14289_, _14288_, _06869_);
  or (_14290_, _14289_, _14285_);
  or (_14291_, _07296_, _07295_);
  nand (_14292_, _14291_, _07353_);
  or (_14293_, _14291_, _07353_);
  and (_14294_, _14293_, _14292_);
  or (_14295_, _14294_, _06875_);
  and (_14296_, _14295_, _03710_);
  and (_14297_, _14296_, _14290_);
  nor (_14298_, _12256_, _07391_);
  or (_14299_, _14298_, _14267_);
  and (_14300_, _14299_, _03505_);
  or (_14301_, _14300_, _07390_);
  or (_14302_, _14301_, _14297_);
  or (_14303_, _14274_, _06838_);
  and (_14304_, _14303_, _14302_);
  or (_14305_, _14304_, _04481_);
  and (_14306_, _06501_, _05248_);
  or (_14307_, _14272_, _07400_);
  or (_14308_, _14307_, _14306_);
  and (_14309_, _14308_, _03589_);
  and (_14310_, _14309_, _14305_);
  nand (_14311_, _12313_, _05248_);
  and (_14312_, _14252_, _03222_);
  and (_14313_, _14312_, _14311_);
  or (_14314_, _14313_, _07405_);
  or (_14315_, _14314_, _14310_);
  and (_14316_, _07760_, _07707_);
  nor (_14317_, _07755_, _07754_);
  or (_14318_, _14317_, _07756_);
  nor (_14319_, _14318_, _07760_);
  or (_14320_, _14319_, _14316_);
  or (_14321_, _14320_, _07411_);
  and (_14322_, _14321_, _05886_);
  and (_14323_, _14322_, _14315_);
  nand (_14324_, _05248_, _04303_);
  and (_14325_, _14324_, _03601_);
  and (_14326_, _14325_, _14252_);
  or (_14327_, _14326_, _14323_);
  and (_14328_, _14327_, _07766_);
  or (_14329_, _12327_, _06830_);
  and (_14330_, _14252_, _03600_);
  and (_14331_, _14330_, _14329_);
  or (_14332_, _14331_, _14328_);
  and (_14333_, _14332_, _07778_);
  or (_14334_, _12333_, _06830_);
  and (_14335_, _14252_, _03780_);
  and (_14336_, _14335_, _14334_);
  or (_14337_, _14336_, _14333_);
  and (_14338_, _14337_, _07777_);
  or (_14339_, _12207_, _06830_);
  and (_14340_, _14252_, _03622_);
  and (_14341_, _14340_, _14339_);
  or (_14342_, _14341_, _14338_);
  and (_14343_, _14342_, _06828_);
  or (_14344_, _14272_, _05618_);
  and (_14345_, _14258_, _03790_);
  and (_14346_, _14345_, _14344_);
  or (_14347_, _14346_, _14343_);
  and (_14348_, _14347_, _03786_);
  or (_14349_, _14324_, _05618_);
  and (_14350_, _14252_, _03624_);
  and (_14351_, _14350_, _14349_);
  or (_14352_, _14257_, _05618_);
  and (_14353_, _14252_, _03785_);
  and (_14354_, _14353_, _14352_);
  or (_14355_, _14354_, _03815_);
  or (_14356_, _14355_, _14351_);
  or (_14357_, _14356_, _14348_);
  or (_14358_, _14255_, _04246_);
  and (_14359_, _14358_, _03823_);
  and (_14360_, _14359_, _14357_);
  and (_14361_, _14282_, _03453_);
  or (_14362_, _14361_, _03447_);
  or (_14363_, _14362_, _14360_);
  or (_14364_, _14272_, _03514_);
  or (_14365_, _14364_, _14253_);
  and (_14366_, _14365_, _43000_);
  and (_14367_, _14366_, _14363_);
  or (_14368_, _14367_, _14251_);
  and (_43481_, _14368_, _41806_);
  nor (_14369_, _43000_, _07426_);
  nor (_14370_, _05248_, _07426_);
  nor (_14371_, _06830_, _04875_);
  or (_14372_, _14371_, _14370_);
  or (_14373_, _14372_, _06838_);
  and (_14374_, _12411_, _05910_);
  and (_14375_, _14374_, _12443_);
  nor (_14376_, _05910_, _07426_);
  or (_14377_, _14376_, _06840_);
  or (_14378_, _14377_, _14375_);
  or (_14379_, _14372_, _03996_);
  nor (_14380_, _12416_, _06830_);
  or (_14381_, _14380_, _14370_);
  or (_14382_, _14381_, _04081_);
  and (_14383_, _05248_, \oc8051_golden_model_1.ACC [2]);
  or (_14384_, _14383_, _14370_);
  and (_14385_, _14384_, _04409_);
  nor (_14386_, _04409_, _07426_);
  or (_14387_, _14386_, _03610_);
  or (_14388_, _14387_, _14385_);
  and (_14389_, _14388_, _04055_);
  and (_14390_, _14389_, _14382_);
  or (_14391_, _14376_, _14374_);
  and (_14392_, _14391_, _03715_);
  or (_14393_, _14392_, _03723_);
  or (_14394_, _14393_, _14390_);
  and (_14395_, _14394_, _14379_);
  or (_14396_, _14395_, _03729_);
  or (_14397_, _14384_, _03737_);
  and (_14398_, _14397_, _03736_);
  and (_14399_, _14398_, _14396_);
  and (_14400_, _12409_, _05910_);
  or (_14401_, _14400_, _14376_);
  and (_14402_, _14401_, _03714_);
  or (_14403_, _14402_, _03719_);
  or (_14404_, _14403_, _14399_);
  and (_14405_, _14404_, _14378_);
  or (_14406_, _14405_, _06869_);
  nor (_14407_, _07355_, _07252_);
  nor (_14408_, _14407_, _07356_);
  or (_14409_, _14408_, _06875_);
  and (_14410_, _14409_, _03710_);
  and (_14411_, _14410_, _14406_);
  nor (_14412_, _12461_, _07391_);
  or (_14413_, _14412_, _14376_);
  and (_14414_, _14413_, _03505_);
  or (_14415_, _14414_, _07390_);
  or (_14416_, _14415_, _14411_);
  and (_14417_, _14416_, _14373_);
  or (_14418_, _14417_, _04481_);
  and (_14419_, _06637_, _05248_);
  or (_14420_, _14370_, _07400_);
  or (_14421_, _14420_, _14419_);
  and (_14422_, _14421_, _14418_);
  or (_14423_, _14422_, _03222_);
  nor (_14424_, _12519_, _06830_);
  or (_14425_, _14370_, _03589_);
  or (_14426_, _14425_, _14424_);
  and (_14427_, _14426_, _07411_);
  and (_14428_, _14427_, _14423_);
  not (_14429_, _07760_);
  or (_14430_, _14429_, _07697_);
  nor (_14431_, _07756_, _07708_);
  not (_14432_, _14431_);
  and (_14433_, _14432_, _07700_);
  nor (_14434_, _14432_, _07700_);
  nor (_14435_, _14434_, _14433_);
  or (_14436_, _14435_, _07760_);
  and (_14437_, _14436_, _07405_);
  and (_14438_, _14437_, _14430_);
  or (_14439_, _14438_, _08828_);
  or (_14440_, _14439_, _14428_);
  and (_14441_, _12533_, _05248_);
  or (_14442_, _14370_, _07766_);
  or (_14443_, _14442_, _14441_);
  and (_14444_, _05248_, _06332_);
  or (_14445_, _14444_, _14370_);
  or (_14446_, _14445_, _05886_);
  and (_14447_, _14446_, _07778_);
  and (_14448_, _14447_, _14443_);
  and (_14449_, _14448_, _14440_);
  and (_14450_, _12539_, _05248_);
  or (_14451_, _14450_, _14370_);
  and (_14452_, _14451_, _03780_);
  or (_14453_, _14452_, _14449_);
  and (_14454_, _14453_, _07777_);
  or (_14455_, _14370_, _05718_);
  and (_14456_, _14445_, _03622_);
  and (_14457_, _14456_, _14455_);
  or (_14458_, _14457_, _14454_);
  and (_14459_, _14458_, _06828_);
  and (_14460_, _14384_, _03790_);
  and (_14461_, _14460_, _14455_);
  or (_14462_, _14461_, _03624_);
  or (_14463_, _14462_, _14459_);
  nor (_14464_, _12532_, _06830_);
  or (_14465_, _14370_, _07795_);
  or (_14466_, _14465_, _14464_);
  and (_14467_, _14466_, _07793_);
  and (_14468_, _14467_, _14463_);
  nor (_14469_, _12538_, _06830_);
  or (_14470_, _14469_, _14370_);
  and (_14471_, _14470_, _03785_);
  or (_14472_, _14471_, _03815_);
  or (_14473_, _14472_, _14468_);
  or (_14474_, _14381_, _04246_);
  and (_14475_, _14474_, _03823_);
  and (_14476_, _14475_, _14473_);
  and (_14477_, _14401_, _03453_);
  or (_14478_, _14477_, _03447_);
  or (_14479_, _14478_, _14476_);
  and (_14480_, _12592_, _05248_);
  or (_14481_, _14370_, _03514_);
  or (_14482_, _14481_, _14480_);
  and (_14483_, _14482_, _43000_);
  and (_14484_, _14483_, _14479_);
  or (_14485_, _14484_, _14369_);
  and (_43482_, _14485_, _41806_);
  nor (_14486_, _43000_, _07427_);
  nor (_14487_, _05248_, _07427_);
  nor (_14488_, _12718_, _06830_);
  or (_14489_, _14488_, _14487_);
  and (_14490_, _14489_, _03222_);
  nor (_14491_, _05910_, _07427_);
  and (_14492_, _12631_, _05910_);
  or (_14493_, _14492_, _14491_);
  or (_14494_, _14491_, _12648_);
  and (_14495_, _14494_, _14493_);
  or (_14496_, _14495_, _06840_);
  nor (_14497_, _12627_, _06830_);
  or (_14498_, _14497_, _14487_);
  or (_14499_, _14498_, _04081_);
  and (_14500_, _05248_, \oc8051_golden_model_1.ACC [3]);
  or (_14501_, _14500_, _14487_);
  and (_14502_, _14501_, _04409_);
  nor (_14503_, _04409_, _07427_);
  or (_14504_, _14503_, _03610_);
  or (_14505_, _14504_, _14502_);
  and (_14506_, _14505_, _04055_);
  and (_14507_, _14506_, _14499_);
  and (_14508_, _14493_, _03715_);
  or (_14509_, _14508_, _03723_);
  or (_14510_, _14509_, _14507_);
  nor (_14511_, _06830_, _05005_);
  or (_14512_, _14511_, _14487_);
  or (_14513_, _14512_, _03996_);
  and (_14514_, _14513_, _14510_);
  or (_14515_, _14514_, _03729_);
  or (_14516_, _14501_, _03737_);
  and (_14517_, _14516_, _03736_);
  and (_14518_, _14517_, _14515_);
  and (_14519_, _12641_, _05910_);
  or (_14520_, _14519_, _14491_);
  and (_14521_, _14520_, _03714_);
  or (_14522_, _14521_, _03719_);
  or (_14523_, _14522_, _14518_);
  and (_14524_, _14523_, _14496_);
  or (_14525_, _14524_, _06869_);
  nor (_14526_, _07358_, _07194_);
  nor (_14527_, _14526_, _07359_);
  or (_14528_, _14527_, _06875_);
  and (_14529_, _14528_, _03710_);
  and (_14530_, _14529_, _14525_);
  nor (_14531_, _12612_, _07391_);
  or (_14532_, _14531_, _14491_);
  and (_14533_, _14532_, _03505_);
  or (_14534_, _14533_, _07390_);
  or (_14535_, _14534_, _14530_);
  or (_14536_, _14512_, _06838_);
  and (_14537_, _14536_, _14535_);
  or (_14538_, _14537_, _04481_);
  and (_14539_, _06592_, _05248_);
  or (_14540_, _14487_, _07400_);
  or (_14541_, _14540_, _14539_);
  and (_14542_, _14541_, _03589_);
  and (_14543_, _14542_, _14538_);
  or (_14544_, _14543_, _14490_);
  and (_14545_, _14544_, _07411_);
  nand (_14546_, _07760_, _07689_);
  nor (_14547_, _14433_, _07699_);
  nor (_14548_, _14547_, _07692_);
  and (_14549_, _14547_, _07692_);
  or (_14550_, _14549_, _14548_);
  or (_14551_, _14550_, _07760_);
  and (_14552_, _14551_, _07405_);
  and (_14553_, _14552_, _14546_);
  or (_14554_, _14553_, _08828_);
  or (_14555_, _14554_, _14545_);
  and (_14556_, _12733_, _05248_);
  or (_14557_, _14487_, _07766_);
  or (_14558_, _14557_, _14556_);
  and (_14559_, _05248_, _06276_);
  or (_14560_, _14559_, _14487_);
  or (_14561_, _14560_, _05886_);
  and (_14562_, _14561_, _07778_);
  and (_14563_, _14562_, _14558_);
  and (_14564_, _14563_, _14555_);
  and (_14565_, _12739_, _05248_);
  or (_14566_, _14565_, _14487_);
  and (_14567_, _14566_, _03780_);
  or (_14568_, _14567_, _14564_);
  and (_14569_, _14568_, _07777_);
  or (_14570_, _14487_, _05567_);
  and (_14571_, _14560_, _03622_);
  and (_14572_, _14571_, _14570_);
  or (_14573_, _14572_, _14569_);
  and (_14574_, _14573_, _06828_);
  and (_14575_, _14501_, _03790_);
  and (_14576_, _14575_, _14570_);
  or (_14577_, _14576_, _03624_);
  or (_14578_, _14577_, _14574_);
  nor (_14579_, _12732_, _06830_);
  or (_14580_, _14487_, _07795_);
  or (_14581_, _14580_, _14579_);
  and (_14582_, _14581_, _07793_);
  and (_14583_, _14582_, _14578_);
  nor (_14584_, _12738_, _06830_);
  or (_14585_, _14584_, _14487_);
  and (_14586_, _14585_, _03785_);
  or (_14587_, _14586_, _03815_);
  or (_14588_, _14587_, _14583_);
  or (_14589_, _14498_, _04246_);
  and (_14590_, _14589_, _03823_);
  and (_14591_, _14590_, _14588_);
  and (_14592_, _14520_, _03453_);
  or (_14593_, _14592_, _03447_);
  or (_14594_, _14593_, _14591_);
  and (_14595_, _12794_, _05248_);
  or (_14596_, _14487_, _03514_);
  or (_14597_, _14596_, _14595_);
  and (_14598_, _14597_, _43000_);
  and (_14599_, _14598_, _14594_);
  or (_14600_, _14599_, _14486_);
  and (_43485_, _14600_, _41806_);
  nor (_14601_, _43000_, _07550_);
  nor (_14602_, _05248_, _07550_);
  nor (_14603_, _12933_, _06830_);
  or (_14604_, _14603_, _14602_);
  and (_14605_, _14604_, _03222_);
  nor (_14606_, _05777_, _06830_);
  or (_14607_, _14606_, _14602_);
  or (_14608_, _14607_, _06838_);
  nor (_14609_, _05910_, _07550_);
  and (_14610_, _12827_, _05910_);
  or (_14611_, _14610_, _14609_);
  and (_14612_, _14611_, _03714_);
  nor (_14613_, _12841_, _06830_);
  or (_14614_, _14613_, _14602_);
  or (_14615_, _14614_, _04081_);
  and (_14616_, _05248_, \oc8051_golden_model_1.ACC [4]);
  or (_14617_, _14616_, _14602_);
  and (_14618_, _14617_, _04409_);
  nor (_14619_, _04409_, _07550_);
  or (_14620_, _14619_, _03610_);
  or (_14621_, _14620_, _14618_);
  and (_14622_, _14621_, _04055_);
  and (_14623_, _14622_, _14615_);
  and (_14624_, _12845_, _05910_);
  or (_14625_, _14624_, _14609_);
  and (_14626_, _14625_, _03715_);
  or (_14627_, _14626_, _03723_);
  or (_14628_, _14627_, _14623_);
  or (_14629_, _14607_, _03996_);
  and (_14630_, _14629_, _14628_);
  or (_14631_, _14630_, _03729_);
  or (_14632_, _14617_, _03737_);
  and (_14633_, _14632_, _03736_);
  and (_14634_, _14633_, _14631_);
  or (_14635_, _14634_, _14612_);
  and (_14636_, _14635_, _06840_);
  or (_14637_, _14609_, _12860_);
  and (_14638_, _14637_, _03719_);
  and (_14639_, _14638_, _14625_);
  or (_14640_, _14639_, _06869_);
  or (_14641_, _14640_, _14636_);
  nor (_14642_, _07363_, _07361_);
  nor (_14643_, _14642_, _07364_);
  or (_14644_, _14643_, _06875_);
  and (_14645_, _14644_, _03710_);
  and (_14646_, _14645_, _14641_);
  nor (_14647_, _12825_, _07391_);
  or (_14648_, _14647_, _14609_);
  and (_14649_, _14648_, _03505_);
  or (_14650_, _14649_, _07390_);
  or (_14651_, _14650_, _14646_);
  and (_14652_, _14651_, _14608_);
  or (_14653_, _14652_, _04481_);
  and (_14654_, _06730_, _05248_);
  or (_14655_, _14602_, _07400_);
  or (_14656_, _14655_, _14654_);
  and (_14657_, _14656_, _03589_);
  and (_14658_, _14657_, _14653_);
  or (_14659_, _14658_, _14605_);
  and (_14660_, _14659_, _07411_);
  or (_14661_, _14429_, _07727_);
  nor (_14662_, _14547_, _07691_);
  or (_14663_, _14662_, _07690_);
  nand (_14664_, _14663_, _07730_);
  or (_14665_, _14663_, _07730_);
  and (_14666_, _14665_, _14664_);
  or (_14667_, _14666_, _07760_);
  and (_14668_, _14667_, _07405_);
  and (_14669_, _14668_, _14661_);
  or (_14670_, _14669_, _08828_);
  or (_14671_, _14670_, _14660_);
  and (_14672_, _12821_, _05248_);
  or (_14673_, _14602_, _07766_);
  or (_14674_, _14673_, _14672_);
  and (_14675_, _06298_, _05248_);
  or (_14676_, _14675_, _14602_);
  or (_14677_, _14676_, _05886_);
  and (_14678_, _14677_, _07778_);
  and (_14679_, _14678_, _14674_);
  and (_14680_, _14679_, _14671_);
  and (_14681_, _12817_, _05248_);
  or (_14682_, _14681_, _14602_);
  and (_14683_, _14682_, _03780_);
  or (_14684_, _14683_, _14680_);
  and (_14685_, _14684_, _07777_);
  or (_14686_, _14602_, _05825_);
  and (_14687_, _14676_, _03622_);
  and (_14688_, _14687_, _14686_);
  or (_14689_, _14688_, _14685_);
  and (_14690_, _14689_, _06828_);
  and (_14691_, _14617_, _03790_);
  and (_14692_, _14691_, _14686_);
  or (_14693_, _14692_, _03624_);
  or (_14694_, _14693_, _14690_);
  nor (_14695_, _12819_, _06830_);
  or (_14696_, _14602_, _07795_);
  or (_14697_, _14696_, _14695_);
  and (_14698_, _14697_, _07793_);
  and (_14699_, _14698_, _14694_);
  nor (_14700_, _12816_, _06830_);
  or (_14701_, _14700_, _14602_);
  and (_14702_, _14701_, _03785_);
  or (_14703_, _14702_, _03815_);
  or (_14704_, _14703_, _14699_);
  or (_14705_, _14614_, _04246_);
  and (_14706_, _14705_, _03823_);
  and (_14707_, _14706_, _14704_);
  and (_14708_, _14611_, _03453_);
  or (_14709_, _14708_, _03447_);
  or (_14710_, _14709_, _14707_);
  and (_14711_, _13003_, _05248_);
  or (_14712_, _14602_, _03514_);
  or (_14713_, _14712_, _14711_);
  and (_14714_, _14713_, _43000_);
  and (_14715_, _14714_, _14710_);
  or (_14716_, _14715_, _14601_);
  and (_43486_, _14716_, _41806_);
  nor (_14717_, _43000_, _07541_);
  nor (_14718_, _05248_, _07541_);
  nor (_14719_, _13127_, _06830_);
  or (_14720_, _14719_, _14718_);
  and (_14721_, _14720_, _03222_);
  nor (_14722_, _05469_, _06830_);
  or (_14723_, _14722_, _14718_);
  or (_14724_, _14723_, _06838_);
  nor (_14725_, _05910_, _07541_);
  and (_14726_, _13047_, _05910_);
  or (_14727_, _14726_, _14725_);
  and (_14728_, _14727_, _03714_);
  nor (_14729_, _13014_, _06830_);
  or (_14730_, _14729_, _14718_);
  and (_14731_, _14730_, _03610_);
  nor (_14732_, _04409_, _07541_);
  and (_14733_, _05248_, \oc8051_golden_model_1.ACC [5]);
  or (_14734_, _14733_, _14718_);
  and (_14735_, _14734_, _04409_);
  or (_14736_, _14735_, _14732_);
  and (_14737_, _14736_, _04081_);
  or (_14738_, _14737_, _14265_);
  or (_14739_, _14738_, _14731_);
  and (_14740_, _13037_, _05910_);
  or (_14741_, _14740_, _14725_);
  or (_14742_, _14741_, _04055_);
  or (_14743_, _14723_, _03996_);
  and (_14744_, _14743_, _14742_);
  and (_14745_, _14744_, _14739_);
  or (_14746_, _14745_, _03729_);
  or (_14747_, _14734_, _03737_);
  and (_14748_, _14747_, _03736_);
  and (_14749_, _14748_, _14746_);
  or (_14750_, _14749_, _14728_);
  and (_14751_, _14750_, _06840_);
  or (_14752_, _14725_, _13054_);
  and (_14753_, _14752_, _03719_);
  and (_14754_, _14753_, _14741_);
  or (_14755_, _14754_, _06869_);
  or (_14756_, _14755_, _14751_);
  nor (_14757_, _07366_, _07068_);
  nor (_14758_, _14757_, _07367_);
  or (_14759_, _14758_, _06875_);
  and (_14760_, _14759_, _03710_);
  and (_14761_, _14760_, _14756_);
  nor (_14762_, _13020_, _07391_);
  or (_14763_, _14762_, _14725_);
  and (_14764_, _14763_, _03505_);
  or (_14765_, _14764_, _07390_);
  or (_14766_, _14765_, _14761_);
  and (_14767_, _14766_, _14724_);
  or (_14768_, _14767_, _04481_);
  and (_14769_, _06684_, _05248_);
  or (_14770_, _14718_, _07400_);
  or (_14771_, _14770_, _14769_);
  and (_14772_, _14771_, _03589_);
  and (_14773_, _14772_, _14768_);
  or (_14774_, _14773_, _14721_);
  and (_14775_, _14774_, _07411_);
  nand (_14776_, _07760_, _07737_);
  not (_14777_, _07729_);
  and (_14778_, _14664_, _14777_);
  and (_14779_, _14778_, _07740_);
  nor (_14780_, _14778_, _07740_);
  or (_14781_, _14780_, _14779_);
  or (_14782_, _14781_, _07760_);
  and (_14783_, _14782_, _07405_);
  and (_14784_, _14783_, _14776_);
  or (_14785_, _14784_, _08828_);
  or (_14786_, _14785_, _14775_);
  and (_14787_, _13141_, _05248_);
  or (_14788_, _14718_, _07766_);
  or (_14789_, _14788_, _14787_);
  and (_14790_, _06306_, _05248_);
  or (_14791_, _14790_, _14718_);
  or (_14792_, _14791_, _05886_);
  and (_14793_, _14792_, _07778_);
  and (_14794_, _14793_, _14789_);
  and (_14795_, _14794_, _14786_);
  and (_14796_, _13147_, _05248_);
  or (_14797_, _14796_, _14718_);
  and (_14798_, _14797_, _03780_);
  or (_14799_, _14798_, _14795_);
  and (_14800_, _14799_, _07777_);
  or (_14801_, _14718_, _05518_);
  and (_14802_, _14791_, _03622_);
  and (_14803_, _14802_, _14801_);
  or (_14804_, _14803_, _14800_);
  and (_14805_, _14804_, _06828_);
  and (_14806_, _14734_, _03790_);
  and (_14807_, _14806_, _14801_);
  or (_14808_, _14807_, _03624_);
  or (_14809_, _14808_, _14805_);
  nor (_14810_, _13140_, _06830_);
  or (_14811_, _14718_, _07795_);
  or (_14812_, _14811_, _14810_);
  and (_14813_, _14812_, _07793_);
  and (_14814_, _14813_, _14809_);
  nor (_14815_, _13146_, _06830_);
  or (_14816_, _14815_, _14718_);
  and (_14817_, _14816_, _03785_);
  or (_14818_, _14817_, _03815_);
  or (_14819_, _14818_, _14814_);
  or (_14820_, _14730_, _04246_);
  and (_14821_, _14820_, _03823_);
  and (_14822_, _14821_, _14819_);
  and (_14823_, _14727_, _03453_);
  or (_14824_, _14823_, _03447_);
  or (_14825_, _14824_, _14822_);
  and (_14826_, _13199_, _05248_);
  or (_14827_, _14718_, _03514_);
  or (_14828_, _14827_, _14826_);
  and (_14829_, _14828_, _43000_);
  and (_14830_, _14829_, _14825_);
  or (_14831_, _14830_, _14717_);
  and (_43487_, _14831_, _41806_);
  nor (_14832_, _43000_, _07673_);
  nor (_14833_, _05248_, _07673_);
  nor (_14834_, _13332_, _06830_);
  or (_14835_, _14834_, _14833_);
  and (_14836_, _14835_, _03222_);
  nor (_14837_, _05363_, _06830_);
  or (_14838_, _14837_, _14833_);
  or (_14839_, _14838_, _06838_);
  nor (_14840_, _05910_, _07673_);
  and (_14841_, _13253_, _05910_);
  or (_14842_, _14841_, _14840_);
  and (_14843_, _14842_, _03714_);
  nor (_14844_, _13242_, _06830_);
  or (_14845_, _14844_, _14833_);
  or (_14846_, _14845_, _04081_);
  and (_14847_, _05248_, \oc8051_golden_model_1.ACC [6]);
  or (_14848_, _14847_, _14833_);
  and (_14849_, _14848_, _04409_);
  nor (_14850_, _04409_, _07673_);
  or (_14851_, _14850_, _03610_);
  or (_14852_, _14851_, _14849_);
  and (_14853_, _14852_, _04055_);
  and (_14854_, _14853_, _14846_);
  and (_14855_, _13229_, _05910_);
  or (_14856_, _14855_, _14840_);
  and (_14857_, _14856_, _03715_);
  or (_14858_, _14857_, _03723_);
  or (_14859_, _14858_, _14854_);
  or (_14860_, _14838_, _03996_);
  and (_14861_, _14860_, _14859_);
  or (_14862_, _14861_, _03729_);
  or (_14863_, _14848_, _03737_);
  and (_14864_, _14863_, _03736_);
  and (_14865_, _14864_, _14862_);
  or (_14866_, _14865_, _14843_);
  and (_14867_, _14866_, _06840_);
  or (_14868_, _14840_, _13260_);
  and (_14869_, _14868_, _03719_);
  and (_14870_, _14869_, _14856_);
  or (_14871_, _14870_, _06869_);
  or (_14872_, _14871_, _14867_);
  nor (_14873_, _07382_, _07369_);
  nor (_14874_, _14873_, _07383_);
  or (_14875_, _14874_, _06875_);
  and (_14876_, _14875_, _03710_);
  and (_14877_, _14876_, _14872_);
  nor (_14878_, _13226_, _07391_);
  or (_14879_, _14878_, _14840_);
  and (_14880_, _14879_, _03505_);
  or (_14881_, _14880_, _07390_);
  or (_14882_, _14881_, _14877_);
  and (_14883_, _14882_, _14839_);
  or (_14884_, _14883_, _04481_);
  and (_14885_, _06455_, _05248_);
  or (_14886_, _14833_, _07400_);
  or (_14887_, _14886_, _14885_);
  and (_14888_, _14887_, _03589_);
  and (_14889_, _14888_, _14884_);
  or (_14890_, _14889_, _14836_);
  and (_14891_, _14890_, _07411_);
  nor (_14892_, _14778_, _07738_);
  or (_14893_, _14892_, _07739_);
  and (_14894_, _14893_, _07721_);
  nor (_14895_, _14893_, _07721_);
  or (_14896_, _14895_, _14894_);
  or (_14897_, _14896_, _07760_);
  or (_14898_, _14429_, _07679_);
  and (_14899_, _14898_, _07405_);
  and (_14900_, _14899_, _14897_);
  or (_14901_, _14900_, _08828_);
  or (_14902_, _14901_, _14891_);
  and (_14903_, _13347_, _05248_);
  or (_14904_, _14833_, _07766_);
  or (_14905_, _14904_, _14903_);
  and (_14906_, _13339_, _05248_);
  or (_14907_, _14906_, _14833_);
  or (_14908_, _14907_, _05886_);
  and (_14909_, _14908_, _07778_);
  and (_14910_, _14909_, _14905_);
  and (_14911_, _14910_, _14902_);
  and (_14912_, _13353_, _05248_);
  or (_14913_, _14912_, _14833_);
  and (_14914_, _14913_, _03780_);
  or (_14915_, _14914_, _14911_);
  and (_14916_, _14915_, _07777_);
  or (_14917_, _14833_, _05412_);
  and (_14918_, _14907_, _03622_);
  and (_14919_, _14918_, _14917_);
  or (_14920_, _14919_, _14916_);
  and (_14921_, _14920_, _06828_);
  and (_14922_, _14848_, _03790_);
  and (_14923_, _14922_, _14917_);
  or (_14924_, _14923_, _03624_);
  or (_14925_, _14924_, _14921_);
  nor (_14926_, _13346_, _06830_);
  or (_14927_, _14833_, _07795_);
  or (_14928_, _14927_, _14926_);
  and (_14929_, _14928_, _07793_);
  and (_14930_, _14929_, _14925_);
  nor (_14931_, _13352_, _06830_);
  or (_14932_, _14931_, _14833_);
  and (_14933_, _14932_, _03785_);
  or (_14934_, _14933_, _03815_);
  or (_14935_, _14934_, _14930_);
  or (_14936_, _14845_, _04246_);
  and (_14937_, _14936_, _03823_);
  and (_14938_, _14937_, _14935_);
  and (_14939_, _14842_, _03453_);
  or (_14940_, _14939_, _03447_);
  or (_14941_, _14940_, _14938_);
  and (_14942_, _13402_, _05248_);
  or (_14943_, _14833_, _03514_);
  or (_14944_, _14943_, _14942_);
  and (_14945_, _14944_, _43000_);
  and (_14946_, _14945_, _14941_);
  or (_14947_, _14946_, _14832_);
  and (_43488_, _14947_, _41806_);
  nor (_14948_, _43000_, _03335_);
  and (_14949_, _08780_, \oc8051_golden_model_1.ACC [1]);
  nand (_14950_, _08732_, _06075_);
  nand (_14951_, _08318_, _03517_);
  and (_14952_, _14951_, _08734_);
  and (_14953_, _03605_, _03202_);
  and (_14954_, _03616_, _03202_);
  nand (_14955_, _08458_, _10057_);
  nor (_14956_, _05666_, _07908_);
  nor (_14957_, _05254_, _03335_);
  and (_14958_, _05254_, _06274_);
  nor (_14959_, _14958_, _14957_);
  nor (_14960_, _14959_, _14956_);
  and (_14961_, _14960_, _03622_);
  nor (_14962_, _04198_, _04197_);
  or (_14963_, _14962_, _08681_);
  and (_14964_, _12124_, _05254_);
  nor (_14965_, _14964_, _14957_);
  nand (_14966_, _14965_, _03600_);
  or (_14967_, _12128_, _03779_);
  and (_14968_, _14967_, _07905_);
  nand (_14969_, _04048_, _03216_);
  and (_14970_, _05254_, _04620_);
  nor (_14971_, _14970_, _14957_);
  nand (_14972_, _14971_, _07390_);
  nand (_14973_, _07974_, _07913_);
  or (_14974_, _08063_, _04620_);
  nor (_14975_, _08066_, _04422_);
  or (_14976_, _14975_, _06546_);
  and (_14977_, _08079_, _04620_);
  or (_14978_, _04064_, \oc8051_golden_model_1.ACC [0]);
  nand (_14979_, _04064_, \oc8051_golden_model_1.ACC [0]);
  and (_14980_, _14979_, _14978_);
  and (_14981_, _14980_, _08078_);
  or (_14982_, _14981_, _08066_);
  or (_14983_, _14982_, _14977_);
  and (_14984_, _14983_, _03235_);
  or (_14985_, _14984_, _04422_);
  and (_14986_, _14985_, _04081_);
  and (_14987_, _14986_, _14976_);
  nor (_14988_, _14957_, _14956_);
  nor (_14989_, _14988_, _04081_);
  or (_14990_, _14989_, _03715_);
  or (_14991_, _14990_, _14987_);
  nor (_14992_, _05903_, _03335_);
  and (_14993_, _12021_, _05903_);
  nor (_14994_, _14993_, _14992_);
  nand (_14995_, _14994_, _03715_);
  and (_14996_, _14995_, _03996_);
  and (_14997_, _14996_, _14991_);
  nor (_14998_, _14971_, _03996_);
  or (_14999_, _14998_, _08064_);
  or (_15000_, _14999_, _14997_);
  and (_15001_, _15000_, _14974_);
  or (_15002_, _15001_, _04443_);
  or (_15003_, _06546_, _08128_);
  and (_15004_, _15003_, _03737_);
  and (_15005_, _15004_, _15002_);
  nor (_15006_, _08285_, _03737_);
  or (_15007_, _15006_, _08132_);
  or (_15008_, _15007_, _15005_);
  nand (_15009_, _08132_, _07484_);
  and (_15010_, _15009_, _15008_);
  or (_15011_, _15010_, _03714_);
  or (_15012_, _14957_, _03736_);
  and (_15013_, _15012_, _06840_);
  and (_15014_, _15013_, _15011_);
  nor (_15015_, _14988_, _06840_);
  or (_15016_, _15015_, _06869_);
  or (_15017_, _15016_, _15014_);
  nand (_15018_, _03494_, _03223_);
  or (_15019_, _15018_, _12559_);
  not (_15020_, _07330_);
  nand (_15021_, _15020_, _06869_);
  and (_15022_, _15021_, _15019_);
  and (_15023_, _15022_, _08058_);
  and (_15024_, _15023_, _15017_);
  nor (_15025_, _08170_, _08059_);
  or (_15026_, _15025_, _08051_);
  or (_15027_, _15026_, _15024_);
  nor (_15028_, _08035_, _03335_);
  nor (_15029_, _15028_, _08036_);
  nand (_15030_, _08051_, _15029_);
  and (_15031_, _15030_, _03766_);
  and (_15032_, _15031_, _15027_);
  nor (_15033_, _08566_, _03335_);
  nor (_15034_, _15033_, _10217_);
  nand (_15035_, _15034_, _07914_);
  and (_15036_, _15035_, _08187_);
  or (_15037_, _15036_, _15032_);
  and (_15038_, _15037_, _14973_);
  or (_15039_, _15038_, _07912_);
  nand (_15040_, _04048_, _07912_);
  and (_15041_, _15040_, _03710_);
  and (_15042_, _15041_, _15039_);
  nor (_15043_, _12052_, _08339_);
  nor (_15044_, _15043_, _14992_);
  nor (_15045_, _15044_, _03710_);
  or (_15046_, _15045_, _07390_);
  or (_15047_, _15046_, _15042_);
  and (_15048_, _15047_, _14972_);
  or (_15049_, _15048_, _04481_);
  and (_15050_, _06546_, _05254_);
  nor (_15051_, _15050_, _14957_);
  nand (_15052_, _15051_, _04481_);
  and (_15053_, _15052_, _03589_);
  and (_15054_, _15053_, _15049_);
  nor (_15055_, _12109_, _07908_);
  nor (_15056_, _15055_, _14957_);
  nor (_15057_, _15056_, _03589_);
  or (_15058_, _15057_, _07405_);
  or (_15059_, _15058_, _15054_);
  nand (_15060_, _07760_, _07405_);
  and (_15061_, _15060_, _15059_);
  or (_15062_, _15061_, _03216_);
  and (_15063_, _15062_, _14969_);
  or (_15064_, _15063_, _03601_);
  nand (_15065_, _14959_, _03601_);
  and (_15066_, _15065_, _08364_);
  and (_15067_, _15066_, _15064_);
  nor (_15068_, _08364_, _04048_);
  or (_15069_, _15068_, _08371_);
  or (_15070_, _15069_, _15067_);
  and (_15071_, _04634_, _03335_);
  nor (_15072_, _15071_, _08681_);
  or (_15073_, _08377_, _15072_);
  and (_15074_, _15073_, _08383_);
  and (_15075_, _15074_, _15070_);
  or (_15076_, _08386_, _15072_);
  and (_15077_, _15076_, _08388_);
  or (_15078_, _15077_, _15075_);
  or (_15079_, _08394_, _15072_);
  and (_15080_, _15079_, _08393_);
  and (_15081_, _15080_, _15078_);
  nor (_15082_, _06546_, \oc8051_golden_model_1.ACC [0]);
  nor (_15083_, _15082_, _08645_);
  and (_15084_, _08392_, _15083_);
  or (_15085_, _15084_, _03778_);
  or (_15086_, _15085_, _15081_);
  and (_15087_, _15086_, _14968_);
  and (_15088_, _10058_, _07904_);
  or (_15089_, _15088_, _03600_);
  or (_15090_, _15089_, _15087_);
  and (_15091_, _15090_, _14966_);
  or (_15092_, _15091_, _03780_);
  not (_15093_, _03592_);
  and (_15094_, _08070_, _15093_);
  nor (_15095_, _15094_, _04193_);
  nor (_15096_, _15095_, _03982_);
  or (_15097_, _14957_, _07778_);
  and (_15098_, _15097_, _15096_);
  and (_15099_, _15098_, _15092_);
  nor (_15100_, _10321_, _04193_);
  not (_15101_, _15100_);
  and (_15102_, _15096_, _15101_);
  not (_15103_, _15102_);
  or (_15104_, _15100_, _08681_);
  and (_15105_, _15104_, _15103_);
  or (_15106_, _15105_, _04199_);
  or (_15107_, _15106_, _15099_);
  and (_15108_, _15107_, _14963_);
  or (_15109_, _15108_, _08420_);
  or (_15110_, _08425_, _08645_);
  and (_15111_, _15110_, _03789_);
  and (_15112_, _15111_, _15109_);
  or (_15113_, _12005_, _08429_);
  and (_15114_, _15113_, _08431_);
  or (_15115_, _15114_, _15112_);
  or (_15116_, _08435_, _08751_);
  and (_15117_, _15116_, _07777_);
  and (_15118_, _15117_, _15115_);
  or (_15119_, _15118_, _14961_);
  nor (_15120_, _07895_, _04190_);
  not (_15121_, _15120_);
  and (_15122_, _15121_, _15119_);
  nor (_15123_, _10321_, _04190_);
  nor (_15124_, _15121_, _15071_);
  or (_15125_, _15124_, _15123_);
  or (_15126_, _15125_, _15122_);
  and (_15127_, _04058_, _03200_);
  not (_15128_, _15127_);
  nand (_15129_, _15123_, _15071_);
  and (_15130_, _15129_, _15128_);
  and (_15131_, _15130_, _15126_);
  nor (_15132_, _15071_, _15128_);
  or (_15133_, _15132_, _08450_);
  or (_15134_, _15133_, _15131_);
  nand (_15135_, _08450_, _15082_);
  and (_15136_, _15135_, _03784_);
  and (_15137_, _15136_, _15134_);
  nand (_15138_, _12003_, _08461_);
  and (_15139_, _15138_, _08460_);
  or (_15140_, _15139_, _15137_);
  and (_15141_, _15140_, _14955_);
  or (_15142_, _15141_, _03624_);
  nor (_15143_, _12122_, _07908_);
  nor (_15144_, _15143_, _14957_);
  nand (_15145_, _15144_, _03624_);
  and (_15146_, _15145_, _07898_);
  and (_15147_, _15146_, _15142_);
  nor (_15148_, _08170_, _07898_);
  or (_15149_, _15148_, _08475_);
  or (_15150_, _15149_, _15147_);
  nand (_15151_, _08475_, _15029_);
  and (_15152_, _15151_, _15150_);
  or (_15153_, _15152_, _03776_);
  nand (_15154_, _15034_, _03776_);
  and (_15155_, _15154_, _08589_);
  and (_15156_, _15155_, _15153_);
  nor (_15157_, _08589_, _07974_);
  or (_15158_, _15157_, _08587_);
  or (_15159_, _15158_, _15156_);
  nand (_15160_, _08587_, _07871_);
  and (_15161_, _15160_, _08617_);
  and (_15162_, _15161_, _15159_);
  and (_15163_, _08618_, _15072_);
  nor (_15164_, _15163_, _15162_);
  or (_15165_, _15164_, _14954_);
  nand (_15166_, _14954_, _15083_);
  and (_15167_, _15166_, _15165_);
  nor (_15168_, _15167_, _14953_);
  and (_15169_, _15083_, _14953_);
  or (_15170_, _15169_, _03517_);
  or (_15171_, _15170_, _15168_);
  and (_15172_, _15171_, _14952_);
  and (_15173_, _08701_, _10058_);
  or (_15174_, _15173_, _08732_);
  or (_15175_, _15174_, _15172_);
  and (_15176_, _15175_, _14950_);
  or (_15177_, _15176_, _03815_);
  nand (_15178_, _14988_, _03815_);
  and (_15179_, _15178_, _08776_);
  and (_15180_, _15179_, _15177_);
  and (_15181_, _08775_, _03335_);
  or (_15182_, _15181_, _15180_);
  and (_15183_, _15182_, _10359_);
  or (_15184_, _15183_, _14949_);
  and (_15185_, _15184_, _03823_);
  and (_15186_, _14957_, _03453_);
  or (_15187_, _15186_, _03447_);
  or (_15188_, _15187_, _15185_);
  nand (_15189_, _14988_, _03447_);
  and (_15190_, _15189_, _08799_);
  and (_15191_, _15190_, _15188_);
  and (_15192_, _08798_, _03335_);
  or (_15193_, _15192_, _08805_);
  or (_15194_, _15193_, _15191_);
  nand (_15195_, _08805_, _03274_);
  and (_15196_, _15195_, _43000_);
  and (_15197_, _15196_, _15194_);
  or (_15198_, _15197_, _14948_);
  and (_43491_, _15198_, _41806_);
  nor (_15199_, _43000_, _03274_);
  nand (_15200_, _08732_, _03335_);
  nor (_15201_, _08645_, _08644_);
  nor (_15202_, _15201_, _08646_);
  or (_15203_, _15202_, _08624_);
  nor (_15204_, _05254_, _03274_);
  and (_15205_, _12207_, _05254_);
  nor (_15206_, _15205_, _15204_);
  nor (_15207_, _15206_, _07777_);
  and (_15208_, _12327_, _05254_);
  nor (_15209_, _15208_, _15204_);
  and (_15210_, _15209_, _03600_);
  nand (_15211_, _03414_, _03216_);
  and (_15212_, _05254_, _06764_);
  nor (_15213_, _15212_, _15204_);
  nand (_15214_, _15213_, _07390_);
  or (_15215_, _08063_, _06764_);
  or (_15216_, _08078_, _06764_);
  nor (_15217_, _04064_, _03274_);
  and (_15218_, _04064_, _03274_);
  nor (_15219_, _15218_, _15217_);
  nand (_15220_, _15219_, _08078_);
  and (_15221_, _15220_, _08067_);
  and (_15222_, _15221_, _15216_);
  or (_15223_, _15222_, _08066_);
  and (_15224_, _15223_, _03235_);
  or (_15225_, _15224_, _04422_);
  and (_15226_, _15222_, _05966_);
  or (_15227_, _15226_, _06501_);
  and (_15228_, _15227_, _15225_);
  or (_15229_, _15228_, _03610_);
  nor (_15230_, _05254_, \oc8051_golden_model_1.ACC [1]);
  and (_15231_, _12213_, _05254_);
  nor (_15232_, _15231_, _15230_);
  or (_15233_, _15232_, _04081_);
  and (_15234_, _15233_, _15229_);
  or (_15235_, _15234_, _08089_);
  nor (_15236_, _08096_, \oc8051_golden_model_1.PSW [6]);
  nor (_15237_, _15236_, \oc8051_golden_model_1.ACC [1]);
  and (_15238_, _15236_, \oc8051_golden_model_1.ACC [1]);
  nor (_15239_, _15238_, _15237_);
  nand (_15240_, _15239_, _08089_);
  and (_15241_, _15240_, _03730_);
  and (_15242_, _15241_, _15235_);
  nor (_15243_, _05903_, _03274_);
  and (_15244_, _12224_, _05903_);
  nor (_15245_, _15244_, _15243_);
  nor (_15246_, _15245_, _04055_);
  nor (_15247_, _15213_, _03996_);
  or (_15248_, _15247_, _08064_);
  or (_15249_, _15248_, _15246_);
  or (_15250_, _15249_, _15242_);
  and (_15251_, _15250_, _15215_);
  or (_15252_, _15251_, _04443_);
  or (_15253_, _06501_, _08128_);
  and (_15254_, _15253_, _03737_);
  and (_15255_, _15254_, _15252_);
  nor (_15256_, _08271_, _03737_);
  or (_15257_, _15256_, _08132_);
  or (_15258_, _15257_, _15255_);
  nand (_15259_, _08132_, _07478_);
  and (_15260_, _15259_, _15258_);
  or (_15261_, _15260_, _03714_);
  and (_15262_, _12211_, _05903_);
  nor (_15263_, _15262_, _15243_);
  nand (_15264_, _15263_, _03714_);
  and (_15265_, _15264_, _06840_);
  and (_15266_, _15265_, _15261_);
  and (_15267_, _15244_, _12239_);
  nor (_15268_, _15267_, _15243_);
  nor (_15269_, _15268_, _06840_);
  or (_15270_, _15269_, _06869_);
  or (_15271_, _15270_, _15266_);
  and (_15272_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_15273_, _15272_, _07703_);
  nor (_15274_, _15273_, _07331_);
  or (_15275_, _15274_, _06875_);
  and (_15276_, _15275_, _08059_);
  and (_15277_, _15276_, _15271_);
  and (_15278_, \oc8051_golden_model_1.PSW [7], _03335_);
  and (_15279_, _07871_, \oc8051_golden_model_1.ACC [0]);
  not (_15280_, _15279_);
  and (_15281_, _15280_, _04620_);
  nor (_15282_, _15281_, _15278_);
  and (_15283_, _15282_, _08680_);
  nor (_15284_, _15282_, _08680_);
  or (_15285_, _15284_, _15283_);
  nor (_15286_, _15285_, _08051_);
  nor (_15287_, _15286_, _11350_);
  or (_15288_, _15287_, _15277_);
  and (_15289_, _15280_, _06546_);
  nor (_15290_, _15289_, _15278_);
  and (_15291_, _15290_, _08644_);
  nor (_15292_, _15290_, _08644_);
  or (_15293_, _15292_, _15291_);
  or (_15294_, _10201_, _15293_);
  and (_15295_, _15294_, _15288_);
  or (_15296_, _15295_, _03761_);
  nor (_15297_, _08285_, _15279_);
  nor (_15298_, _15297_, _15278_);
  and (_15299_, _15298_, _08316_);
  nor (_15300_, _15298_, _08316_);
  or (_15301_, _15300_, _15299_);
  nand (_15302_, _15301_, _03761_);
  and (_15303_, _15302_, _07914_);
  and (_15304_, _15303_, _15296_);
  nor (_15305_, _15279_, _04048_);
  nor (_15306_, _15305_, _15278_);
  and (_15307_, _15306_, _08753_);
  nor (_15308_, _15306_, _08753_);
  or (_15309_, _15308_, _15307_);
  and (_15310_, _15309_, _07913_);
  or (_15311_, _15310_, _07912_);
  or (_15312_, _15311_, _15304_);
  nand (_15313_, _03414_, _07912_);
  and (_15314_, _15313_, _03710_);
  and (_15315_, _15314_, _15312_);
  nor (_15316_, _12256_, _08339_);
  nor (_15317_, _15316_, _15243_);
  nor (_15318_, _15317_, _03710_);
  or (_15319_, _15318_, _07390_);
  or (_15320_, _15319_, _15315_);
  and (_15321_, _15320_, _15214_);
  or (_15322_, _15321_, _04481_);
  and (_15323_, _06501_, _05254_);
  nor (_15324_, _15323_, _15204_);
  nand (_15325_, _15324_, _04481_);
  and (_15326_, _15325_, _03589_);
  and (_15327_, _15326_, _15322_);
  nor (_15328_, _12313_, _07908_);
  nor (_15329_, _15328_, _15204_);
  nor (_15330_, _15329_, _03589_);
  or (_15331_, _15330_, _07405_);
  or (_15332_, _15331_, _15327_);
  or (_15333_, _07668_, _07411_);
  and (_15334_, _15333_, _15332_);
  or (_15335_, _15334_, _03216_);
  and (_15336_, _15335_, _15211_);
  or (_15337_, _15336_, _03601_);
  and (_15338_, _05254_, _04303_);
  nor (_15339_, _15338_, _15230_);
  or (_15340_, _15339_, _05886_);
  and (_15341_, _15340_, _08364_);
  and (_15342_, _15341_, _15337_);
  nor (_15343_, _08364_, _03414_);
  or (_15344_, _15343_, _11344_);
  or (_15345_, _15344_, _15342_);
  or (_15346_, _11343_, _08680_);
  and (_15347_, _15346_, _08393_);
  and (_15348_, _15347_, _15345_);
  and (_15349_, _08392_, _08644_);
  or (_15350_, _15349_, _03778_);
  or (_15351_, _15350_, _15348_);
  or (_15352_, _12333_, _03779_);
  and (_15353_, _15352_, _07905_);
  nand (_15354_, _15353_, _15351_);
  nand (_15355_, _08753_, _07904_);
  and (_15356_, _15355_, _07766_);
  and (_15357_, _15356_, _15354_);
  or (_15358_, _15357_, _15210_);
  and (_15359_, _15358_, _07778_);
  nor (_15360_, _15204_, _07778_);
  or (_15361_, _15360_, _15103_);
  nor (_15362_, _15361_, _15359_);
  or (_15363_, _08678_, _04199_);
  and (_15364_, _15363_, _08421_);
  or (_15365_, _15364_, _15362_);
  and (_15366_, _04058_, _03191_);
  not (_15367_, _15366_);
  or (_15368_, _08678_, _15367_);
  and (_15369_, _15368_, _15365_);
  or (_15370_, _15369_, _08420_);
  or (_15371_, _08425_, _08642_);
  and (_15372_, _15371_, _03789_);
  and (_15373_, _15372_, _15370_);
  or (_15374_, _12331_, _08429_);
  and (_15375_, _15374_, _08431_);
  or (_15376_, _15375_, _15373_);
  or (_15377_, _08435_, _08750_);
  and (_15378_, _15377_, _07777_);
  and (_15379_, _15378_, _15376_);
  or (_15380_, _15379_, _15207_);
  and (_15381_, _15380_, _15121_);
  nor (_15382_, _15121_, _08679_);
  or (_15383_, _15382_, _15123_);
  or (_15384_, _15383_, _15381_);
  nand (_15385_, _15123_, _08679_);
  and (_15386_, _15385_, _15128_);
  and (_15387_, _15386_, _15384_);
  nor (_15388_, _08679_, _15128_);
  or (_15389_, _15388_, _08450_);
  or (_15390_, _15389_, _15387_);
  nand (_15391_, _08450_, _08643_);
  and (_15392_, _15391_, _03784_);
  and (_15393_, _15392_, _15390_);
  nor (_15394_, _12332_, _03784_);
  or (_15395_, _15394_, _08458_);
  or (_15396_, _15395_, _15393_);
  nand (_15397_, _08458_, _08752_);
  and (_15398_, _15397_, _15396_);
  or (_15399_, _15398_, _03624_);
  nor (_15400_, _12326_, _07908_);
  or (_15401_, _15400_, _15204_);
  or (_15402_, _15401_, _07795_);
  and (_15403_, _15402_, _07898_);
  and (_15404_, _15403_, _15399_);
  and (_15405_, _07875_, _07870_);
  nor (_15406_, _15405_, _07876_);
  and (_15407_, _15406_, _08468_);
  or (_15408_, _15407_, _08475_);
  or (_15409_, _15408_, _15404_);
  and (_15410_, _08487_, _08485_);
  nor (_15411_, _15410_, _08488_);
  or (_15412_, _15411_, _08477_);
  and (_15413_, _15412_, _03777_);
  and (_15414_, _15413_, _15409_);
  and (_15415_, _08568_, _08564_);
  nor (_15416_, _15415_, _08569_);
  and (_15417_, _15416_, _03776_);
  or (_15418_, _15417_, _15414_);
  and (_15419_, _15418_, _08589_);
  and (_15420_, _08598_, _07972_);
  nor (_15421_, _15420_, _08599_);
  and (_15422_, _15421_, _08506_);
  or (_15423_, _15422_, _08587_);
  or (_15424_, _15423_, _15419_);
  nand (_15425_, _08587_, _03335_);
  and (_15426_, _15425_, _08617_);
  and (_15427_, _15426_, _15424_);
  nor (_15428_, _08681_, _08680_);
  nor (_15429_, _15428_, _08682_);
  and (_15430_, _15429_, _08618_);
  or (_15431_, _15430_, _08620_);
  or (_15432_, _15431_, _15427_);
  and (_15433_, _15432_, _15203_);
  or (_15434_, _15433_, _03517_);
  and (_15435_, _08711_, _08316_);
  nor (_15436_, _15435_, _08712_);
  or (_15437_, _15436_, _03518_);
  and (_15438_, _15437_, _08734_);
  and (_15439_, _15438_, _15434_);
  nor (_15440_, _08753_, _08751_);
  nor (_15441_, _15440_, _08754_);
  and (_15442_, _15441_, _08701_);
  or (_15443_, _15442_, _08732_);
  or (_15444_, _15443_, _15439_);
  and (_15445_, _15444_, _15200_);
  or (_15446_, _15445_, _03815_);
  or (_15447_, _15232_, _04246_);
  and (_15448_, _15447_, _08776_);
  and (_15449_, _15448_, _15446_);
  nor (_15450_, _08806_, _08781_);
  nor (_15451_, _15450_, _08776_);
  or (_15452_, _15451_, _08780_);
  or (_15453_, _15452_, _15449_);
  nand (_15454_, _08780_, _07584_);
  and (_15455_, _15454_, _03823_);
  and (_15456_, _15455_, _15453_);
  nor (_15457_, _15263_, _03823_);
  or (_15458_, _15457_, _03447_);
  or (_15459_, _15458_, _15456_);
  nor (_15460_, _15231_, _15204_);
  nand (_15461_, _15460_, _03447_);
  and (_15462_, _15461_, _08799_);
  and (_15463_, _15462_, _15459_);
  and (_15464_, _15450_, _08798_);
  or (_15465_, _15464_, _08805_);
  or (_15466_, _15465_, _15463_);
  nand (_15467_, _08805_, _07584_);
  and (_15468_, _15467_, _43000_);
  and (_15469_, _15468_, _15466_);
  or (_15470_, _15469_, _15199_);
  and (_43492_, _15470_, _41806_);
  nor (_15471_, _43000_, _07584_);
  nor (_15472_, _05254_, _07584_);
  and (_15473_, _12533_, _05254_);
  nor (_15474_, _15473_, _15472_);
  nand (_15475_, _15474_, _03600_);
  not (_15476_, _04182_);
  or (_15477_, _08640_, _15476_);
  and (_15478_, _04058_, _03181_);
  nand (_15479_, _03904_, _03216_);
  nor (_15480_, _07908_, _04875_);
  nor (_15481_, _15480_, _15472_);
  nand (_15482_, _15481_, _07390_);
  nand (_15483_, _08064_, _04875_);
  or (_15484_, _14975_, _06637_);
  nor (_15485_, _08078_, _04875_);
  nor (_15486_, _04064_, _07584_);
  and (_15487_, _04064_, _07584_);
  or (_15488_, _15487_, _15486_);
  and (_15489_, _15488_, _08078_);
  or (_15490_, _15489_, _08066_);
  or (_15491_, _15490_, _15485_);
  and (_15492_, _15491_, _03235_);
  or (_15493_, _15492_, _04422_);
  and (_15494_, _15493_, _15484_);
  and (_15495_, _15494_, _04081_);
  nor (_15496_, _12416_, _07908_);
  nor (_15497_, _15496_, _15472_);
  nor (_15498_, _15497_, _04081_);
  or (_15499_, _15498_, _08089_);
  or (_15500_, _15499_, _15495_);
  nand (_15501_, _15236_, \oc8051_golden_model_1.ACC [2]);
  and (_15502_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_15503_, _15502_, _08095_);
  or (_15504_, _15503_, _15236_);
  and (_15505_, _15504_, _15501_);
  nand (_15506_, _15505_, _08089_);
  and (_15507_, _15506_, _03730_);
  and (_15508_, _15507_, _15500_);
  nor (_15509_, _05903_, _07584_);
  and (_15510_, _12411_, _05903_);
  nor (_15511_, _15510_, _15509_);
  nor (_15512_, _15511_, _04055_);
  nor (_15513_, _15481_, _03996_);
  or (_15514_, _15513_, _08064_);
  or (_15515_, _15514_, _15512_);
  or (_15516_, _15515_, _15508_);
  and (_15517_, _15516_, _15483_);
  or (_15518_, _15517_, _04443_);
  or (_15519_, _06637_, _08128_);
  and (_15520_, _15519_, _03737_);
  and (_15521_, _15520_, _15518_);
  nor (_15522_, _08260_, _03737_);
  or (_15523_, _15522_, _08132_);
  or (_15524_, _15523_, _15521_);
  nand (_15525_, _08132_, _07433_);
  and (_15526_, _15525_, _15524_);
  or (_15527_, _15526_, _03714_);
  and (_15528_, _12409_, _05903_);
  nor (_15529_, _15528_, _15509_);
  nand (_15530_, _15529_, _03714_);
  and (_15531_, _15530_, _06840_);
  and (_15532_, _15531_, _15527_);
  and (_15533_, _15510_, _12443_);
  nor (_15534_, _15533_, _15509_);
  nor (_15535_, _15534_, _06840_);
  or (_15536_, _15535_, _06869_);
  or (_15537_, _15536_, _15532_);
  nor (_15538_, _07333_, _07331_);
  nor (_15539_, _15538_, _07334_);
  or (_15540_, _15539_, _06875_);
  and (_15541_, _15540_, _15537_);
  or (_15542_, _15541_, _08060_);
  and (_15543_, _04406_, \oc8051_golden_model_1.ACC [1]);
  and (_15544_, _04620_, _03335_);
  nor (_15545_, _15544_, _08680_);
  nor (_15546_, _15545_, _15543_);
  nor (_15547_, _08676_, _15546_);
  and (_15548_, _08676_, _15546_);
  nor (_15549_, _15548_, _15547_);
  nor (_15550_, _15072_, _08680_);
  not (_15551_, _15550_);
  or (_15552_, _15551_, _15549_);
  and (_15553_, _15552_, \oc8051_golden_model_1.PSW [7]);
  nor (_15554_, _15549_, \oc8051_golden_model_1.PSW [7]);
  or (_15555_, _15554_, _15553_);
  nand (_15556_, _15551_, _15549_);
  and (_15557_, _15556_, _15555_);
  nor (_15558_, _15557_, _08051_);
  or (_15559_, _15558_, _11350_);
  and (_15560_, _15559_, _15542_);
  nor (_15561_, _06501_, _03274_);
  and (_15562_, _06546_, _03335_);
  nor (_15563_, _15562_, _08644_);
  nor (_15564_, _15563_, _15561_);
  nor (_15565_, _08640_, _15564_);
  and (_15566_, _08640_, _15564_);
  nor (_15567_, _15566_, _15565_);
  nor (_15568_, _15083_, _08644_);
  and (_15569_, _15568_, \oc8051_golden_model_1.PSW [7]);
  not (_15570_, _15569_);
  nor (_15571_, _15570_, _15567_);
  and (_15572_, _15570_, _15567_);
  nor (_15573_, _15572_, _15571_);
  nor (_15574_, _15573_, _10201_);
  or (_15575_, _15574_, _03761_);
  or (_15576_, _15575_, _15560_);
  nor (_15577_, _08290_, _08288_);
  nor (_15578_, _15577_, _08291_);
  and (_15579_, _08319_, \oc8051_golden_model_1.PSW [7]);
  not (_15580_, _15579_);
  nor (_15581_, _15580_, _15578_);
  and (_15582_, _15580_, _15578_);
  nor (_15583_, _15582_, _15581_);
  nand (_15584_, _15583_, _03761_);
  and (_15585_, _15584_, _07914_);
  and (_15586_, _15585_, _15576_);
  nor (_15587_, _04048_, \oc8051_golden_model_1.ACC [0]);
  nor (_15588_, _08753_, _15587_);
  nor (_15589_, _15588_, _10033_);
  nor (_15590_, _08748_, _15589_);
  and (_15591_, _08748_, _15589_);
  nor (_15592_, _15591_, _15590_);
  not (_15593_, _10059_);
  or (_15594_, _15593_, _15592_);
  and (_15595_, _15594_, \oc8051_golden_model_1.PSW [7]);
  nor (_15596_, _15592_, \oc8051_golden_model_1.PSW [7]);
  or (_15597_, _15596_, _15595_);
  nand (_15598_, _15593_, _15592_);
  and (_15599_, _15598_, _15597_);
  nor (_15600_, _15599_, _07914_);
  or (_15601_, _15600_, _07912_);
  or (_15602_, _15601_, _15586_);
  nand (_15603_, _03904_, _07912_);
  and (_15604_, _15603_, _03710_);
  and (_15605_, _15604_, _15602_);
  nor (_15606_, _12461_, _08339_);
  nor (_15607_, _15606_, _15509_);
  nor (_15608_, _15607_, _03710_);
  or (_15609_, _15608_, _07390_);
  or (_15610_, _15609_, _15605_);
  and (_15611_, _15610_, _15482_);
  or (_15612_, _15611_, _04481_);
  and (_15613_, _06637_, _05254_);
  nor (_15614_, _15613_, _15472_);
  nand (_15615_, _15614_, _04481_);
  and (_15616_, _15615_, _03589_);
  and (_15617_, _15616_, _15612_);
  nor (_15618_, _12519_, _07908_);
  nor (_15619_, _15618_, _15472_);
  nor (_15620_, _15619_, _03589_);
  or (_15621_, _15620_, _07405_);
  or (_15622_, _15621_, _15617_);
  or (_15623_, _07604_, _07411_);
  and (_15624_, _15623_, _15622_);
  or (_15626_, _15624_, _03216_);
  and (_15627_, _15626_, _15479_);
  or (_15628_, _15627_, _03601_);
  and (_15629_, _05254_, _06332_);
  nor (_15630_, _15629_, _15472_);
  nand (_15631_, _15630_, _03601_);
  and (_15632_, _15631_, _08364_);
  and (_15633_, _15632_, _15628_);
  nor (_15634_, _08364_, _03904_);
  or (_15635_, _15634_, _08371_);
  or (_15637_, _15635_, _15633_);
  or (_15638_, _08377_, _08676_);
  and (_15639_, _15638_, _08383_);
  and (_15640_, _15639_, _15637_);
  and (_15641_, _04488_, _03181_);
  nor (_15642_, _08383_, _08677_);
  or (_15643_, _15642_, _15641_);
  or (_15644_, _15643_, _15640_);
  nand (_15645_, _15641_, _08677_);
  and (_15646_, _15645_, _15644_);
  or (_15648_, _15646_, _15478_);
  and (_15649_, _03616_, _03181_);
  not (_15650_, _15649_);
  not (_15651_, _15478_);
  or (_15652_, _08676_, _15651_);
  and (_15653_, _15652_, _15650_);
  and (_15654_, _15653_, _15648_);
  or (_15655_, _08640_, _04182_);
  and (_15656_, _15655_, _08392_);
  or (_15657_, _15656_, _15654_);
  and (_15659_, _15657_, _15477_);
  or (_15660_, _15659_, _03778_);
  or (_15661_, _12539_, _03779_);
  and (_15662_, _15661_, _07905_);
  and (_15663_, _15662_, _15660_);
  and (_15664_, _08748_, _07904_);
  or (_15665_, _15664_, _03600_);
  or (_15666_, _15665_, _15663_);
  and (_15667_, _15666_, _15475_);
  or (_15668_, _15667_, _03780_);
  or (_15670_, _15472_, _07778_);
  and (_15671_, _15670_, _08417_);
  and (_15672_, _15671_, _15668_);
  and (_15673_, _08421_, _08674_);
  or (_15674_, _15673_, _08420_);
  or (_15675_, _15674_, _15672_);
  or (_15676_, _08425_, _08638_);
  and (_15677_, _15676_, _03789_);
  and (_15678_, _15677_, _15675_);
  and (_15679_, _12537_, _03788_);
  or (_15681_, _15679_, _08429_);
  or (_15682_, _15681_, _15678_);
  or (_15683_, _08435_, _08746_);
  and (_15684_, _15683_, _07777_);
  and (_15685_, _15684_, _15682_);
  not (_15686_, _11332_);
  or (_15687_, _15630_, _12538_);
  nor (_15688_, _15687_, _07777_);
  or (_15689_, _15688_, _15686_);
  or (_15690_, _15689_, _15685_);
  nor (_15692_, _08675_, _11333_);
  or (_15693_, _15692_, _08447_);
  and (_15694_, _15693_, _15690_);
  not (_15695_, _11333_);
  nor (_15696_, _08675_, _15695_);
  or (_15697_, _15696_, _08450_);
  or (_15698_, _15697_, _15694_);
  nand (_15699_, _08450_, _08639_);
  and (_15700_, _15699_, _03784_);
  and (_15701_, _15700_, _15698_);
  nor (_15703_, _12538_, _03784_);
  or (_15704_, _15703_, _08458_);
  or (_15705_, _15704_, _15701_);
  nand (_15706_, _08458_, _08747_);
  and (_15707_, _15706_, _15705_);
  or (_15708_, _15707_, _03624_);
  nor (_15709_, _12532_, _07908_);
  nor (_15710_, _15709_, _15472_);
  nand (_15711_, _15710_, _03624_);
  and (_15712_, _15711_, _07898_);
  and (_15714_, _15712_, _15708_);
  and (_15715_, _07877_, _07863_);
  nor (_15716_, _15715_, _07878_);
  and (_15717_, _15716_, _08468_);
  or (_15718_, _15717_, _15714_);
  and (_15719_, _15718_, _08477_);
  and (_15720_, _08489_, _08027_);
  nor (_15721_, _15720_, _08490_);
  and (_15722_, _15721_, _08475_);
  or (_15723_, _15722_, _03776_);
  or (_15725_, _15723_, _15719_);
  and (_15726_, _08570_, _08558_);
  nor (_15727_, _15726_, _08571_);
  or (_15728_, _15727_, _03777_);
  and (_15729_, _15728_, _08589_);
  and (_15730_, _15729_, _15725_);
  and (_15731_, _08600_, _07953_);
  nor (_15732_, _15731_, _08601_);
  and (_15733_, _15732_, _08506_);
  or (_15734_, _15733_, _08587_);
  or (_15736_, _15734_, _15730_);
  nand (_15737_, _08587_, _03274_);
  and (_15738_, _15737_, _08617_);
  and (_15739_, _15738_, _15736_);
  and (_15740_, _08683_, _08677_);
  nor (_15741_, _15740_, _08684_);
  and (_15742_, _15741_, _08618_);
  or (_15743_, _15742_, _08620_);
  or (_15744_, _15743_, _15739_);
  and (_15745_, _08647_, _08641_);
  nor (_15747_, _15745_, _08648_);
  or (_15748_, _15747_, _08624_);
  and (_15749_, _15748_, _03518_);
  and (_15750_, _15749_, _15744_);
  and (_15751_, _08713_, _08290_);
  nor (_15752_, _15751_, _08714_);
  or (_15753_, _15752_, _08701_);
  and (_15754_, _15753_, _08703_);
  or (_15755_, _15754_, _15750_);
  and (_15756_, _08755_, _08749_);
  nor (_15758_, _15756_, _08756_);
  or (_15759_, _15758_, _08734_);
  and (_15760_, _15759_, _08733_);
  and (_15761_, _15760_, _15755_);
  and (_15762_, _08732_, \oc8051_golden_model_1.ACC [1]);
  or (_15763_, _15762_, _03815_);
  or (_15764_, _15763_, _15761_);
  nand (_15765_, _15497_, _03815_);
  and (_15766_, _15765_, _08776_);
  and (_15767_, _15766_, _15764_);
  and (_15769_, _08095_, _03335_);
  nor (_15770_, _08781_, _07584_);
  or (_15771_, _15770_, _15769_);
  and (_15772_, _15771_, _08775_);
  or (_15773_, _15772_, _08780_);
  or (_15774_, _15773_, _15767_);
  nand (_15775_, _08780_, _07578_);
  and (_15776_, _15775_, _03823_);
  and (_15777_, _15776_, _15774_);
  nor (_15778_, _15529_, _03823_);
  or (_15780_, _15778_, _03447_);
  or (_15781_, _15780_, _15777_);
  and (_15782_, _12592_, _05254_);
  nor (_15783_, _15782_, _15472_);
  nand (_15784_, _15783_, _03447_);
  and (_15785_, _15784_, _08799_);
  and (_15786_, _15785_, _15781_);
  and (_15787_, _08806_, \oc8051_golden_model_1.ACC [2]);
  nor (_15788_, _08806_, \oc8051_golden_model_1.ACC [2]);
  nor (_15789_, _15788_, _15787_);
  nor (_15791_, _15789_, _08805_);
  nor (_15792_, _15791_, _11964_);
  or (_15793_, _15792_, _15786_);
  nand (_15794_, _08805_, _07578_);
  and (_15795_, _15794_, _43000_);
  and (_15796_, _15795_, _15793_);
  or (_15797_, _15796_, _15471_);
  and (_43493_, _15797_, _41806_);
  nor (_15798_, _43000_, _07578_);
  nor (_15799_, _08673_, _08671_);
  nor (_15800_, _08685_, _15799_);
  and (_15801_, _08685_, _15799_);
  nor (_15802_, _15801_, _15800_);
  nand (_15803_, _15802_, _08618_);
  and (_15804_, _07879_, _07857_);
  nor (_15805_, _15804_, _07880_);
  or (_15806_, _15805_, _07898_);
  nand (_15807_, _15686_, _08673_);
  and (_15808_, _15807_, _15695_);
  or (_15809_, _14962_, _08671_);
  nor (_15811_, _05254_, _07578_);
  and (_15812_, _12733_, _05254_);
  nor (_15813_, _15812_, _15811_);
  nand (_15814_, _15813_, _03600_);
  nor (_15815_, _08364_, _03581_);
  nand (_15816_, _03581_, _03216_);
  nor (_15817_, _07908_, _05005_);
  nor (_15818_, _15817_, _15811_);
  nand (_15819_, _15818_, _07390_);
  and (_15820_, _03904_, \oc8051_golden_model_1.ACC [2]);
  nor (_15822_, _15590_, _15820_);
  nor (_15823_, _10030_, _15822_);
  and (_15824_, _10030_, _15822_);
  nor (_15825_, _15824_, _15823_);
  and (_15826_, _15825_, \oc8051_golden_model_1.PSW [7]);
  nor (_15827_, _15825_, \oc8051_golden_model_1.PSW [7]);
  nor (_15828_, _15827_, _15826_);
  and (_15829_, _15828_, _15595_);
  nor (_15830_, _15828_, _15595_);
  or (_15831_, _15830_, _15829_);
  nand (_15833_, _15831_, _07913_);
  nor (_15834_, _05903_, _07578_);
  and (_15835_, _12631_, _05903_);
  and (_15836_, _15835_, _12648_);
  nor (_15837_, _15836_, _15834_);
  nor (_15838_, _15837_, _06840_);
  nand (_15839_, _08064_, _05005_);
  or (_15840_, _14975_, _06592_);
  nand (_15841_, _08079_, _05005_);
  nor (_15842_, _04064_, _07578_);
  and (_15844_, _04064_, _07578_);
  nor (_15845_, _15844_, _15842_);
  nand (_15846_, _15845_, _08078_);
  and (_15847_, _15846_, _15841_);
  or (_15848_, _15847_, _08066_);
  and (_15849_, _15848_, _03235_);
  or (_15850_, _15849_, _04422_);
  and (_15851_, _15850_, _04081_);
  and (_15852_, _15851_, _15840_);
  nor (_15853_, _12627_, _07908_);
  nor (_15855_, _15853_, _15811_);
  nor (_15856_, _15855_, _04081_);
  or (_15857_, _15856_, _08089_);
  or (_15858_, _15857_, _15852_);
  not (_15859_, \oc8051_golden_model_1.PSW [6]);
  nor (_15860_, _08095_, _15859_);
  nor (_15861_, _15860_, \oc8051_golden_model_1.ACC [3]);
  or (_15862_, _15861_, _08096_);
  nand (_15863_, _15862_, _08089_);
  and (_15864_, _15863_, _15858_);
  or (_15866_, _15864_, _03715_);
  nor (_15867_, _15835_, _15834_);
  nand (_15868_, _15867_, _03715_);
  and (_15869_, _15868_, _03996_);
  and (_15870_, _15869_, _15866_);
  nor (_15871_, _15818_, _03996_);
  or (_15872_, _15871_, _08064_);
  or (_15873_, _15872_, _15870_);
  and (_15874_, _15873_, _15839_);
  or (_15875_, _15874_, _04443_);
  or (_15877_, _06592_, _08128_);
  and (_15878_, _15877_, _03737_);
  and (_15879_, _15878_, _15875_);
  nor (_15880_, _08248_, _03737_);
  or (_15881_, _15880_, _08132_);
  or (_15882_, _15881_, _15879_);
  nand (_15883_, _08132_, _06075_);
  and (_15884_, _15883_, _15882_);
  or (_15885_, _15884_, _03714_);
  and (_15886_, _12641_, _05903_);
  nor (_15888_, _15886_, _15834_);
  nand (_15889_, _15888_, _03714_);
  and (_15890_, _15889_, _06840_);
  and (_15891_, _15890_, _15885_);
  or (_15892_, _15891_, _15838_);
  and (_15893_, _15892_, _06875_);
  nor (_15894_, _07336_, _07334_);
  nor (_15895_, _15894_, _07337_);
  nand (_15896_, _15895_, _06869_);
  nand (_15897_, _15896_, _08059_);
  or (_15899_, _15897_, _15893_);
  and (_15900_, _04875_, \oc8051_golden_model_1.ACC [2]);
  nor (_15901_, _15547_, _15900_);
  nor (_15902_, _15799_, _15901_);
  and (_15903_, _15799_, _15901_);
  nor (_15904_, _15903_, _15902_);
  and (_15905_, _15904_, \oc8051_golden_model_1.PSW [7]);
  nor (_15906_, _15904_, \oc8051_golden_model_1.PSW [7]);
  nor (_15907_, _15906_, _15905_);
  and (_15908_, _15907_, _15553_);
  nor (_15910_, _15907_, _15553_);
  or (_15911_, _15910_, _15908_);
  nand (_15912_, _15911_, _08060_);
  and (_15913_, _15912_, _15899_);
  or (_15914_, _15913_, _08051_);
  not (_15915_, _15568_);
  or (_15916_, _15915_, _15567_);
  and (_15917_, _15916_, \oc8051_golden_model_1.PSW [7]);
  nor (_15918_, _06637_, _07584_);
  nor (_15919_, _15565_, _15918_);
  nor (_15921_, _08637_, _08635_);
  nor (_15922_, _15921_, _15919_);
  and (_15923_, _15921_, _15919_);
  nor (_15924_, _15923_, _15922_);
  and (_15925_, _15924_, \oc8051_golden_model_1.PSW [7]);
  nor (_15926_, _15924_, \oc8051_golden_model_1.PSW [7]);
  nor (_15927_, _15926_, _15925_);
  and (_15928_, _15927_, _15917_);
  nor (_15929_, _15927_, _15917_);
  or (_15930_, _15929_, _15928_);
  nand (_15932_, _15930_, _08051_);
  and (_15933_, _15932_, _03766_);
  and (_15934_, _15933_, _15914_);
  nor (_15935_, _08314_, _08292_);
  and (_15936_, _08314_, _08292_);
  or (_15937_, _15936_, _15935_);
  not (_15938_, _15581_);
  and (_15939_, _15938_, _15937_);
  nor (_15940_, _15939_, _08321_);
  nand (_15941_, _15940_, _07914_);
  and (_15943_, _15941_, _08187_);
  or (_15944_, _15943_, _15934_);
  and (_15945_, _15944_, _15833_);
  or (_15946_, _15945_, _07912_);
  nand (_15947_, _03581_, _07912_);
  and (_15948_, _15947_, _03710_);
  and (_15949_, _15948_, _15946_);
  nor (_15950_, _12612_, _08339_);
  nor (_15951_, _15950_, _15834_);
  nor (_15952_, _15951_, _03710_);
  or (_15954_, _15952_, _07390_);
  or (_15955_, _15954_, _15949_);
  and (_15956_, _15955_, _15819_);
  or (_15957_, _15956_, _04481_);
  and (_15958_, _06592_, _05254_);
  nor (_15959_, _15958_, _15811_);
  nand (_15960_, _15959_, _04481_);
  and (_15961_, _15960_, _03589_);
  and (_15962_, _15961_, _15957_);
  nor (_15963_, _12718_, _07908_);
  nor (_15965_, _15963_, _15811_);
  nor (_15966_, _15965_, _03589_);
  or (_15967_, _15966_, _07405_);
  or (_15968_, _15967_, _15962_);
  or (_15969_, _07547_, _07411_);
  and (_15970_, _15969_, _15968_);
  or (_15971_, _15970_, _03216_);
  and (_15972_, _15971_, _15816_);
  or (_15973_, _15972_, _03601_);
  and (_15974_, _05254_, _06276_);
  nor (_15976_, _15974_, _15811_);
  nand (_15977_, _15976_, _03601_);
  and (_15978_, _15977_, _08364_);
  and (_15979_, _15978_, _15973_);
  or (_15980_, _15979_, _15815_);
  and (_15981_, _15980_, _11343_);
  and (_15982_, _11344_, _15799_);
  or (_15983_, _15982_, _15981_);
  and (_15984_, _15983_, _08393_);
  and (_15985_, _08392_, _15921_);
  or (_15987_, _15985_, _03778_);
  or (_15988_, _15987_, _15984_);
  or (_15989_, _12739_, _03779_);
  and (_15990_, _15989_, _07905_);
  and (_15991_, _15990_, _15988_);
  and (_15992_, _10030_, _07904_);
  or (_15993_, _15992_, _03600_);
  or (_15994_, _15993_, _15991_);
  and (_15995_, _15994_, _15814_);
  or (_15996_, _15995_, _03780_);
  or (_15998_, _15811_, _07778_);
  and (_15999_, _15998_, _15096_);
  and (_16000_, _15999_, _15996_);
  or (_16001_, _15100_, _08671_);
  and (_16002_, _16001_, _15103_);
  or (_16003_, _16002_, _04199_);
  or (_16004_, _16003_, _16000_);
  and (_16005_, _16004_, _15809_);
  or (_16006_, _16005_, _08420_);
  or (_16007_, _08425_, _08635_);
  and (_16009_, _16007_, _03789_);
  and (_16010_, _16009_, _16006_);
  or (_16011_, _12737_, _08429_);
  and (_16012_, _16011_, _08431_);
  or (_16013_, _16012_, _16010_);
  or (_16014_, _08435_, _08744_);
  and (_16015_, _16014_, _07777_);
  and (_16016_, _16015_, _16013_);
  or (_16017_, _15976_, _12738_);
  nor (_16018_, _16017_, _07777_);
  or (_16020_, _16018_, _15686_);
  or (_16021_, _16020_, _16016_);
  and (_16022_, _16021_, _15808_);
  nor (_16023_, _08673_, _15695_);
  or (_16024_, _16023_, _08450_);
  or (_16025_, _16024_, _16022_);
  nand (_16026_, _08450_, _08637_);
  and (_16027_, _16026_, _03784_);
  and (_16028_, _16027_, _16025_);
  nand (_16029_, _12738_, _08461_);
  and (_16031_, _16029_, _08460_);
  or (_16032_, _16031_, _16028_);
  nand (_16033_, _08458_, _08745_);
  and (_16034_, _16033_, _07795_);
  and (_16035_, _16034_, _16032_);
  nor (_16036_, _12732_, _07908_);
  nor (_16037_, _16036_, _15811_);
  nor (_16038_, _16037_, _07795_);
  or (_16039_, _16038_, _08468_);
  or (_16040_, _16039_, _16035_);
  and (_16042_, _16040_, _15806_);
  or (_16043_, _16042_, _08475_);
  and (_16044_, _08491_, _08022_);
  nor (_16045_, _16044_, _08492_);
  or (_16046_, _16045_, _08477_);
  and (_16047_, _16046_, _03777_);
  and (_16048_, _16047_, _16043_);
  and (_16049_, _08572_, _08552_);
  nor (_16050_, _16049_, _08573_);
  and (_16051_, _16050_, _03776_);
  or (_16053_, _16051_, _08506_);
  or (_16054_, _16053_, _16048_);
  and (_16055_, _08602_, _07948_);
  nor (_16056_, _16055_, _08603_);
  or (_16057_, _16056_, _08589_);
  and (_16058_, _16057_, _08588_);
  and (_16059_, _16058_, _16054_);
  and (_16060_, _08587_, \oc8051_golden_model_1.ACC [2]);
  or (_16061_, _16060_, _08618_);
  or (_16062_, _16061_, _16059_);
  and (_16064_, _16062_, _15803_);
  or (_16065_, _16064_, _08620_);
  nor (_16066_, _08649_, _15921_);
  and (_16067_, _08649_, _15921_);
  nor (_16068_, _16067_, _16066_);
  nand (_16069_, _16068_, _08620_);
  and (_16070_, _16069_, _03518_);
  and (_16071_, _16070_, _16065_);
  nor (_16072_, _08715_, _08314_);
  and (_16073_, _08715_, _08314_);
  nor (_16075_, _16073_, _16072_);
  and (_16076_, _16075_, _03517_);
  or (_16077_, _16076_, _08701_);
  or (_16078_, _16077_, _16071_);
  nor (_16079_, _08757_, _10030_);
  and (_16080_, _08757_, _10030_);
  nor (_16081_, _16080_, _16079_);
  nand (_16082_, _16081_, _08701_);
  and (_16083_, _16082_, _08733_);
  and (_16084_, _16083_, _16078_);
  and (_16086_, _08732_, \oc8051_golden_model_1.ACC [2]);
  or (_16087_, _16086_, _03815_);
  or (_16088_, _16087_, _16084_);
  nand (_16089_, _15855_, _03815_);
  and (_16090_, _16089_, _08776_);
  and (_16091_, _16090_, _16088_);
  nor (_16092_, _15769_, _07578_);
  or (_16093_, _16092_, _08782_);
  and (_16094_, _16093_, _08775_);
  or (_16095_, _16094_, _08780_);
  or (_16097_, _16095_, _16091_);
  nand (_16098_, _08780_, _07484_);
  and (_16099_, _16098_, _03823_);
  and (_16100_, _16099_, _16097_);
  nor (_16101_, _15888_, _03823_);
  or (_16102_, _16101_, _03447_);
  or (_16103_, _16102_, _16100_);
  and (_16104_, _12794_, _05254_);
  nor (_16105_, _16104_, _15811_);
  nand (_16106_, _16105_, _03447_);
  and (_16108_, _16106_, _08799_);
  and (_16109_, _16108_, _16103_);
  or (_16110_, _15787_, \oc8051_golden_model_1.ACC [3]);
  and (_16111_, _16110_, _08807_);
  and (_16112_, _16111_, _08798_);
  or (_16113_, _16112_, _08805_);
  or (_16114_, _16113_, _16109_);
  nand (_16115_, _08805_, _07484_);
  and (_16116_, _16115_, _43000_);
  and (_16117_, _16116_, _16114_);
  or (_16119_, _16117_, _15798_);
  and (_43494_, _16119_, _41806_);
  nor (_16120_, _43000_, _07484_);
  nand (_16121_, _08732_, _07578_);
  nor (_16122_, _05254_, _07484_);
  and (_16123_, _12821_, _05254_);
  nor (_16124_, _16123_, _16122_);
  nand (_16125_, _16124_, _03600_);
  and (_16126_, _08669_, _08381_);
  nor (_16127_, _08364_, _03486_);
  nand (_16129_, _03486_, _03216_);
  nor (_16130_, _05777_, _07908_);
  nor (_16131_, _16130_, _16122_);
  nand (_16132_, _16131_, _07390_);
  and (_16133_, _08322_, _08313_);
  nor (_16134_, _16133_, _08323_);
  nand (_16135_, _16134_, _03761_);
  and (_16136_, _16135_, _07914_);
  or (_16137_, _15928_, _15925_);
  and (_16138_, _06592_, _07578_);
  or (_16140_, _06592_, _07578_);
  and (_16141_, _16140_, _15919_);
  or (_16142_, _16141_, _16138_);
  nor (_16143_, _08634_, _16142_);
  and (_16144_, _08634_, _16142_);
  nor (_16145_, _16144_, _16143_);
  and (_16146_, _16145_, \oc8051_golden_model_1.PSW [7]);
  nor (_16147_, _16145_, \oc8051_golden_model_1.PSW [7]);
  nor (_16148_, _16147_, _16146_);
  and (_16149_, _16148_, _16137_);
  nor (_16151_, _16148_, _16137_);
  nor (_16152_, _16151_, _16149_);
  and (_16153_, _16152_, _08051_);
  nand (_16154_, _08064_, _05777_);
  or (_16155_, _08067_, _06730_);
  nor (_16156_, _08078_, _05777_);
  or (_16157_, _04064_, \oc8051_golden_model_1.ACC [4]);
  nand (_16158_, _04064_, \oc8051_golden_model_1.ACC [4]);
  and (_16159_, _16158_, _16157_);
  and (_16160_, _16159_, _08078_);
  or (_16162_, _16160_, _08066_);
  or (_16163_, _16162_, _16156_);
  and (_16164_, _16163_, _08069_);
  and (_16165_, _16164_, _16155_);
  nor (_16166_, _12841_, _07908_);
  nor (_16167_, _16166_, _16122_);
  nor (_16168_, _16167_, _04081_);
  or (_16169_, _16168_, _08089_);
  or (_16170_, _16169_, _16165_);
  nor (_16171_, _08096_, \oc8051_golden_model_1.ACC [4]);
  or (_16173_, _16171_, _08102_);
  nand (_16174_, _16173_, _08089_);
  and (_16175_, _16174_, _03730_);
  and (_16176_, _16175_, _16170_);
  nor (_16177_, _05903_, _07484_);
  and (_16178_, _12845_, _05903_);
  nor (_16179_, _16178_, _16177_);
  nor (_16180_, _16179_, _04055_);
  nor (_16181_, _16131_, _03996_);
  or (_16182_, _16181_, _08064_);
  or (_16184_, _16182_, _16180_);
  or (_16185_, _16184_, _16176_);
  and (_16186_, _16185_, _16154_);
  or (_16187_, _16186_, _04443_);
  or (_16188_, _06730_, _08128_);
  and (_16189_, _16188_, _03737_);
  and (_16190_, _16189_, _16187_);
  nor (_16191_, _08235_, _03737_);
  or (_16192_, _16191_, _08132_);
  or (_16193_, _16192_, _16190_);
  nand (_16195_, _08132_, _03335_);
  and (_16196_, _16195_, _16193_);
  or (_16197_, _16196_, _03714_);
  and (_16198_, _12827_, _05903_);
  nor (_16199_, _16198_, _16177_);
  nand (_16200_, _16199_, _03714_);
  and (_16201_, _16200_, _06840_);
  and (_16202_, _16201_, _16197_);
  and (_16203_, _16178_, _12860_);
  nor (_16204_, _16203_, _16177_);
  nor (_16206_, _16204_, _06840_);
  or (_16207_, _16206_, _06869_);
  or (_16208_, _16207_, _16202_);
  nor (_16209_, _07339_, _07337_);
  nor (_16210_, _16209_, _07340_);
  or (_16211_, _16210_, _06875_);
  and (_16212_, _16211_, _16208_);
  or (_16213_, _16212_, _08060_);
  or (_16214_, _15908_, _15905_);
  nor (_16215_, _05005_, \oc8051_golden_model_1.ACC [3]);
  nand (_16217_, _05005_, \oc8051_golden_model_1.ACC [3]);
  and (_16218_, _16217_, _15901_);
  or (_16219_, _16218_, _16215_);
  nor (_16220_, _08669_, _16219_);
  and (_16221_, _08669_, _16219_);
  nor (_16222_, _16221_, _16220_);
  and (_16223_, _16222_, \oc8051_golden_model_1.PSW [7]);
  nor (_16224_, _16222_, \oc8051_golden_model_1.PSW [7]);
  nor (_16225_, _16224_, _16223_);
  and (_16226_, _16225_, _16214_);
  nor (_16228_, _16225_, _16214_);
  nor (_16229_, _16228_, _16226_);
  or (_16230_, _16229_, _08059_);
  and (_16231_, _16230_, _10201_);
  and (_16232_, _16231_, _16213_);
  or (_16233_, _16232_, _03761_);
  or (_16234_, _16233_, _16153_);
  and (_16235_, _16234_, _16136_);
  or (_16236_, _15829_, _15826_);
  or (_16237_, _15822_, _10039_);
  and (_16239_, _16237_, _10038_);
  nor (_16240_, _08743_, _16239_);
  and (_16241_, _08743_, _16239_);
  nor (_16242_, _16241_, _16240_);
  and (_16243_, _16242_, \oc8051_golden_model_1.PSW [7]);
  nor (_16244_, _16242_, \oc8051_golden_model_1.PSW [7]);
  nor (_16245_, _16244_, _16243_);
  and (_16246_, _16245_, _16236_);
  nor (_16247_, _16245_, _16236_);
  nor (_16248_, _16247_, _16246_);
  and (_16250_, _16248_, _07913_);
  or (_16251_, _16250_, _07912_);
  or (_16252_, _16251_, _16235_);
  nand (_16253_, _03486_, _07912_);
  and (_16254_, _16253_, _03710_);
  and (_16255_, _16254_, _16252_);
  nor (_16256_, _12825_, _08339_);
  nor (_16257_, _16256_, _16177_);
  nor (_16258_, _16257_, _03710_);
  or (_16259_, _16258_, _07390_);
  or (_16261_, _16259_, _16255_);
  and (_16262_, _16261_, _16132_);
  or (_16263_, _16262_, _04481_);
  and (_16264_, _06730_, _05254_);
  nor (_16265_, _16264_, _16122_);
  nand (_16266_, _16265_, _04481_);
  and (_16267_, _16266_, _03589_);
  and (_16268_, _16267_, _16263_);
  nor (_16269_, _12933_, _07908_);
  nor (_16270_, _16269_, _16122_);
  nor (_16272_, _16270_, _03589_);
  or (_16273_, _16272_, _07405_);
  or (_16274_, _16273_, _16268_);
  or (_16275_, _07493_, _07411_);
  and (_16276_, _16275_, _16274_);
  or (_16277_, _16276_, _03216_);
  and (_16278_, _16277_, _16129_);
  or (_16279_, _16278_, _03601_);
  and (_16280_, _06298_, _05254_);
  nor (_16281_, _16280_, _16122_);
  nand (_16283_, _16281_, _03601_);
  and (_16284_, _16283_, _08364_);
  and (_16285_, _16284_, _16279_);
  or (_16286_, _16285_, _16127_);
  and (_16287_, _16286_, _08377_);
  and (_16288_, _08371_, _08669_);
  or (_16289_, _16288_, _08380_);
  or (_16290_, _16289_, _16287_);
  not (_16291_, _08381_);
  and (_16292_, _08669_, _16291_);
  or (_16294_, _16292_, _08382_);
  and (_16295_, _16294_, _16290_);
  or (_16296_, _16295_, _16126_);
  and (_16297_, _16296_, _08387_);
  nor (_16298_, _08387_, _08670_);
  or (_16299_, _16298_, _15649_);
  or (_16300_, _16299_, _16297_);
  or (_16301_, _15650_, _08634_);
  and (_16302_, _16301_, _15476_);
  and (_16303_, _16302_, _16300_);
  and (_16305_, _08634_, _04182_);
  or (_16306_, _16305_, _03778_);
  or (_16307_, _16306_, _16303_);
  or (_16308_, _12817_, _03779_);
  and (_16309_, _16308_, _07905_);
  and (_16310_, _16309_, _16307_);
  and (_16311_, _08743_, _07904_);
  or (_16312_, _16311_, _03600_);
  or (_16313_, _16312_, _16310_);
  and (_16314_, _16313_, _16125_);
  or (_16316_, _16314_, _03780_);
  or (_16317_, _16122_, _07778_);
  and (_16318_, _16317_, _08417_);
  and (_16319_, _16318_, _16316_);
  and (_16320_, _08421_, _08667_);
  or (_16321_, _16320_, _08420_);
  or (_16322_, _16321_, _16319_);
  or (_16323_, _08425_, _08632_);
  and (_16324_, _16323_, _03789_);
  and (_16325_, _16324_, _16322_);
  or (_16327_, _12815_, _08429_);
  and (_16328_, _16327_, _08431_);
  or (_16329_, _16328_, _16325_);
  or (_16330_, _08435_, _08741_);
  and (_16331_, _16330_, _07777_);
  and (_16332_, _16331_, _16329_);
  or (_16333_, _16281_, _12816_);
  nor (_16334_, _16333_, _07777_);
  or (_16335_, _16334_, _08446_);
  or (_16336_, _16335_, _16332_);
  nand (_16338_, _08446_, _08668_);
  and (_16339_, _16338_, _16336_);
  or (_16340_, _16339_, _08450_);
  nand (_16341_, _08450_, _08633_);
  and (_16342_, _16341_, _03784_);
  and (_16343_, _16342_, _16340_);
  nor (_16344_, _12816_, _03784_);
  or (_16345_, _16344_, _08458_);
  or (_16346_, _16345_, _16343_);
  nand (_16347_, _08458_, _08742_);
  and (_16349_, _16347_, _16346_);
  or (_16350_, _16349_, _03624_);
  nor (_16351_, _12819_, _07908_);
  nor (_16352_, _16351_, _16122_);
  nand (_16353_, _16352_, _03624_);
  and (_16354_, _16353_, _07898_);
  and (_16355_, _16354_, _16350_);
  and (_16356_, _07881_, _07847_);
  nor (_16357_, _16356_, _07882_);
  and (_16358_, _16357_, _08468_);
  or (_16360_, _16358_, _08475_);
  or (_16361_, _16360_, _16355_);
  and (_16362_, _08493_, _08014_);
  nor (_16363_, _16362_, _08494_);
  or (_16364_, _16363_, _08477_);
  and (_16365_, _16364_, _16361_);
  or (_16366_, _16365_, _03776_);
  and (_16367_, _08574_, _08546_);
  nor (_16368_, _16367_, _08575_);
  or (_16369_, _16368_, _03777_);
  and (_16371_, _16369_, _08589_);
  and (_16372_, _16371_, _16366_);
  and (_16373_, _08604_, _07941_);
  nor (_16374_, _16373_, _08605_);
  and (_16375_, _16374_, _08506_);
  or (_16376_, _16375_, _08587_);
  or (_16377_, _16376_, _16372_);
  nand (_16378_, _08587_, _07578_);
  and (_16379_, _16378_, _08617_);
  and (_16380_, _16379_, _16377_);
  and (_16382_, _08687_, _08670_);
  nor (_16383_, _16382_, _08688_);
  and (_16384_, _16383_, _08618_);
  or (_16385_, _16384_, _16380_);
  and (_16386_, _16385_, _08624_);
  nor (_16387_, _08651_, _08634_);
  nor (_16388_, _16387_, _08652_);
  and (_16389_, _16388_, _08620_);
  or (_16390_, _16389_, _03517_);
  or (_16391_, _16390_, _16386_);
  nor (_16393_, _08719_, _08707_);
  nor (_16394_, _16393_, _08720_);
  or (_16395_, _16394_, _03518_);
  and (_16396_, _16395_, _08734_);
  and (_16397_, _16396_, _16391_);
  nor (_16398_, _08759_, _08743_);
  nor (_16399_, _16398_, _08760_);
  and (_16400_, _16399_, _08701_);
  or (_16401_, _16400_, _08732_);
  or (_16402_, _16401_, _16397_);
  and (_16404_, _16402_, _16121_);
  or (_16405_, _16404_, _03815_);
  nand (_16406_, _16167_, _03815_);
  and (_16407_, _16406_, _08776_);
  and (_16408_, _16407_, _16405_);
  and (_16409_, _08782_, _07484_);
  nor (_16410_, _08782_, _07484_);
  nor (_16411_, _16410_, _16409_);
  not (_16412_, _16411_);
  and (_16413_, _16412_, _08775_);
  or (_16415_, _16413_, _08780_);
  or (_16416_, _16415_, _16408_);
  nand (_16417_, _08780_, _07478_);
  and (_16418_, _16417_, _03823_);
  and (_16419_, _16418_, _16416_);
  nor (_16420_, _16199_, _03823_);
  or (_16421_, _16420_, _03447_);
  or (_16422_, _16421_, _16419_);
  and (_16423_, _13003_, _05254_);
  nor (_16424_, _16423_, _16122_);
  nand (_16426_, _16424_, _03447_);
  and (_16427_, _16426_, _08799_);
  and (_16428_, _16427_, _16422_);
  and (_16429_, _08807_, _07484_);
  nor (_16430_, _16429_, _08808_);
  and (_16431_, _16430_, _08798_);
  or (_16432_, _16431_, _08805_);
  or (_16433_, _16432_, _16428_);
  nand (_16434_, _08805_, _07478_);
  and (_16435_, _16434_, _43000_);
  and (_16437_, _16435_, _16433_);
  or (_16438_, _16437_, _16120_);
  and (_43495_, _16438_, _41806_);
  nor (_16439_, _43000_, _07478_);
  nor (_16440_, _05254_, _07478_);
  nor (_16441_, _13140_, _07908_);
  nor (_16442_, _16441_, _16440_);
  nor (_16443_, _16442_, _07795_);
  and (_16444_, _06306_, _05254_);
  nor (_16445_, _16444_, _16440_);
  or (_16447_, _16445_, _13146_);
  nor (_16448_, _16447_, _07777_);
  and (_16449_, _13141_, _05254_);
  nor (_16450_, _16449_, _16440_);
  nand (_16451_, _16450_, _03600_);
  or (_16452_, _08630_, _15476_);
  nor (_16453_, _08665_, _08666_);
  nor (_16454_, _15641_, _04181_);
  and (_16455_, _16454_, _08382_);
  and (_16456_, _16455_, _08377_);
  or (_16458_, _16456_, _16453_);
  nand (_16459_, _03860_, _03216_);
  nor (_16460_, _05469_, _07908_);
  nor (_16461_, _16460_, _16440_);
  nand (_16462_, _16461_, _07390_);
  and (_16463_, _03486_, \oc8051_golden_model_1.ACC [4]);
  nor (_16464_, _16240_, _16463_);
  nor (_16465_, _10026_, _16464_);
  and (_16466_, _10026_, _16464_);
  nor (_16467_, _16466_, _16465_);
  and (_16469_, _16467_, \oc8051_golden_model_1.PSW [7]);
  nor (_16470_, _16467_, \oc8051_golden_model_1.PSW [7]);
  nor (_16471_, _16470_, _16469_);
  nor (_16472_, _16246_, _16243_);
  not (_16473_, _16472_);
  and (_16474_, _16473_, _16471_);
  nor (_16475_, _16473_, _16471_);
  nor (_16476_, _16475_, _16474_);
  or (_16477_, _16476_, _07914_);
  nor (_16478_, _05903_, _07478_);
  and (_16480_, _13037_, _05903_);
  and (_16481_, _16480_, _13054_);
  nor (_16482_, _16481_, _16478_);
  nor (_16483_, _16482_, _06840_);
  nand (_16484_, _08064_, _05469_);
  or (_16485_, _08067_, _06684_);
  nor (_16486_, _08078_, _05469_);
  and (_16487_, _04064_, _07478_);
  nor (_16488_, _04064_, _07478_);
  or (_16489_, _16488_, _16487_);
  and (_16491_, _16489_, _08078_);
  or (_16492_, _16491_, _08066_);
  or (_16493_, _16492_, _16486_);
  and (_16494_, _16493_, _08069_);
  and (_16495_, _16494_, _16485_);
  nor (_16496_, _13014_, _07908_);
  nor (_16497_, _16496_, _16440_);
  nor (_16498_, _16497_, _04081_);
  or (_16499_, _16498_, _08089_);
  or (_16500_, _16499_, _16495_);
  and (_16502_, _09893_, _08104_);
  nor (_16503_, _09893_, _08104_);
  nor (_16504_, _16503_, _16502_);
  nand (_16505_, _16504_, _08089_);
  and (_16506_, _16505_, _16500_);
  or (_16507_, _16506_, _03715_);
  nor (_16508_, _16480_, _16478_);
  nand (_16509_, _16508_, _03715_);
  and (_16510_, _16509_, _03996_);
  and (_16511_, _16510_, _16507_);
  nor (_16513_, _16461_, _03996_);
  or (_16514_, _16513_, _08064_);
  or (_16515_, _16514_, _16511_);
  and (_16516_, _16515_, _16484_);
  or (_16517_, _16516_, _04443_);
  or (_16518_, _06684_, _08128_);
  and (_16519_, _16518_, _03737_);
  and (_16520_, _16519_, _16517_);
  nor (_16521_, _08218_, _03737_);
  or (_16522_, _16521_, _08132_);
  or (_16524_, _16522_, _16520_);
  nand (_16525_, _08132_, _03274_);
  and (_16526_, _16525_, _16524_);
  or (_16527_, _16526_, _03714_);
  and (_16528_, _13047_, _05903_);
  nor (_16529_, _16528_, _16478_);
  nand (_16530_, _16529_, _03714_);
  and (_16531_, _16530_, _06840_);
  and (_16532_, _16531_, _16527_);
  or (_16533_, _16532_, _16483_);
  and (_16535_, _16533_, _06875_);
  nor (_16536_, _07342_, _07340_);
  nor (_16537_, _16536_, _07343_);
  and (_16538_, _16537_, _06869_);
  or (_16539_, _16538_, _10170_);
  or (_16540_, _16539_, _16535_);
  and (_16541_, _05777_, \oc8051_golden_model_1.ACC [4]);
  nor (_16542_, _16220_, _16541_);
  nor (_16543_, _16453_, _16542_);
  and (_16544_, _16453_, _16542_);
  nor (_16546_, _16544_, _16543_);
  and (_16547_, _16546_, \oc8051_golden_model_1.PSW [7]);
  nor (_16548_, _16546_, \oc8051_golden_model_1.PSW [7]);
  nor (_16549_, _16548_, _16547_);
  nor (_16550_, _16226_, _16223_);
  not (_16551_, _16550_);
  and (_16552_, _16551_, _16549_);
  nor (_16553_, _16551_, _16549_);
  nor (_16554_, _16553_, _16552_);
  or (_16555_, _16554_, _08058_);
  and (_16558_, _16555_, _08054_);
  and (_16559_, _16558_, _16540_);
  and (_16560_, _16554_, _08053_);
  or (_16561_, _16560_, _08051_);
  or (_16562_, _16561_, _16559_);
  nor (_16563_, _06730_, _07484_);
  nor (_16564_, _16143_, _16563_);
  nor (_16565_, _08630_, _16564_);
  and (_16566_, _08630_, _16564_);
  nor (_16567_, _16566_, _16565_);
  and (_16569_, _16567_, \oc8051_golden_model_1.PSW [7]);
  nor (_16570_, _16567_, \oc8051_golden_model_1.PSW [7]);
  nor (_16571_, _16570_, _16569_);
  nor (_16572_, _16149_, _16146_);
  not (_16573_, _16572_);
  and (_16574_, _16573_, _16571_);
  nor (_16575_, _16573_, _16571_);
  nor (_16576_, _16575_, _16574_);
  or (_16577_, _16576_, _10201_);
  and (_16578_, _16577_, _03766_);
  and (_16580_, _16578_, _16562_);
  and (_16581_, _08324_, _08311_);
  nor (_16582_, _16581_, _08325_);
  nor (_16583_, _16582_, _03766_);
  or (_16584_, _16583_, _07913_);
  or (_16585_, _16584_, _16580_);
  and (_16586_, _16585_, _16477_);
  or (_16587_, _16586_, _07912_);
  nand (_16588_, _03860_, _07912_);
  and (_16589_, _16588_, _03710_);
  and (_16591_, _16589_, _16587_);
  nor (_16592_, _13020_, _08339_);
  nor (_16593_, _16592_, _16478_);
  nor (_16594_, _16593_, _03710_);
  or (_16595_, _16594_, _07390_);
  or (_16596_, _16595_, _16591_);
  and (_16597_, _16596_, _16462_);
  or (_16598_, _16597_, _04481_);
  and (_16599_, _06684_, _05254_);
  nor (_16600_, _16599_, _16440_);
  nand (_16602_, _16600_, _04481_);
  and (_16603_, _16602_, _03589_);
  and (_16604_, _16603_, _16598_);
  nor (_16605_, _13127_, _07908_);
  nor (_16606_, _16605_, _16440_);
  nor (_16607_, _16606_, _03589_);
  or (_16608_, _16607_, _07405_);
  or (_16609_, _16608_, _16604_);
  or (_16610_, _07463_, _07411_);
  and (_16611_, _16610_, _16609_);
  or (_16613_, _16611_, _03216_);
  and (_16614_, _16613_, _16459_);
  or (_16615_, _16614_, _03601_);
  nand (_16616_, _16445_, _03601_);
  and (_16617_, _16616_, _08364_);
  and (_16618_, _16617_, _16615_);
  or (_16619_, _08364_, _03860_);
  nand (_16620_, _16619_, _16456_);
  or (_16621_, _16620_, _16618_);
  and (_16622_, _16621_, _16458_);
  or (_16624_, _16622_, _15478_);
  or (_16625_, _16453_, _15651_);
  and (_16626_, _16625_, _15650_);
  and (_16627_, _16626_, _16624_);
  or (_16628_, _08630_, _04182_);
  and (_16629_, _16628_, _08392_);
  or (_16630_, _16629_, _16627_);
  and (_16631_, _16630_, _16452_);
  or (_16632_, _16631_, _03778_);
  or (_16633_, _13147_, _03779_);
  and (_16635_, _16633_, _07905_);
  and (_16636_, _16635_, _16632_);
  and (_16637_, _10026_, _07904_);
  or (_16638_, _16637_, _03600_);
  or (_16639_, _16638_, _16636_);
  and (_16640_, _16639_, _16451_);
  or (_16641_, _16640_, _03780_);
  or (_16642_, _16440_, _07778_);
  and (_16643_, _16642_, _08417_);
  and (_16644_, _16643_, _16641_);
  and (_16646_, _08421_, _08665_);
  or (_16647_, _16646_, _08420_);
  or (_16648_, _16647_, _16644_);
  or (_16649_, _08425_, _08628_);
  and (_16650_, _16649_, _03789_);
  and (_16651_, _16650_, _16648_);
  or (_16652_, _13145_, _08429_);
  and (_16653_, _16652_, _08431_);
  or (_16654_, _16653_, _16651_);
  or (_16655_, _08435_, _08739_);
  and (_16657_, _16655_, _07777_);
  and (_16658_, _16657_, _16654_);
  or (_16659_, _16658_, _16448_);
  and (_16660_, _16659_, _15121_);
  nor (_16661_, _15121_, _08666_);
  or (_16662_, _16661_, _15123_);
  or (_16663_, _16662_, _16660_);
  nand (_16664_, _15123_, _08666_);
  and (_16665_, _16664_, _15128_);
  and (_16666_, _16665_, _16663_);
  nor (_16668_, _08666_, _15128_);
  or (_16669_, _16668_, _08450_);
  or (_16670_, _16669_, _16666_);
  nand (_16671_, _08450_, _08629_);
  and (_16672_, _16671_, _03784_);
  and (_16673_, _16672_, _16670_);
  nor (_16674_, _13146_, _03784_);
  or (_16675_, _16674_, _08458_);
  or (_16676_, _16675_, _16673_);
  nand (_16677_, _08458_, _08740_);
  and (_16679_, _16677_, _07795_);
  and (_16680_, _16679_, _16676_);
  or (_16681_, _16680_, _16443_);
  and (_16682_, _16681_, _07898_);
  and (_16683_, _07883_, _07841_);
  nor (_16684_, _16683_, _07884_);
  and (_16685_, _16684_, _08468_);
  or (_16686_, _16685_, _08475_);
  or (_16687_, _16686_, _16682_);
  and (_16688_, _08495_, _08012_);
  nor (_16690_, _16688_, _08496_);
  or (_16691_, _16690_, _08477_);
  and (_16692_, _16691_, _03777_);
  and (_16693_, _16692_, _16687_);
  and (_16694_, _08576_, _08540_);
  nor (_16695_, _16694_, _08577_);
  or (_16696_, _16695_, _08506_);
  and (_16697_, _16696_, _08508_);
  or (_16698_, _16697_, _16693_);
  and (_16699_, _08606_, _07939_);
  nor (_16701_, _16699_, _08607_);
  or (_16702_, _16701_, _08589_);
  and (_16703_, _16702_, _08588_);
  and (_16704_, _16703_, _16698_);
  not (_16705_, _04226_);
  and (_16706_, _10320_, _16705_);
  nand (_16707_, _08587_, \oc8051_golden_model_1.ACC [4]);
  nand (_16708_, _16707_, _16706_);
  or (_16709_, _16708_, _16704_);
  and (_16710_, _03494_, _03202_);
  not (_16712_, _16710_);
  nor (_16713_, _08689_, _16453_);
  and (_16714_, _08689_, _16453_);
  or (_16715_, _16714_, _16713_);
  or (_16716_, _16715_, _16706_);
  and (_16717_, _16716_, _16712_);
  and (_16718_, _16717_, _16709_);
  and (_16719_, _16715_, _16710_);
  or (_16720_, _16719_, _08620_);
  or (_16721_, _16720_, _16718_);
  and (_16723_, _08653_, _08631_);
  nor (_16724_, _16723_, _08654_);
  or (_16725_, _16724_, _08624_);
  and (_16726_, _16725_, _03518_);
  and (_16727_, _16726_, _16721_);
  and (_16728_, _08721_, _08308_);
  nor (_16729_, _16728_, _08722_);
  or (_16730_, _16729_, _08701_);
  and (_16731_, _16730_, _08703_);
  or (_16732_, _16731_, _16727_);
  not (_16734_, _10026_);
  nor (_16735_, _08761_, _16734_);
  and (_16736_, _08761_, _16734_);
  nor (_16737_, _16736_, _16735_);
  or (_16738_, _16737_, _08734_);
  and (_16739_, _16738_, _08733_);
  and (_16740_, _16739_, _16732_);
  and (_16741_, _08732_, \oc8051_golden_model_1.ACC [4]);
  or (_16742_, _16741_, _03815_);
  or (_16743_, _16742_, _16740_);
  nand (_16745_, _16497_, _03815_);
  and (_16746_, _16745_, _08776_);
  and (_16747_, _16746_, _16743_);
  nor (_16748_, _16409_, _07478_);
  or (_16749_, _16748_, _08783_);
  and (_16750_, _16749_, _08775_);
  or (_16751_, _16750_, _08780_);
  or (_16752_, _16751_, _16747_);
  nand (_16753_, _08780_, _07433_);
  and (_16754_, _16753_, _03823_);
  and (_16756_, _16754_, _16752_);
  nor (_16757_, _16529_, _03823_);
  or (_16758_, _16757_, _03447_);
  or (_16759_, _16758_, _16756_);
  and (_16760_, _13199_, _05254_);
  nor (_16761_, _16760_, _16440_);
  nand (_16762_, _16761_, _03447_);
  and (_16763_, _16762_, _08799_);
  and (_16764_, _16763_, _16759_);
  nor (_16765_, _08808_, \oc8051_golden_model_1.ACC [5]);
  nor (_16767_, _16765_, _08809_);
  nor (_16768_, _16767_, _08805_);
  nor (_16769_, _16768_, _11964_);
  or (_16770_, _16769_, _16764_);
  nand (_16771_, _08805_, _07433_);
  and (_16772_, _16771_, _43000_);
  and (_16773_, _16772_, _16770_);
  or (_16774_, _16773_, _16439_);
  and (_43496_, _16774_, _41806_);
  nor (_16775_, _43000_, _07433_);
  nand (_16777_, _08732_, _07478_);
  nor (_16778_, _05254_, _07433_);
  and (_16779_, _13339_, _05254_);
  nor (_16780_, _16779_, _16778_);
  or (_16781_, _16780_, _13352_);
  nor (_16782_, _16781_, _07777_);
  and (_16783_, _13347_, _05254_);
  nor (_16784_, _16783_, _16778_);
  nand (_16785_, _16784_, _03600_);
  and (_16786_, _08387_, _16291_);
  not (_16788_, _16786_);
  and (_16789_, _16788_, _08664_);
  or (_16790_, _08377_, _08664_);
  nand (_16791_, _03549_, _03216_);
  nor (_16792_, _05363_, _07908_);
  nor (_16793_, _16792_, _16778_);
  nand (_16794_, _16793_, _07390_);
  and (_16795_, _08326_, _08307_);
  nor (_16796_, _16795_, _08327_);
  nand (_16797_, _16796_, _03761_);
  and (_16799_, _16797_, _07914_);
  or (_16800_, _06684_, _07478_);
  and (_16801_, _06684_, _07478_);
  or (_16802_, _16564_, _16801_);
  and (_16803_, _16802_, _16800_);
  nor (_16804_, _16803_, _08627_);
  and (_16805_, _16803_, _08627_);
  nor (_16806_, _16805_, _16804_);
  nor (_16807_, _16574_, _16569_);
  and (_16808_, _16807_, \oc8051_golden_model_1.PSW [7]);
  nor (_16810_, _16808_, _16806_);
  and (_16811_, _16808_, _16806_);
  nor (_16812_, _16811_, _16810_);
  and (_16813_, _16812_, _08051_);
  nand (_16814_, _08064_, _05363_);
  nor (_16815_, _13242_, _07908_);
  nor (_16816_, _16815_, _16778_);
  nor (_16817_, _16816_, _04081_);
  or (_16818_, _08067_, _06455_);
  nor (_16819_, _08078_, _05363_);
  and (_16821_, _04064_, _07433_);
  nor (_16822_, _04064_, _07433_);
  or (_16823_, _16822_, _16821_);
  and (_16824_, _16823_, _08078_);
  or (_16825_, _16824_, _08066_);
  or (_16826_, _16825_, _16819_);
  and (_16827_, _16826_, _08069_);
  and (_16828_, _16827_, _16818_);
  or (_16829_, _16828_, _16817_);
  and (_16830_, _16829_, _09882_);
  not (_16832_, _08106_);
  nor (_16833_, _16503_, _16832_);
  and (_16834_, _09892_, _08107_);
  nor (_16835_, _16834_, _16833_);
  nor (_16836_, _16835_, _09882_);
  or (_16837_, _16836_, _03715_);
  or (_16838_, _16837_, _16830_);
  nor (_16839_, _05903_, _07433_);
  and (_16840_, _13229_, _05903_);
  nor (_16841_, _16840_, _16839_);
  nand (_16843_, _16841_, _03715_);
  and (_16844_, _16843_, _03996_);
  and (_16845_, _16844_, _16838_);
  nor (_16846_, _16793_, _03996_);
  or (_16847_, _16846_, _08064_);
  or (_16848_, _16847_, _16845_);
  and (_16849_, _16848_, _16814_);
  or (_16850_, _16849_, _04443_);
  or (_16851_, _06455_, _08128_);
  and (_16852_, _16851_, _03737_);
  and (_16854_, _16852_, _16850_);
  nor (_16855_, _08203_, _03737_);
  or (_16856_, _16855_, _08132_);
  or (_16857_, _16856_, _16854_);
  nand (_16858_, _08132_, _07584_);
  and (_16859_, _16858_, _16857_);
  or (_16860_, _16859_, _03714_);
  and (_16861_, _13253_, _05903_);
  nor (_16862_, _16861_, _16839_);
  nand (_16863_, _16862_, _03714_);
  and (_16865_, _16863_, _06840_);
  and (_16866_, _16865_, _16860_);
  and (_16867_, _16840_, _13260_);
  nor (_16868_, _16867_, _16839_);
  nor (_16869_, _16868_, _06840_);
  or (_16870_, _16869_, _06869_);
  or (_16871_, _16870_, _16866_);
  nor (_16872_, _07345_, _07343_);
  nor (_16873_, _16872_, _07346_);
  or (_16874_, _16873_, _06875_);
  and (_16876_, _16874_, _16871_);
  or (_16877_, _16876_, _08060_);
  nand (_16878_, _05469_, \oc8051_golden_model_1.ACC [5]);
  nor (_16879_, _05469_, \oc8051_golden_model_1.ACC [5]);
  or (_16880_, _16542_, _16879_);
  and (_16881_, _16880_, _16878_);
  nor (_16882_, _16881_, _08664_);
  and (_16883_, _16881_, _08664_);
  nor (_16884_, _16883_, _16882_);
  nor (_16885_, _16552_, _16547_);
  and (_16887_, _16885_, \oc8051_golden_model_1.PSW [7]);
  or (_16888_, _16887_, _16884_);
  nand (_16889_, _16887_, _16884_);
  and (_16890_, _16889_, _16888_);
  and (_16891_, _16890_, _10201_);
  or (_16892_, _16891_, _11350_);
  and (_16893_, _16892_, _16877_);
  or (_16894_, _16893_, _03761_);
  or (_16895_, _16894_, _16813_);
  and (_16896_, _16895_, _16799_);
  or (_16898_, _16464_, _10046_);
  and (_16899_, _16898_, _10045_);
  nor (_16900_, _16899_, _08738_);
  and (_16901_, _16899_, _08738_);
  nor (_16902_, _16901_, _16900_);
  nor (_16903_, _16474_, _16469_);
  and (_16904_, _16903_, \oc8051_golden_model_1.PSW [7]);
  or (_16905_, _16904_, _16902_);
  nand (_16906_, _16904_, _16902_);
  and (_16907_, _16906_, _16905_);
  and (_16909_, _16907_, _07913_);
  or (_16910_, _16909_, _07912_);
  or (_16911_, _16910_, _16896_);
  nand (_16912_, _03549_, _07912_);
  and (_16913_, _16912_, _03710_);
  and (_16914_, _16913_, _16911_);
  nor (_16915_, _13226_, _08339_);
  nor (_16916_, _16915_, _16839_);
  nor (_16917_, _16916_, _03710_);
  or (_16918_, _16917_, _07390_);
  or (_16920_, _16918_, _16914_);
  and (_16921_, _16920_, _16794_);
  or (_16922_, _16921_, _04481_);
  and (_16923_, _06455_, _05254_);
  nor (_16924_, _16923_, _16778_);
  nand (_16925_, _16924_, _04481_);
  and (_16926_, _16925_, _03589_);
  and (_16927_, _16926_, _16922_);
  nor (_16928_, _13332_, _07908_);
  nor (_16929_, _16928_, _16778_);
  nor (_16931_, _16929_, _03589_);
  or (_16932_, _16931_, _07405_);
  or (_16933_, _16932_, _16927_);
  not (_16934_, _07434_);
  and (_16935_, _07437_, _16934_);
  or (_16936_, _16935_, _07411_);
  and (_16937_, _16936_, _16933_);
  or (_16938_, _16937_, _03216_);
  and (_16939_, _16938_, _16791_);
  or (_16940_, _16939_, _03601_);
  nand (_16942_, _16780_, _03601_);
  and (_16943_, _16942_, _08364_);
  and (_16944_, _16943_, _16940_);
  nor (_16945_, _08364_, _03549_);
  or (_16946_, _16945_, _08371_);
  or (_16947_, _16946_, _16944_);
  and (_16948_, _16947_, _16790_);
  or (_16949_, _16948_, _08380_);
  or (_16950_, _08664_, _04180_);
  and (_16951_, _16950_, _16786_);
  and (_16953_, _16951_, _16949_);
  or (_16954_, _16953_, _16789_);
  and (_16955_, _16954_, _08393_);
  and (_16956_, _08392_, _08627_);
  or (_16957_, _16956_, _03778_);
  or (_16958_, _16957_, _16955_);
  or (_16959_, _13353_, _03779_);
  and (_16960_, _16959_, _07905_);
  and (_16961_, _16960_, _16958_);
  nor (_16962_, _08737_, _07905_);
  or (_16964_, _16962_, _03600_);
  or (_16965_, _16964_, _16961_);
  nand (_16966_, _16965_, _16785_);
  and (_16967_, _16966_, _07778_);
  nor (_16968_, _16778_, _07778_);
  or (_16969_, _16968_, _15103_);
  nor (_16970_, _16969_, _16967_);
  or (_16971_, _08662_, _04199_);
  and (_16972_, _16971_, _08421_);
  or (_16973_, _16972_, _16970_);
  or (_16975_, _08662_, _15367_);
  and (_16976_, _16975_, _16973_);
  or (_16977_, _16976_, _08420_);
  or (_16978_, _08425_, _08625_);
  and (_16979_, _16978_, _03789_);
  and (_16980_, _16979_, _16977_);
  or (_16981_, _13351_, _08429_);
  and (_16982_, _16981_, _08431_);
  or (_16983_, _16982_, _16980_);
  or (_16984_, _08435_, _08735_);
  and (_16986_, _16984_, _07777_);
  and (_16987_, _16986_, _16983_);
  or (_16988_, _16987_, _16782_);
  and (_16989_, _16988_, _08447_);
  nor (_16990_, _08447_, _08663_);
  or (_16991_, _16990_, _08450_);
  or (_16992_, _16991_, _16989_);
  nand (_16993_, _08450_, _08626_);
  and (_16994_, _16993_, _03784_);
  and (_16995_, _16994_, _16992_);
  nor (_16997_, _13352_, _03784_);
  or (_16998_, _16997_, _08458_);
  or (_16999_, _16998_, _16995_);
  nand (_17000_, _08458_, _08736_);
  and (_17001_, _17000_, _16999_);
  or (_17002_, _17001_, _03624_);
  nor (_17003_, _13346_, _07908_);
  nor (_17004_, _17003_, _16778_);
  nand (_17005_, _17004_, _03624_);
  and (_17006_, _17005_, _07898_);
  and (_17008_, _17006_, _17002_);
  and (_17009_, _07885_, _07832_);
  nor (_17010_, _17009_, _07886_);
  or (_17011_, _17010_, _08475_);
  and (_17012_, _17011_, _11885_);
  or (_17013_, _17012_, _17008_);
  and (_17014_, _08497_, _08479_);
  nor (_17015_, _17014_, _08498_);
  or (_17016_, _17015_, _08477_);
  and (_17017_, _17016_, _17013_);
  or (_17019_, _17017_, _03776_);
  and (_17020_, _08578_, _08531_);
  nor (_17021_, _17020_, _08579_);
  or (_17022_, _17021_, _03777_);
  and (_17023_, _17022_, _08589_);
  and (_17024_, _17023_, _17019_);
  and (_17025_, _08608_, _08591_);
  nor (_17026_, _17025_, _08609_);
  and (_17027_, _17026_, _08506_);
  or (_17028_, _17027_, _08587_);
  or (_17030_, _17028_, _17024_);
  nand (_17031_, _08587_, _07478_);
  and (_17032_, _17031_, _08617_);
  and (_17033_, _17032_, _17030_);
  nor (_17034_, _08691_, _08664_);
  nor (_17035_, _17034_, _08692_);
  and (_17036_, _17035_, _08618_);
  or (_17037_, _17036_, _17033_);
  and (_17038_, _17037_, _08624_);
  nor (_17039_, _08655_, _08627_);
  nor (_17041_, _17039_, _08656_);
  and (_17042_, _17041_, _08620_);
  or (_17043_, _17042_, _03517_);
  or (_17044_, _17043_, _17038_);
  and (_17045_, _08723_, _08206_);
  nor (_17046_, _17045_, _08724_);
  or (_17047_, _17046_, _03518_);
  and (_17048_, _17047_, _08734_);
  and (_17049_, _17048_, _17044_);
  nor (_17050_, _08763_, _08738_);
  nor (_17052_, _17050_, _08764_);
  and (_17053_, _17052_, _08701_);
  or (_17054_, _17053_, _08732_);
  or (_17055_, _17054_, _17049_);
  and (_17056_, _17055_, _16777_);
  or (_17057_, _17056_, _03815_);
  nand (_17058_, _16816_, _03815_);
  and (_17059_, _17058_, _08776_);
  and (_17060_, _17059_, _17057_);
  nor (_17061_, _08783_, _07433_);
  or (_17063_, _17061_, _08784_);
  and (_17064_, _17063_, _08775_);
  or (_17065_, _17064_, _08780_);
  or (_17066_, _17065_, _17060_);
  nand (_17067_, _08780_, _06075_);
  and (_17068_, _17067_, _03823_);
  and (_17069_, _17068_, _17066_);
  nor (_17070_, _16862_, _03823_);
  or (_17071_, _17070_, _03447_);
  or (_17072_, _17071_, _17069_);
  and (_17074_, _13402_, _05254_);
  nor (_17075_, _17074_, _16778_);
  nand (_17076_, _17075_, _03447_);
  and (_17077_, _17076_, _08799_);
  and (_17078_, _17077_, _17072_);
  nor (_17079_, _08809_, \oc8051_golden_model_1.ACC [6]);
  nor (_17080_, _17079_, _08810_);
  nor (_17081_, _17080_, _08805_);
  nor (_17082_, _17081_, _11964_);
  or (_17083_, _17082_, _17078_);
  nand (_17085_, _08805_, _06075_);
  and (_17086_, _17085_, _43000_);
  and (_17087_, _17086_, _17083_);
  or (_17088_, _17087_, _16775_);
  and (_43497_, _17088_, _41806_);
  not (_17089_, \oc8051_golden_model_1.DPL [0]);
  nor (_17090_, _43000_, _17089_);
  nor (_17091_, _05303_, _17089_);
  and (_17092_, _05303_, _04620_);
  or (_17093_, _17092_, _17091_);
  or (_17095_, _17093_, _06838_);
  and (_17096_, _05303_, \oc8051_golden_model_1.ACC [0]);
  or (_17097_, _17096_, _17091_);
  or (_17098_, _17097_, _03737_);
  nor (_17099_, _05666_, _08824_);
  or (_17100_, _17099_, _17091_);
  or (_17101_, _17100_, _04081_);
  and (_17102_, _17097_, _04409_);
  nor (_17103_, _04409_, _17089_);
  or (_17104_, _17103_, _03610_);
  or (_17106_, _17104_, _17102_);
  and (_17107_, _17106_, _03996_);
  and (_17108_, _17107_, _17101_);
  and (_17109_, _17093_, _03723_);
  or (_17110_, _17109_, _03729_);
  or (_17111_, _17110_, _17108_);
  and (_17112_, _17111_, _17098_);
  or (_17113_, _17112_, _08847_);
  nand (_17114_, _08847_, \oc8051_golden_model_1.DPL [0]);
  and (_17115_, _17114_, _08832_);
  and (_17117_, _17115_, _17113_);
  nor (_17118_, _04163_, _08832_);
  or (_17119_, _17118_, _07390_);
  or (_17120_, _17119_, _17117_);
  and (_17121_, _17120_, _17095_);
  or (_17122_, _17121_, _04481_);
  and (_17123_, _06546_, _05303_);
  or (_17124_, _17091_, _07400_);
  or (_17125_, _17124_, _17123_);
  and (_17126_, _17125_, _17122_);
  or (_17128_, _17126_, _03222_);
  nor (_17129_, _12109_, _08824_);
  or (_17130_, _17129_, _17091_);
  or (_17131_, _17130_, _03589_);
  and (_17132_, _17131_, _05886_);
  and (_17133_, _17132_, _17128_);
  and (_17134_, _05303_, _06274_);
  or (_17135_, _17134_, _17091_);
  and (_17136_, _17135_, _03601_);
  or (_17137_, _17136_, _03600_);
  or (_17139_, _17137_, _17133_);
  and (_17140_, _12124_, _05303_);
  or (_17141_, _17140_, _17091_);
  or (_17142_, _17141_, _07766_);
  and (_17143_, _17142_, _17139_);
  or (_17144_, _17143_, _03780_);
  and (_17145_, _12128_, _05303_);
  or (_17146_, _17145_, _17091_);
  or (_17147_, _17146_, _07778_);
  and (_17148_, _17147_, _07777_);
  and (_17150_, _17148_, _17144_);
  nand (_17151_, _17135_, _03622_);
  nor (_17152_, _17151_, _17099_);
  or (_17153_, _17152_, _17150_);
  and (_17154_, _17153_, _06828_);
  or (_17155_, _17091_, _05666_);
  and (_17156_, _17097_, _03790_);
  and (_17157_, _17156_, _17155_);
  or (_17158_, _17157_, _03624_);
  or (_17159_, _17158_, _17154_);
  nor (_17161_, _12122_, _08824_);
  or (_17162_, _17091_, _07795_);
  or (_17163_, _17162_, _17161_);
  and (_17164_, _17163_, _07793_);
  and (_17165_, _17164_, _17159_);
  not (_17166_, _03909_);
  nor (_17167_, _12003_, _08824_);
  or (_17168_, _17167_, _17091_);
  and (_17169_, _17168_, _03785_);
  or (_17170_, _17169_, _17166_);
  or (_17172_, _17170_, _17165_);
  or (_17173_, _17100_, _03909_);
  and (_17174_, _17173_, _43000_);
  and (_17175_, _17174_, _17172_);
  or (_17176_, _17175_, _17090_);
  and (_43498_, _17176_, _41806_);
  not (_17177_, \oc8051_golden_model_1.DPL [1]);
  nor (_17178_, _43000_, _17177_);
  nor (_17179_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_17180_, _17179_, _08852_);
  and (_17182_, _17180_, _08847_);
  or (_17183_, _05303_, \oc8051_golden_model_1.DPL [1]);
  and (_17184_, _12213_, _05303_);
  not (_17185_, _17184_);
  and (_17186_, _17185_, _17183_);
  or (_17187_, _17186_, _04081_);
  nand (_17188_, _05303_, _03274_);
  and (_17189_, _17188_, _17183_);
  and (_17190_, _17189_, _04409_);
  nor (_17191_, _04409_, _17177_);
  or (_17193_, _17191_, _03610_);
  or (_17194_, _17193_, _17190_);
  and (_17195_, _17194_, _03996_);
  and (_17196_, _17195_, _17187_);
  nor (_17197_, _05303_, _17177_);
  and (_17198_, _05303_, _06764_);
  or (_17199_, _17198_, _17197_);
  and (_17200_, _17199_, _03723_);
  or (_17201_, _17200_, _03729_);
  or (_17202_, _17201_, _17196_);
  or (_17204_, _17189_, _03737_);
  and (_17205_, _17204_, _08848_);
  and (_17206_, _17205_, _17202_);
  or (_17207_, _17206_, _17182_);
  and (_17208_, _17207_, _08832_);
  nor (_17209_, _04303_, _08832_);
  or (_17210_, _17209_, _07390_);
  or (_17211_, _17210_, _17208_);
  or (_17212_, _17199_, _06838_);
  and (_17213_, _17212_, _17211_);
  or (_17215_, _17213_, _04481_);
  and (_17216_, _06501_, _05303_);
  or (_17217_, _17197_, _07400_);
  or (_17218_, _17217_, _17216_);
  and (_17219_, _17218_, _03589_);
  and (_17220_, _17219_, _17215_);
  nor (_17221_, _12313_, _08824_);
  or (_17222_, _17221_, _17197_);
  and (_17223_, _17222_, _03222_);
  or (_17224_, _17223_, _17220_);
  and (_17226_, _17224_, _03602_);
  nand (_17227_, _05303_, _04303_);
  and (_17228_, _17183_, _03601_);
  and (_17229_, _17228_, _17227_);
  or (_17230_, _12327_, _08824_);
  and (_17231_, _17183_, _03600_);
  and (_17232_, _17231_, _17230_);
  or (_17233_, _17232_, _17229_);
  or (_17234_, _17233_, _17226_);
  and (_17235_, _17234_, _07778_);
  or (_17237_, _12333_, _08824_);
  and (_17238_, _17183_, _03780_);
  and (_17239_, _17238_, _17237_);
  or (_17240_, _17239_, _17235_);
  and (_17241_, _17240_, _07777_);
  or (_17242_, _12207_, _08824_);
  and (_17243_, _17183_, _03622_);
  and (_17244_, _17243_, _17242_);
  or (_17245_, _17244_, _17241_);
  and (_17246_, _17245_, _06828_);
  or (_17248_, _17197_, _05618_);
  and (_17249_, _17189_, _03790_);
  and (_17250_, _17249_, _17248_);
  or (_17251_, _17250_, _17246_);
  and (_17252_, _17251_, _03786_);
  or (_17253_, _17227_, _05618_);
  and (_17254_, _17183_, _03624_);
  and (_17255_, _17254_, _17253_);
  or (_17256_, _17188_, _05618_);
  and (_17257_, _17183_, _03785_);
  and (_17259_, _17257_, _17256_);
  or (_17260_, _17259_, _03815_);
  or (_17261_, _17260_, _17255_);
  or (_17262_, _17261_, _17252_);
  or (_17263_, _17186_, _04246_);
  and (_17264_, _17263_, _17262_);
  or (_17265_, _17264_, _03447_);
  or (_17266_, _17197_, _03514_);
  or (_17267_, _17266_, _17184_);
  and (_17268_, _17267_, _43000_);
  and (_17269_, _17268_, _17265_);
  or (_17270_, _17269_, _17178_);
  and (_43499_, _17270_, _41806_);
  not (_17271_, \oc8051_golden_model_1.DPL [2]);
  nor (_17272_, _43000_, _17271_);
  nor (_17273_, _05303_, _17271_);
  nor (_17274_, _12538_, _08824_);
  or (_17275_, _17274_, _17273_);
  and (_17276_, _17275_, _03785_);
  and (_17277_, _12539_, _05303_);
  or (_17280_, _17277_, _17273_);
  and (_17281_, _17280_, _03780_);
  nor (_17282_, _08824_, _04875_);
  or (_17283_, _17282_, _17273_);
  or (_17284_, _17283_, _03996_);
  nor (_17285_, _12416_, _08824_);
  or (_17286_, _17285_, _17273_);
  and (_17287_, _17286_, _03610_);
  nor (_17288_, _04409_, _17271_);
  and (_17289_, _05303_, \oc8051_golden_model_1.ACC [2]);
  or (_17290_, _17289_, _17273_);
  and (_17291_, _17290_, _04409_);
  or (_17292_, _17291_, _17288_);
  and (_17293_, _17292_, _04081_);
  or (_17294_, _17293_, _03723_);
  or (_17295_, _17294_, _17287_);
  and (_17296_, _17295_, _17284_);
  or (_17297_, _17296_, _03729_);
  or (_17298_, _17290_, _03737_);
  and (_17299_, _17298_, _08848_);
  and (_17302_, _17299_, _17297_);
  nor (_17303_, _08852_, \oc8051_golden_model_1.DPL [2]);
  nor (_17304_, _17303_, _08853_);
  and (_17305_, _17304_, _08847_);
  or (_17306_, _17305_, _17302_);
  and (_17307_, _17306_, _08832_);
  nor (_17308_, _03946_, _08832_);
  or (_17309_, _17308_, _07390_);
  or (_17310_, _17309_, _17307_);
  or (_17311_, _17283_, _06838_);
  and (_17313_, _17311_, _17310_);
  or (_17314_, _17313_, _04481_);
  and (_17315_, _06637_, _05303_);
  or (_17316_, _17273_, _07400_);
  or (_17317_, _17316_, _17315_);
  and (_17318_, _17317_, _03589_);
  and (_17319_, _17318_, _17314_);
  nor (_17320_, _12519_, _08824_);
  or (_17321_, _17320_, _17273_);
  and (_17322_, _17321_, _03222_);
  or (_17324_, _17322_, _08828_);
  or (_17325_, _17324_, _17319_);
  and (_17326_, _12533_, _05303_);
  or (_17327_, _17273_, _07766_);
  or (_17328_, _17327_, _17326_);
  and (_17329_, _05303_, _06332_);
  or (_17330_, _17329_, _17273_);
  or (_17331_, _17330_, _05886_);
  and (_17332_, _17331_, _07778_);
  and (_17333_, _17332_, _17328_);
  and (_17335_, _17333_, _17325_);
  or (_17336_, _17335_, _17281_);
  and (_17337_, _17336_, _07777_);
  or (_17338_, _17273_, _05718_);
  and (_17339_, _17330_, _03622_);
  and (_17340_, _17339_, _17338_);
  or (_17341_, _17340_, _17337_);
  and (_17342_, _17341_, _06828_);
  and (_17343_, _17290_, _03790_);
  and (_17344_, _17343_, _17338_);
  or (_17346_, _17344_, _03624_);
  or (_17347_, _17346_, _17342_);
  nor (_17348_, _12532_, _08824_);
  or (_17349_, _17273_, _07795_);
  or (_17350_, _17349_, _17348_);
  and (_17351_, _17350_, _07793_);
  and (_17352_, _17351_, _17347_);
  or (_17353_, _17352_, _17276_);
  and (_17354_, _17353_, _04246_);
  and (_17355_, _17286_, _03815_);
  or (_17357_, _17355_, _03447_);
  or (_17358_, _17357_, _17354_);
  and (_17359_, _12592_, _05303_);
  or (_17360_, _17273_, _03514_);
  or (_17361_, _17360_, _17359_);
  and (_17362_, _17361_, _43000_);
  and (_17363_, _17362_, _17358_);
  or (_17364_, _17363_, _17272_);
  and (_43500_, _17364_, _41806_);
  not (_17365_, \oc8051_golden_model_1.DPL [3]);
  nor (_17367_, _43000_, _17365_);
  nor (_17368_, _05303_, _17365_);
  nor (_17369_, _12738_, _08824_);
  or (_17370_, _17369_, _17368_);
  and (_17371_, _17370_, _03785_);
  and (_17372_, _12739_, _05303_);
  or (_17373_, _17372_, _17368_);
  and (_17374_, _17373_, _03780_);
  nor (_17375_, _08853_, \oc8051_golden_model_1.DPL [3]);
  nor (_17376_, _17375_, _08854_);
  and (_17378_, _17376_, _08847_);
  nor (_17379_, _12627_, _08824_);
  or (_17380_, _17379_, _17368_);
  or (_17381_, _17380_, _04081_);
  and (_17382_, _05303_, \oc8051_golden_model_1.ACC [3]);
  or (_17383_, _17382_, _17368_);
  and (_17384_, _17383_, _04409_);
  nor (_17385_, _04409_, _17365_);
  or (_17386_, _17385_, _03610_);
  or (_17387_, _17386_, _17384_);
  and (_17389_, _17387_, _03996_);
  and (_17390_, _17389_, _17381_);
  nor (_17391_, _08824_, _05005_);
  or (_17392_, _17391_, _17368_);
  and (_17393_, _17392_, _03723_);
  or (_17394_, _17393_, _03729_);
  or (_17395_, _17394_, _17390_);
  or (_17396_, _17383_, _03737_);
  and (_17397_, _17396_, _08848_);
  and (_17398_, _17397_, _17395_);
  or (_17400_, _17398_, _17378_);
  and (_17401_, _17400_, _08832_);
  nor (_17402_, _03708_, _08832_);
  or (_17403_, _17402_, _07390_);
  or (_17404_, _17403_, _17401_);
  or (_17405_, _17392_, _06838_);
  and (_17406_, _17405_, _17404_);
  or (_17407_, _17406_, _04481_);
  and (_17408_, _06592_, _05303_);
  or (_17409_, _17368_, _07400_);
  or (_17411_, _17409_, _17408_);
  and (_17412_, _17411_, _03589_);
  and (_17413_, _17412_, _17407_);
  nor (_17414_, _12718_, _08824_);
  or (_17415_, _17414_, _17368_);
  and (_17416_, _17415_, _03222_);
  or (_17417_, _17416_, _08828_);
  or (_17418_, _17417_, _17413_);
  and (_17419_, _12733_, _05303_);
  or (_17420_, _17368_, _07766_);
  or (_17422_, _17420_, _17419_);
  and (_17423_, _05303_, _06276_);
  or (_17424_, _17423_, _17368_);
  or (_17425_, _17424_, _05886_);
  and (_17426_, _17425_, _07778_);
  and (_17427_, _17426_, _17422_);
  and (_17428_, _17427_, _17418_);
  or (_17429_, _17428_, _17374_);
  and (_17430_, _17429_, _07777_);
  or (_17431_, _17368_, _05567_);
  and (_17433_, _17424_, _03622_);
  and (_17434_, _17433_, _17431_);
  or (_17435_, _17434_, _17430_);
  and (_17436_, _17435_, _06828_);
  and (_17437_, _17383_, _03790_);
  and (_17438_, _17437_, _17431_);
  or (_17439_, _17438_, _03624_);
  or (_17440_, _17439_, _17436_);
  nor (_17441_, _12732_, _08824_);
  or (_17442_, _17368_, _07795_);
  or (_17444_, _17442_, _17441_);
  and (_17445_, _17444_, _07793_);
  and (_17446_, _17445_, _17440_);
  or (_17447_, _17446_, _17371_);
  and (_17448_, _17447_, _04246_);
  and (_17449_, _17380_, _03815_);
  or (_17450_, _17449_, _03447_);
  or (_17451_, _17450_, _17448_);
  and (_17452_, _12794_, _05303_);
  or (_17453_, _17368_, _03514_);
  or (_17455_, _17453_, _17452_);
  and (_17456_, _17455_, _43000_);
  and (_17457_, _17456_, _17451_);
  or (_17458_, _17457_, _17367_);
  and (_43501_, _17458_, _41806_);
  not (_17459_, \oc8051_golden_model_1.DPL [4]);
  nor (_17460_, _43000_, _17459_);
  nor (_17461_, _05303_, _17459_);
  nor (_17462_, _12816_, _08824_);
  or (_17463_, _17462_, _17461_);
  and (_17465_, _17463_, _03785_);
  nor (_17466_, _05777_, _08824_);
  or (_17467_, _17466_, _17461_);
  or (_17468_, _17467_, _06838_);
  nor (_17469_, _12841_, _08824_);
  or (_17470_, _17469_, _17461_);
  or (_17471_, _17470_, _04081_);
  and (_17472_, _05303_, \oc8051_golden_model_1.ACC [4]);
  or (_17473_, _17472_, _17461_);
  and (_17474_, _17473_, _04409_);
  nor (_17476_, _04409_, _17459_);
  or (_17477_, _17476_, _03610_);
  or (_17478_, _17477_, _17474_);
  and (_17479_, _17478_, _03996_);
  and (_17480_, _17479_, _17471_);
  and (_17481_, _17467_, _03723_);
  or (_17482_, _17481_, _03729_);
  or (_17483_, _17482_, _17480_);
  or (_17484_, _17473_, _03737_);
  and (_17485_, _17484_, _08848_);
  and (_17487_, _17485_, _17483_);
  nor (_17488_, _08854_, \oc8051_golden_model_1.DPL [4]);
  nor (_17489_, _17488_, _08855_);
  and (_17490_, _17489_, _08847_);
  or (_17491_, _17490_, _17487_);
  and (_17492_, _17491_, _08832_);
  nor (_17493_, _06236_, _08832_);
  or (_17494_, _17493_, _07390_);
  or (_17495_, _17494_, _17492_);
  and (_17496_, _17495_, _17468_);
  or (_17498_, _17496_, _04481_);
  and (_17499_, _06730_, _05303_);
  or (_17500_, _17461_, _07400_);
  or (_17501_, _17500_, _17499_);
  and (_17502_, _17501_, _03589_);
  and (_17503_, _17502_, _17498_);
  nor (_17504_, _12933_, _08824_);
  or (_17505_, _17504_, _17461_);
  and (_17506_, _17505_, _03222_);
  or (_17507_, _17506_, _17503_);
  or (_17509_, _17507_, _08828_);
  and (_17510_, _12821_, _05303_);
  or (_17511_, _17461_, _07766_);
  or (_17512_, _17511_, _17510_);
  and (_17513_, _06298_, _05303_);
  or (_17514_, _17513_, _17461_);
  or (_17515_, _17514_, _05886_);
  and (_17516_, _17515_, _07778_);
  and (_17517_, _17516_, _17512_);
  and (_17518_, _17517_, _17509_);
  and (_17520_, _12817_, _05303_);
  or (_17521_, _17520_, _17461_);
  and (_17522_, _17521_, _03780_);
  or (_17523_, _17522_, _17518_);
  and (_17524_, _17523_, _07777_);
  or (_17525_, _17461_, _05825_);
  and (_17526_, _17514_, _03622_);
  and (_17527_, _17526_, _17525_);
  or (_17528_, _17527_, _17524_);
  and (_17529_, _17528_, _06828_);
  and (_17531_, _17473_, _03790_);
  and (_17532_, _17531_, _17525_);
  or (_17533_, _17532_, _03624_);
  or (_17534_, _17533_, _17529_);
  nor (_17535_, _12819_, _08824_);
  or (_17536_, _17461_, _07795_);
  or (_17537_, _17536_, _17535_);
  and (_17538_, _17537_, _07793_);
  and (_17539_, _17538_, _17534_);
  or (_17540_, _17539_, _17465_);
  and (_17542_, _17540_, _04246_);
  and (_17543_, _17470_, _03815_);
  or (_17544_, _17543_, _03447_);
  or (_17545_, _17544_, _17542_);
  and (_17546_, _13003_, _05303_);
  or (_17547_, _17461_, _03514_);
  or (_17548_, _17547_, _17546_);
  and (_17549_, _17548_, _43000_);
  and (_17550_, _17549_, _17545_);
  or (_17551_, _17550_, _17460_);
  and (_43502_, _17551_, _41806_);
  not (_17553_, \oc8051_golden_model_1.DPL [5]);
  nor (_17554_, _43000_, _17553_);
  nor (_17555_, _05303_, _17553_);
  nor (_17556_, _13146_, _08824_);
  or (_17557_, _17556_, _17555_);
  and (_17558_, _17557_, _03785_);
  nor (_17559_, _05469_, _08824_);
  or (_17560_, _17559_, _17555_);
  or (_17561_, _17560_, _06838_);
  nor (_17563_, _13014_, _08824_);
  or (_17564_, _17563_, _17555_);
  or (_17565_, _17564_, _04081_);
  and (_17566_, _05303_, \oc8051_golden_model_1.ACC [5]);
  or (_17567_, _17566_, _17555_);
  and (_17568_, _17567_, _04409_);
  nor (_17569_, _04409_, _17553_);
  or (_17570_, _17569_, _03610_);
  or (_17571_, _17570_, _17568_);
  and (_17572_, _17571_, _03996_);
  and (_17574_, _17572_, _17565_);
  and (_17575_, _17560_, _03723_);
  or (_17576_, _17575_, _03729_);
  or (_17577_, _17576_, _17574_);
  or (_17578_, _17567_, _03737_);
  and (_17579_, _17578_, _08848_);
  and (_17580_, _17579_, _17577_);
  nor (_17581_, _08855_, \oc8051_golden_model_1.DPL [5]);
  nor (_17582_, _17581_, _08856_);
  and (_17583_, _17582_, _08847_);
  or (_17585_, _17583_, _17580_);
  and (_17586_, _17585_, _08832_);
  nor (_17587_, _06267_, _08832_);
  or (_17588_, _17587_, _07390_);
  or (_17589_, _17588_, _17586_);
  and (_17590_, _17589_, _17561_);
  or (_17591_, _17590_, _04481_);
  and (_17592_, _06684_, _05303_);
  or (_17593_, _17555_, _07400_);
  or (_17594_, _17593_, _17592_);
  and (_17596_, _17594_, _03589_);
  and (_17597_, _17596_, _17591_);
  nor (_17598_, _13127_, _08824_);
  or (_17599_, _17598_, _17555_);
  and (_17600_, _17599_, _03222_);
  or (_17601_, _17600_, _17597_);
  or (_17602_, _17601_, _08828_);
  and (_17603_, _13141_, _05303_);
  or (_17604_, _17555_, _07766_);
  or (_17605_, _17604_, _17603_);
  and (_17607_, _06306_, _05303_);
  or (_17608_, _17607_, _17555_);
  or (_17609_, _17608_, _05886_);
  and (_17610_, _17609_, _07778_);
  and (_17611_, _17610_, _17605_);
  and (_17612_, _17611_, _17602_);
  and (_17613_, _13147_, _05303_);
  or (_17614_, _17613_, _17555_);
  and (_17615_, _17614_, _03780_);
  or (_17616_, _17615_, _17612_);
  and (_17618_, _17616_, _07777_);
  or (_17619_, _17555_, _05518_);
  and (_17620_, _17608_, _03622_);
  and (_17621_, _17620_, _17619_);
  or (_17622_, _17621_, _17618_);
  and (_17623_, _17622_, _06828_);
  and (_17624_, _17567_, _03790_);
  and (_17625_, _17624_, _17619_);
  or (_17626_, _17625_, _03624_);
  or (_17627_, _17626_, _17623_);
  nor (_17629_, _13140_, _08824_);
  or (_17630_, _17555_, _07795_);
  or (_17631_, _17630_, _17629_);
  and (_17632_, _17631_, _07793_);
  and (_17633_, _17632_, _17627_);
  or (_17634_, _17633_, _17558_);
  and (_17635_, _17634_, _04246_);
  and (_17636_, _17564_, _03815_);
  or (_17637_, _17636_, _03447_);
  or (_17638_, _17637_, _17635_);
  and (_17640_, _13199_, _05303_);
  or (_17641_, _17555_, _03514_);
  or (_17642_, _17641_, _17640_);
  and (_17643_, _17642_, _43000_);
  and (_17644_, _17643_, _17638_);
  or (_17645_, _17644_, _17554_);
  and (_43505_, _17645_, _41806_);
  not (_17646_, \oc8051_golden_model_1.DPL [6]);
  nor (_17647_, _43000_, _17646_);
  nor (_17648_, _05303_, _17646_);
  nor (_17650_, _13352_, _08824_);
  or (_17651_, _17650_, _17648_);
  and (_17652_, _17651_, _03785_);
  nor (_17653_, _05363_, _08824_);
  or (_17654_, _17653_, _17648_);
  or (_17655_, _17654_, _06838_);
  nor (_17656_, _13242_, _08824_);
  or (_17657_, _17656_, _17648_);
  or (_17658_, _17657_, _04081_);
  and (_17659_, _05303_, \oc8051_golden_model_1.ACC [6]);
  or (_17661_, _17659_, _17648_);
  and (_17662_, _17661_, _04409_);
  nor (_17663_, _04409_, _17646_);
  or (_17664_, _17663_, _03610_);
  or (_17665_, _17664_, _17662_);
  and (_17666_, _17665_, _03996_);
  and (_17667_, _17666_, _17658_);
  and (_17668_, _17654_, _03723_);
  or (_17669_, _17668_, _03729_);
  or (_17670_, _17669_, _17667_);
  or (_17672_, _17661_, _03737_);
  and (_17673_, _17672_, _08848_);
  and (_17674_, _17673_, _17670_);
  nor (_17675_, _08856_, \oc8051_golden_model_1.DPL [6]);
  nor (_17676_, _17675_, _08857_);
  and (_17677_, _17676_, _08847_);
  or (_17678_, _17677_, _17674_);
  and (_17679_, _17678_, _08832_);
  nor (_17680_, _06204_, _08832_);
  or (_17681_, _17680_, _07390_);
  or (_17683_, _17681_, _17679_);
  and (_17684_, _17683_, _17655_);
  or (_17685_, _17684_, _04481_);
  and (_17686_, _06455_, _05303_);
  or (_17687_, _17648_, _07400_);
  or (_17688_, _17687_, _17686_);
  and (_17689_, _17688_, _03589_);
  and (_17690_, _17689_, _17685_);
  nor (_17691_, _13332_, _08824_);
  or (_17692_, _17691_, _17648_);
  and (_17694_, _17692_, _03222_);
  or (_17695_, _17694_, _17690_);
  or (_17696_, _17695_, _08828_);
  and (_17697_, _13347_, _05303_);
  or (_17698_, _17648_, _07766_);
  or (_17699_, _17698_, _17697_);
  and (_17700_, _13339_, _05303_);
  or (_17701_, _17700_, _17648_);
  or (_17702_, _17701_, _05886_);
  and (_17703_, _17702_, _07778_);
  and (_17705_, _17703_, _17699_);
  and (_17706_, _17705_, _17696_);
  and (_17707_, _13353_, _05303_);
  or (_17708_, _17707_, _17648_);
  and (_17709_, _17708_, _03780_);
  or (_17710_, _17709_, _17706_);
  and (_17711_, _17710_, _07777_);
  or (_17712_, _17648_, _05412_);
  and (_17713_, _17701_, _03622_);
  and (_17714_, _17713_, _17712_);
  or (_17716_, _17714_, _17711_);
  and (_17717_, _17716_, _06828_);
  and (_17718_, _17661_, _03790_);
  and (_17719_, _17718_, _17712_);
  or (_17720_, _17719_, _03624_);
  or (_17721_, _17720_, _17717_);
  nor (_17722_, _13346_, _08824_);
  or (_17723_, _17648_, _07795_);
  or (_17724_, _17723_, _17722_);
  and (_17725_, _17724_, _07793_);
  and (_17727_, _17725_, _17721_);
  or (_17728_, _17727_, _17652_);
  and (_17729_, _17728_, _04246_);
  and (_17730_, _17657_, _03815_);
  or (_17731_, _17730_, _03447_);
  or (_17732_, _17731_, _17729_);
  and (_17733_, _13402_, _05303_);
  or (_17734_, _17648_, _03514_);
  or (_17735_, _17734_, _17733_);
  and (_17736_, _17735_, _43000_);
  and (_17738_, _17736_, _17732_);
  or (_17739_, _17738_, _17647_);
  and (_43506_, _17739_, _41806_);
  not (_17740_, \oc8051_golden_model_1.DPH [0]);
  nor (_17741_, _43000_, _17740_);
  nor (_17742_, _08859_, \oc8051_golden_model_1.DPH [0]);
  nor (_17743_, _17742_, _08947_);
  and (_17744_, _17743_, _08847_);
  nor (_17745_, _05297_, _17740_);
  nor (_17746_, _05666_, _08921_);
  or (_17748_, _17746_, _17745_);
  or (_17749_, _17748_, _04081_);
  and (_17750_, _05297_, \oc8051_golden_model_1.ACC [0]);
  or (_17751_, _17750_, _17745_);
  and (_17752_, _17751_, _04409_);
  nor (_17753_, _04409_, _17740_);
  or (_17754_, _17753_, _03610_);
  or (_17755_, _17754_, _17752_);
  and (_17756_, _17755_, _03996_);
  and (_17757_, _17756_, _17749_);
  and (_17759_, _05297_, _04620_);
  or (_17760_, _17759_, _17745_);
  and (_17761_, _17760_, _03723_);
  or (_17762_, _17761_, _03729_);
  or (_17763_, _17762_, _17757_);
  or (_17764_, _17751_, _03737_);
  and (_17765_, _17764_, _08848_);
  and (_17766_, _17765_, _17763_);
  or (_17767_, _17766_, _17744_);
  and (_17768_, _17767_, _08832_);
  nor (_17770_, _04048_, _08832_);
  or (_17771_, _17770_, _07390_);
  or (_17772_, _17771_, _17768_);
  or (_17773_, _17760_, _06838_);
  and (_17774_, _17773_, _17772_);
  or (_17775_, _17774_, _04481_);
  and (_17776_, _06546_, _05297_);
  or (_17777_, _17745_, _07400_);
  or (_17778_, _17777_, _17776_);
  and (_17779_, _17778_, _17775_);
  or (_17781_, _17779_, _03222_);
  nor (_17782_, _12109_, _08921_);
  or (_17783_, _17782_, _17745_);
  or (_17784_, _17783_, _03589_);
  and (_17785_, _17784_, _05886_);
  and (_17786_, _17785_, _17781_);
  and (_17787_, _05297_, _06274_);
  or (_17788_, _17787_, _17745_);
  and (_17789_, _17788_, _03601_);
  or (_17790_, _17789_, _03600_);
  or (_17792_, _17790_, _17786_);
  and (_17793_, _12124_, _05297_);
  or (_17794_, _17793_, _17745_);
  or (_17795_, _17794_, _07766_);
  and (_17796_, _17795_, _17792_);
  or (_17797_, _17796_, _03780_);
  and (_17798_, _12128_, _05297_);
  or (_17799_, _17798_, _17745_);
  or (_17800_, _17799_, _07778_);
  and (_17801_, _17800_, _07777_);
  and (_17803_, _17801_, _17797_);
  nand (_17804_, _17788_, _03622_);
  nor (_17805_, _17804_, _17746_);
  or (_17806_, _17805_, _17803_);
  and (_17807_, _17806_, _06828_);
  or (_17808_, _17745_, _05666_);
  and (_17809_, _17751_, _03790_);
  and (_17810_, _17809_, _17808_);
  or (_17811_, _17810_, _03624_);
  or (_17812_, _17811_, _17807_);
  nor (_17814_, _12122_, _08921_);
  or (_17815_, _17745_, _07795_);
  or (_17816_, _17815_, _17814_);
  and (_17817_, _17816_, _07793_);
  and (_17818_, _17817_, _17812_);
  nor (_17819_, _12003_, _08921_);
  or (_17820_, _17819_, _17745_);
  and (_17821_, _17820_, _03785_);
  or (_17822_, _17821_, _17166_);
  or (_17823_, _17822_, _17818_);
  or (_17825_, _17748_, _03909_);
  and (_17826_, _17825_, _43000_);
  and (_17827_, _17826_, _17823_);
  or (_17828_, _17827_, _17741_);
  and (_43507_, _17828_, _41806_);
  not (_17829_, \oc8051_golden_model_1.DPH [1]);
  nor (_17830_, _43000_, _17829_);
  nor (_17831_, _05297_, _17829_);
  and (_17832_, _05297_, _06764_);
  or (_17833_, _17832_, _17831_);
  or (_17835_, _17833_, _03996_);
  or (_17836_, _05297_, \oc8051_golden_model_1.DPH [1]);
  and (_17837_, _12213_, _05297_);
  not (_17838_, _17837_);
  and (_17839_, _17838_, _17836_);
  and (_17840_, _17839_, _03610_);
  nand (_17841_, _05297_, _03274_);
  and (_17842_, _17841_, _17836_);
  and (_17843_, _17842_, _04409_);
  nor (_17844_, _04409_, _17829_);
  or (_17846_, _17844_, _17843_);
  and (_17847_, _17846_, _04081_);
  or (_17848_, _17847_, _03723_);
  or (_17849_, _17848_, _17840_);
  and (_17850_, _17849_, _17835_);
  or (_17851_, _17850_, _03729_);
  or (_17852_, _17842_, _03737_);
  and (_17853_, _17852_, _08848_);
  and (_17854_, _17853_, _17851_);
  nor (_17855_, _08947_, \oc8051_golden_model_1.DPH [1]);
  nor (_17857_, _17855_, _08948_);
  and (_17858_, _17857_, _08847_);
  or (_17859_, _17858_, _17854_);
  and (_17860_, _17859_, _08832_);
  nor (_17861_, _03414_, _08832_);
  or (_17862_, _17861_, _07390_);
  or (_17863_, _17862_, _17860_);
  or (_17864_, _17833_, _06838_);
  and (_17865_, _17864_, _17863_);
  or (_17866_, _17865_, _04481_);
  and (_17868_, _06501_, _05297_);
  or (_17869_, _17831_, _07400_);
  or (_17870_, _17869_, _17868_);
  and (_17871_, _17870_, _03589_);
  and (_17872_, _17871_, _17866_);
  nand (_17873_, _12313_, _05297_);
  and (_17874_, _17836_, _03222_);
  and (_17875_, _17874_, _17873_);
  or (_17876_, _17875_, _17872_);
  and (_17877_, _17876_, _03602_);
  or (_17879_, _12327_, _08921_);
  and (_17880_, _17879_, _03600_);
  nand (_17881_, _05297_, _04303_);
  and (_17882_, _17881_, _03601_);
  or (_17883_, _17882_, _17880_);
  and (_17884_, _17883_, _17836_);
  or (_17885_, _17884_, _17877_);
  and (_17886_, _17885_, _07778_);
  or (_17887_, _12333_, _08921_);
  and (_17888_, _17836_, _03780_);
  and (_17890_, _17888_, _17887_);
  or (_17891_, _17890_, _17886_);
  and (_17892_, _17891_, _07777_);
  or (_17893_, _12207_, _08921_);
  and (_17894_, _17836_, _03622_);
  and (_17895_, _17894_, _17893_);
  or (_17896_, _17895_, _17892_);
  and (_17897_, _17896_, _06828_);
  or (_17898_, _17831_, _05618_);
  and (_17899_, _17842_, _03790_);
  and (_17901_, _17899_, _17898_);
  or (_17902_, _17901_, _17897_);
  and (_17903_, _17902_, _03786_);
  or (_17904_, _17881_, _05618_);
  and (_17905_, _17836_, _03624_);
  and (_17906_, _17905_, _17904_);
  or (_17907_, _17841_, _05618_);
  and (_17908_, _17836_, _03785_);
  and (_17909_, _17908_, _17907_);
  or (_17910_, _17909_, _03815_);
  or (_17912_, _17910_, _17906_);
  or (_17913_, _17912_, _17903_);
  or (_17914_, _17839_, _04246_);
  and (_17915_, _17914_, _17913_);
  or (_17916_, _17915_, _03447_);
  or (_17917_, _17831_, _03514_);
  or (_17918_, _17917_, _17837_);
  and (_17919_, _17918_, _43000_);
  and (_17920_, _17919_, _17916_);
  or (_17921_, _17920_, _17830_);
  and (_43510_, _17921_, _41806_);
  not (_17923_, \oc8051_golden_model_1.DPH [2]);
  nor (_17924_, _43000_, _17923_);
  nor (_17925_, _05297_, _17923_);
  nor (_17926_, _12538_, _08921_);
  or (_17927_, _17926_, _17925_);
  and (_17928_, _17927_, _03785_);
  and (_17929_, _12539_, _05297_);
  or (_17930_, _17929_, _17925_);
  and (_17931_, _17930_, _03780_);
  nor (_17933_, _08921_, _04875_);
  or (_17934_, _17933_, _17925_);
  or (_17935_, _17934_, _06838_);
  nor (_17936_, _12416_, _08921_);
  or (_17937_, _17936_, _17925_);
  or (_17938_, _17937_, _04081_);
  and (_17939_, _05297_, \oc8051_golden_model_1.ACC [2]);
  or (_17940_, _17939_, _17925_);
  and (_17941_, _17940_, _04409_);
  nor (_17942_, _04409_, _17923_);
  or (_17944_, _17942_, _03610_);
  or (_17945_, _17944_, _17941_);
  and (_17946_, _17945_, _03996_);
  and (_17947_, _17946_, _17938_);
  and (_17948_, _17934_, _03723_);
  or (_17949_, _17948_, _03729_);
  or (_17950_, _17949_, _17947_);
  or (_17951_, _17940_, _03737_);
  and (_17952_, _17951_, _08848_);
  and (_17953_, _17952_, _17950_);
  or (_17955_, _08948_, \oc8051_golden_model_1.DPH [2]);
  nor (_17956_, _08949_, _08848_);
  and (_17957_, _17956_, _17955_);
  or (_17958_, _17957_, _17953_);
  and (_17959_, _17958_, _08832_);
  nor (_17960_, _03904_, _08832_);
  or (_17961_, _17960_, _07390_);
  or (_17962_, _17961_, _17959_);
  and (_17963_, _17962_, _17935_);
  or (_17964_, _17963_, _04481_);
  and (_17966_, _06637_, _05297_);
  or (_17967_, _17925_, _07400_);
  or (_17968_, _17967_, _17966_);
  and (_17969_, _17968_, _03589_);
  and (_17970_, _17969_, _17964_);
  nor (_17971_, _12519_, _08921_);
  or (_17972_, _17971_, _17925_);
  and (_17973_, _17972_, _03222_);
  or (_17974_, _17973_, _17970_);
  or (_17975_, _17974_, _08828_);
  and (_17977_, _12533_, _05297_);
  or (_17978_, _17925_, _07766_);
  or (_17979_, _17978_, _17977_);
  and (_17980_, _05297_, _06332_);
  or (_17981_, _17980_, _17925_);
  or (_17982_, _17981_, _05886_);
  and (_17983_, _17982_, _07778_);
  and (_17984_, _17983_, _17979_);
  and (_17985_, _17984_, _17975_);
  or (_17986_, _17985_, _17931_);
  and (_17988_, _17986_, _07777_);
  or (_17989_, _17925_, _05718_);
  and (_17990_, _17981_, _03622_);
  and (_17991_, _17990_, _17989_);
  or (_17992_, _17991_, _17988_);
  and (_17993_, _17992_, _06828_);
  and (_17994_, _17940_, _03790_);
  and (_17995_, _17994_, _17989_);
  or (_17996_, _17995_, _03624_);
  or (_17997_, _17996_, _17993_);
  nor (_17999_, _12532_, _08921_);
  or (_18000_, _17925_, _07795_);
  or (_18001_, _18000_, _17999_);
  and (_18002_, _18001_, _07793_);
  and (_18003_, _18002_, _17997_);
  or (_18004_, _18003_, _17928_);
  and (_18005_, _18004_, _04246_);
  and (_18006_, _17937_, _03815_);
  or (_18007_, _18006_, _03447_);
  or (_18008_, _18007_, _18005_);
  and (_18010_, _12592_, _05297_);
  or (_18011_, _17925_, _03514_);
  or (_18012_, _18011_, _18010_);
  and (_18013_, _18012_, _43000_);
  and (_18014_, _18013_, _18008_);
  or (_18015_, _18014_, _17924_);
  and (_43511_, _18015_, _41806_);
  not (_18016_, \oc8051_golden_model_1.DPH [3]);
  nor (_18017_, _43000_, _18016_);
  nor (_18018_, _05297_, _18016_);
  nor (_18020_, _12738_, _08921_);
  or (_18021_, _18020_, _18018_);
  and (_18022_, _18021_, _03785_);
  and (_18023_, _12739_, _05297_);
  or (_18024_, _18023_, _18018_);
  and (_18025_, _18024_, _03780_);
  nor (_18026_, _12627_, _08921_);
  or (_18027_, _18026_, _18018_);
  or (_18028_, _18027_, _04081_);
  and (_18029_, _05297_, \oc8051_golden_model_1.ACC [3]);
  or (_18031_, _18029_, _18018_);
  and (_18032_, _18031_, _04409_);
  nor (_18033_, _04409_, _18016_);
  or (_18034_, _18033_, _03610_);
  or (_18035_, _18034_, _18032_);
  and (_18036_, _18035_, _03996_);
  and (_18037_, _18036_, _18028_);
  nor (_18038_, _08921_, _05005_);
  or (_18039_, _18038_, _18018_);
  and (_18040_, _18039_, _03723_);
  or (_18042_, _18040_, _03729_);
  or (_18043_, _18042_, _18037_);
  or (_18044_, _18031_, _03737_);
  and (_18045_, _18044_, _08848_);
  and (_18046_, _18045_, _18043_);
  or (_18047_, _08949_, \oc8051_golden_model_1.DPH [3]);
  nor (_18048_, _08950_, _08848_);
  and (_18049_, _18048_, _18047_);
  or (_18050_, _18049_, _18046_);
  and (_18051_, _18050_, _08832_);
  nor (_18053_, _08832_, _03581_);
  or (_18054_, _18053_, _07390_);
  or (_18055_, _18054_, _18051_);
  or (_18056_, _18039_, _06838_);
  and (_18057_, _18056_, _18055_);
  or (_18058_, _18057_, _04481_);
  and (_18059_, _06592_, _05297_);
  or (_18060_, _18018_, _07400_);
  or (_18061_, _18060_, _18059_);
  and (_18062_, _18061_, _03589_);
  and (_18064_, _18062_, _18058_);
  nor (_18065_, _12718_, _08921_);
  or (_18066_, _18065_, _18018_);
  and (_18067_, _18066_, _03222_);
  or (_18068_, _18067_, _08828_);
  or (_18069_, _18068_, _18064_);
  and (_18070_, _12733_, _05297_);
  or (_18071_, _18018_, _07766_);
  or (_18072_, _18071_, _18070_);
  and (_18073_, _05297_, _06276_);
  or (_18075_, _18073_, _18018_);
  or (_18076_, _18075_, _05886_);
  and (_18077_, _18076_, _07778_);
  and (_18078_, _18077_, _18072_);
  and (_18079_, _18078_, _18069_);
  or (_18080_, _18079_, _18025_);
  and (_18081_, _18080_, _07777_);
  or (_18082_, _18018_, _05567_);
  and (_18083_, _18075_, _03622_);
  and (_18084_, _18083_, _18082_);
  or (_18086_, _18084_, _18081_);
  and (_18087_, _18086_, _06828_);
  and (_18088_, _18031_, _03790_);
  and (_18089_, _18088_, _18082_);
  or (_18090_, _18089_, _03624_);
  or (_18091_, _18090_, _18087_);
  nor (_18092_, _12732_, _08921_);
  or (_18093_, _18018_, _07795_);
  or (_18094_, _18093_, _18092_);
  and (_18095_, _18094_, _07793_);
  and (_18097_, _18095_, _18091_);
  or (_18098_, _18097_, _18022_);
  and (_18099_, _18098_, _04246_);
  and (_18100_, _18027_, _03815_);
  or (_18101_, _18100_, _03447_);
  or (_18102_, _18101_, _18099_);
  and (_18103_, _12794_, _05297_);
  or (_18104_, _18018_, _03514_);
  or (_18105_, _18104_, _18103_);
  and (_18106_, _18105_, _43000_);
  and (_18108_, _18106_, _18102_);
  or (_18109_, _18108_, _18017_);
  and (_43512_, _18109_, _41806_);
  not (_18110_, \oc8051_golden_model_1.DPH [4]);
  nor (_18111_, _43000_, _18110_);
  nor (_18112_, _05297_, _18110_);
  nor (_18113_, _12816_, _08921_);
  or (_18114_, _18113_, _18112_);
  and (_18115_, _18114_, _03785_);
  nor (_18116_, _05777_, _08921_);
  or (_18118_, _18116_, _18112_);
  or (_18119_, _18118_, _06838_);
  nor (_18120_, _12841_, _08921_);
  or (_18121_, _18120_, _18112_);
  or (_18122_, _18121_, _04081_);
  and (_18123_, _05297_, \oc8051_golden_model_1.ACC [4]);
  or (_18124_, _18123_, _18112_);
  and (_18125_, _18124_, _04409_);
  nor (_18126_, _04409_, _18110_);
  or (_18127_, _18126_, _03610_);
  or (_18129_, _18127_, _18125_);
  and (_18130_, _18129_, _03996_);
  and (_18131_, _18130_, _18122_);
  and (_18132_, _18118_, _03723_);
  or (_18133_, _18132_, _03729_);
  or (_18134_, _18133_, _18131_);
  or (_18135_, _18124_, _03737_);
  and (_18136_, _18135_, _08848_);
  and (_18137_, _18136_, _18134_);
  or (_18138_, _08950_, \oc8051_golden_model_1.DPH [4]);
  nor (_18140_, _08951_, _08848_);
  and (_18141_, _18140_, _18138_);
  or (_18142_, _18141_, _18137_);
  and (_18143_, _18142_, _08832_);
  nor (_18144_, _03486_, _08832_);
  or (_18145_, _18144_, _07390_);
  or (_18146_, _18145_, _18143_);
  and (_18147_, _18146_, _18119_);
  or (_18148_, _18147_, _04481_);
  and (_18149_, _06730_, _05297_);
  or (_18151_, _18112_, _07400_);
  or (_18152_, _18151_, _18149_);
  and (_18153_, _18152_, _03589_);
  and (_18154_, _18153_, _18148_);
  nor (_18155_, _12933_, _08921_);
  or (_18156_, _18155_, _18112_);
  and (_18157_, _18156_, _03222_);
  or (_18158_, _18157_, _18154_);
  or (_18159_, _18158_, _08828_);
  and (_18160_, _12821_, _05297_);
  or (_18162_, _18112_, _07766_);
  or (_18163_, _18162_, _18160_);
  and (_18164_, _06298_, _05297_);
  or (_18165_, _18164_, _18112_);
  or (_18166_, _18165_, _05886_);
  and (_18167_, _18166_, _07778_);
  and (_18168_, _18167_, _18163_);
  and (_18169_, _18168_, _18159_);
  and (_18170_, _12817_, _05297_);
  or (_18171_, _18170_, _18112_);
  and (_18173_, _18171_, _03780_);
  or (_18174_, _18173_, _18169_);
  and (_18175_, _18174_, _07777_);
  or (_18176_, _18112_, _05825_);
  and (_18177_, _18165_, _03622_);
  and (_18178_, _18177_, _18176_);
  or (_18179_, _18178_, _18175_);
  and (_18180_, _18179_, _06828_);
  and (_18181_, _18124_, _03790_);
  and (_18182_, _18181_, _18176_);
  or (_18184_, _18182_, _03624_);
  or (_18185_, _18184_, _18180_);
  nor (_18186_, _12819_, _08921_);
  or (_18187_, _18112_, _07795_);
  or (_18188_, _18187_, _18186_);
  and (_18189_, _18188_, _07793_);
  and (_18190_, _18189_, _18185_);
  or (_18191_, _18190_, _18115_);
  and (_18192_, _18191_, _04246_);
  and (_18193_, _18121_, _03815_);
  or (_18195_, _18193_, _03447_);
  or (_18196_, _18195_, _18192_);
  and (_18197_, _13003_, _05297_);
  or (_18198_, _18112_, _03514_);
  or (_18199_, _18198_, _18197_);
  and (_18200_, _18199_, _43000_);
  and (_18201_, _18200_, _18196_);
  or (_18202_, _18201_, _18111_);
  and (_43513_, _18202_, _41806_);
  not (_18203_, \oc8051_golden_model_1.DPH [5]);
  nor (_18205_, _43000_, _18203_);
  nor (_18206_, _05297_, _18203_);
  nor (_18207_, _13146_, _08921_);
  or (_18208_, _18207_, _18206_);
  and (_18209_, _18208_, _03785_);
  nor (_18210_, _05469_, _08921_);
  or (_18211_, _18210_, _18206_);
  or (_18212_, _18211_, _06838_);
  nor (_18213_, _13014_, _08921_);
  or (_18214_, _18213_, _18206_);
  or (_18216_, _18214_, _04081_);
  and (_18217_, _05297_, \oc8051_golden_model_1.ACC [5]);
  or (_18218_, _18217_, _18206_);
  and (_18219_, _18218_, _04409_);
  nor (_18220_, _04409_, _18203_);
  or (_18221_, _18220_, _03610_);
  or (_18222_, _18221_, _18219_);
  and (_18223_, _18222_, _03996_);
  and (_18224_, _18223_, _18216_);
  and (_18225_, _18211_, _03723_);
  or (_18227_, _18225_, _03729_);
  or (_18228_, _18227_, _18224_);
  or (_18229_, _18218_, _03737_);
  and (_18230_, _18229_, _08848_);
  and (_18231_, _18230_, _18228_);
  or (_18232_, _08951_, \oc8051_golden_model_1.DPH [5]);
  nor (_18233_, _08952_, _08848_);
  and (_18234_, _18233_, _18232_);
  or (_18235_, _18234_, _18231_);
  and (_18236_, _18235_, _08832_);
  nor (_18238_, _03860_, _08832_);
  or (_18239_, _18238_, _07390_);
  or (_18240_, _18239_, _18236_);
  and (_18241_, _18240_, _18212_);
  or (_18242_, _18241_, _04481_);
  and (_18243_, _06684_, _05297_);
  or (_18244_, _18206_, _07400_);
  or (_18245_, _18244_, _18243_);
  and (_18246_, _18245_, _03589_);
  and (_18247_, _18246_, _18242_);
  nor (_18249_, _13127_, _08921_);
  or (_18250_, _18249_, _18206_);
  and (_18251_, _18250_, _03222_);
  or (_18252_, _18251_, _18247_);
  or (_18253_, _18252_, _08828_);
  and (_18254_, _13141_, _05297_);
  or (_18255_, _18206_, _07766_);
  or (_18256_, _18255_, _18254_);
  and (_18257_, _06306_, _05297_);
  or (_18258_, _18257_, _18206_);
  or (_18260_, _18258_, _05886_);
  and (_18261_, _18260_, _07778_);
  and (_18262_, _18261_, _18256_);
  and (_18263_, _18262_, _18253_);
  and (_18264_, _13147_, _05297_);
  or (_18265_, _18264_, _18206_);
  and (_18266_, _18265_, _03780_);
  or (_18267_, _18266_, _18263_);
  and (_18268_, _18267_, _07777_);
  or (_18269_, _18206_, _05518_);
  and (_18271_, _18258_, _03622_);
  and (_18272_, _18271_, _18269_);
  or (_18273_, _18272_, _18268_);
  and (_18274_, _18273_, _06828_);
  and (_18275_, _18218_, _03790_);
  and (_18276_, _18275_, _18269_);
  or (_18277_, _18276_, _03624_);
  or (_18278_, _18277_, _18274_);
  nor (_18279_, _13140_, _08921_);
  or (_18280_, _18206_, _07795_);
  or (_18282_, _18280_, _18279_);
  and (_18283_, _18282_, _07793_);
  and (_18284_, _18283_, _18278_);
  or (_18285_, _18284_, _18209_);
  and (_18286_, _18285_, _04246_);
  and (_18287_, _18214_, _03815_);
  or (_18288_, _18287_, _03447_);
  or (_18289_, _18288_, _18286_);
  and (_18290_, _13199_, _05297_);
  or (_18291_, _18206_, _03514_);
  or (_18293_, _18291_, _18290_);
  and (_18294_, _18293_, _43000_);
  and (_18295_, _18294_, _18289_);
  or (_18296_, _18295_, _18205_);
  and (_43514_, _18296_, _41806_);
  not (_18297_, \oc8051_golden_model_1.DPH [6]);
  nor (_18298_, _43000_, _18297_);
  nor (_18299_, _05297_, _18297_);
  nor (_18300_, _13352_, _08921_);
  or (_18301_, _18300_, _18299_);
  and (_18303_, _18301_, _03785_);
  nor (_18304_, _05363_, _08921_);
  or (_18305_, _18304_, _18299_);
  or (_18306_, _18305_, _06838_);
  nor (_18307_, _13242_, _08921_);
  or (_18308_, _18307_, _18299_);
  or (_18309_, _18308_, _04081_);
  and (_18310_, _05297_, \oc8051_golden_model_1.ACC [6]);
  or (_18311_, _18310_, _18299_);
  and (_18312_, _18311_, _04409_);
  nor (_18314_, _04409_, _18297_);
  or (_18315_, _18314_, _03610_);
  or (_18316_, _18315_, _18312_);
  and (_18317_, _18316_, _03996_);
  and (_18318_, _18317_, _18309_);
  and (_18319_, _18305_, _03723_);
  or (_18320_, _18319_, _03729_);
  or (_18321_, _18320_, _18318_);
  or (_18322_, _18311_, _03737_);
  and (_18323_, _18322_, _08848_);
  and (_18325_, _18323_, _18321_);
  or (_18326_, _08952_, \oc8051_golden_model_1.DPH [6]);
  nor (_18327_, _08953_, _08848_);
  and (_18328_, _18327_, _18326_);
  or (_18329_, _18328_, _18325_);
  and (_18330_, _18329_, _08832_);
  nor (_18331_, _08832_, _03549_);
  or (_18332_, _18331_, _07390_);
  or (_18333_, _18332_, _18330_);
  and (_18334_, _18333_, _18306_);
  or (_18336_, _18334_, _04481_);
  and (_18337_, _06455_, _05297_);
  or (_18338_, _18299_, _07400_);
  or (_18339_, _18338_, _18337_);
  and (_18340_, _18339_, _03589_);
  and (_18341_, _18340_, _18336_);
  nor (_18342_, _13332_, _08921_);
  or (_18343_, _18342_, _18299_);
  and (_18344_, _18343_, _03222_);
  or (_18345_, _18344_, _18341_);
  or (_18347_, _18345_, _08828_);
  and (_18348_, _13347_, _05297_);
  or (_18349_, _18299_, _07766_);
  or (_18350_, _18349_, _18348_);
  and (_18351_, _13339_, _05297_);
  or (_18352_, _18351_, _18299_);
  or (_18353_, _18352_, _05886_);
  and (_18354_, _18353_, _07778_);
  and (_18355_, _18354_, _18350_);
  and (_18356_, _18355_, _18347_);
  and (_18358_, _13353_, _05297_);
  or (_18359_, _18358_, _18299_);
  and (_18360_, _18359_, _03780_);
  or (_18361_, _18360_, _18356_);
  and (_18362_, _18361_, _07777_);
  or (_18363_, _18299_, _05412_);
  and (_18364_, _18352_, _03622_);
  and (_18365_, _18364_, _18363_);
  or (_18366_, _18365_, _18362_);
  and (_18367_, _18366_, _06828_);
  and (_18369_, _18311_, _03790_);
  and (_18370_, _18369_, _18363_);
  or (_18371_, _18370_, _03624_);
  or (_18372_, _18371_, _18367_);
  nor (_18373_, _13346_, _08921_);
  or (_18374_, _18299_, _07795_);
  or (_18375_, _18374_, _18373_);
  and (_18376_, _18375_, _07793_);
  and (_18377_, _18376_, _18372_);
  or (_18378_, _18377_, _18303_);
  and (_18380_, _18378_, _04246_);
  and (_18381_, _18308_, _03815_);
  or (_18382_, _18381_, _03447_);
  or (_18383_, _18382_, _18380_);
  and (_18384_, _13402_, _05297_);
  or (_18385_, _18299_, _03514_);
  or (_18386_, _18385_, _18384_);
  and (_18387_, _18386_, _43000_);
  and (_18388_, _18387_, _18383_);
  or (_18389_, _18388_, _18298_);
  and (_43515_, _18389_, _41806_);
  not (_18391_, \oc8051_golden_model_1.IE [0]);
  nor (_18392_, _05229_, _18391_);
  nor (_18393_, _05666_, _09021_);
  nor (_18394_, _18393_, _18392_);
  and (_18395_, _18394_, _03447_);
  and (_18396_, _12128_, _05229_);
  nor (_18397_, _18396_, _18392_);
  nor (_18398_, _18397_, _07778_);
  and (_18399_, _05229_, _06274_);
  nor (_18401_, _18399_, _18392_);
  and (_18402_, _18401_, _03601_);
  and (_18403_, _05229_, _04620_);
  nor (_18404_, _18403_, _18392_);
  and (_18405_, _18404_, _07390_);
  and (_18406_, _05229_, \oc8051_golden_model_1.ACC [0]);
  nor (_18407_, _18406_, _18392_);
  nor (_18408_, _18407_, _09029_);
  nor (_18409_, _04409_, _18391_);
  or (_18410_, _18409_, _18408_);
  and (_18412_, _18410_, _04081_);
  nor (_18413_, _18394_, _04081_);
  or (_18414_, _18413_, _18412_);
  and (_18415_, _18414_, _04055_);
  nor (_18416_, _05924_, _18391_);
  and (_18417_, _12021_, _05924_);
  nor (_18418_, _18417_, _18416_);
  nor (_18419_, _18418_, _04055_);
  nor (_18420_, _18419_, _18415_);
  nor (_18421_, _18420_, _03723_);
  nor (_18423_, _18404_, _03996_);
  or (_18424_, _18423_, _18421_);
  and (_18425_, _18424_, _03737_);
  nor (_18426_, _18407_, _03737_);
  or (_18427_, _18426_, _18425_);
  and (_18428_, _18427_, _03736_);
  and (_18429_, _18392_, _03714_);
  or (_18430_, _18429_, _18428_);
  and (_18431_, _18430_, _06840_);
  nor (_18432_, _18394_, _06840_);
  or (_18434_, _18432_, _18431_);
  and (_18435_, _18434_, _03710_);
  nor (_18436_, _12052_, _09059_);
  nor (_18437_, _18436_, _18416_);
  nor (_18438_, _18437_, _03710_);
  or (_18439_, _18438_, _07390_);
  nor (_18440_, _18439_, _18435_);
  nor (_18441_, _18440_, _18405_);
  nor (_18442_, _18441_, _04481_);
  and (_18443_, _06546_, _05229_);
  nor (_18445_, _18392_, _07400_);
  not (_18446_, _18445_);
  nor (_18447_, _18446_, _18443_);
  or (_18448_, _18447_, _03222_);
  nor (_18449_, _18448_, _18442_);
  nor (_18450_, _12109_, _09021_);
  nor (_18451_, _18450_, _18392_);
  nor (_18452_, _18451_, _03589_);
  or (_18453_, _18452_, _03601_);
  nor (_18454_, _18453_, _18449_);
  nor (_18456_, _18454_, _18402_);
  or (_18457_, _18456_, _03600_);
  and (_18458_, _12124_, _05229_);
  or (_18459_, _18458_, _18392_);
  or (_18460_, _18459_, _07766_);
  and (_18461_, _18460_, _07778_);
  and (_18462_, _18461_, _18457_);
  nor (_18463_, _18462_, _18398_);
  nor (_18464_, _18463_, _03622_);
  or (_18465_, _18401_, _07777_);
  nor (_18467_, _18465_, _18393_);
  nor (_18468_, _18467_, _18464_);
  nor (_18469_, _18468_, _03790_);
  and (_18470_, _12005_, _05229_);
  or (_18471_, _18470_, _18392_);
  and (_18472_, _18471_, _03790_);
  or (_18473_, _18472_, _18469_);
  and (_18474_, _18473_, _07795_);
  nor (_18475_, _12122_, _09021_);
  nor (_18476_, _18475_, _18392_);
  nor (_18478_, _18476_, _07795_);
  or (_18479_, _18478_, _18474_);
  and (_18480_, _18479_, _07793_);
  nor (_18481_, _12003_, _09021_);
  nor (_18482_, _18481_, _18392_);
  nor (_18483_, _18482_, _07793_);
  or (_18484_, _18483_, _18480_);
  and (_18485_, _18484_, _04246_);
  nor (_18486_, _18394_, _04246_);
  or (_18487_, _18486_, _18485_);
  and (_18489_, _18487_, _03823_);
  and (_18490_, _18392_, _03453_);
  nor (_18491_, _18490_, _03447_);
  not (_18492_, _18491_);
  nor (_18493_, _18492_, _18489_);
  nor (_18494_, _18493_, _18395_);
  or (_18495_, _18494_, _43004_);
  or (_18496_, _43000_, \oc8051_golden_model_1.IE [0]);
  and (_18497_, _18496_, _41806_);
  and (_43516_, _18497_, _18495_);
  not (_18499_, _03786_);
  not (_18500_, \oc8051_golden_model_1.IE [1]);
  nor (_18501_, _05229_, _18500_);
  and (_18502_, _06501_, _05229_);
  or (_18503_, _18502_, _18501_);
  and (_18504_, _18503_, _04481_);
  nor (_18505_, _05229_, \oc8051_golden_model_1.IE [1]);
  and (_18506_, _05229_, _03274_);
  nor (_18507_, _18506_, _18505_);
  and (_18508_, _18507_, _04409_);
  nor (_18510_, _04409_, _18500_);
  or (_18511_, _18510_, _18508_);
  and (_18512_, _18511_, _04081_);
  and (_18513_, _12213_, _05229_);
  nor (_18514_, _18513_, _18505_);
  and (_18515_, _18514_, _03610_);
  or (_18516_, _18515_, _18512_);
  and (_18517_, _18516_, _04055_);
  and (_18518_, _12224_, _05924_);
  nor (_18519_, _05924_, _18500_);
  or (_18521_, _18519_, _03723_);
  or (_18522_, _18521_, _18518_);
  and (_18523_, _18522_, _14265_);
  nor (_18524_, _18523_, _18517_);
  and (_18525_, _05229_, _06764_);
  nor (_18526_, _18525_, _18501_);
  and (_18527_, _18526_, _03723_);
  nor (_18528_, _18527_, _18524_);
  and (_18529_, _18528_, _03737_);
  and (_18530_, _18507_, _03729_);
  or (_18532_, _18530_, _18529_);
  and (_18533_, _18532_, _03736_);
  and (_18534_, _12211_, _05924_);
  nor (_18535_, _18534_, _18519_);
  nor (_18536_, _18535_, _03736_);
  or (_18537_, _18536_, _03719_);
  or (_18538_, _18537_, _18533_);
  and (_18539_, _18518_, _12239_);
  or (_18540_, _18519_, _06840_);
  or (_18541_, _18540_, _18539_);
  and (_18543_, _18541_, _18538_);
  and (_18544_, _18543_, _03710_);
  nor (_18545_, _12256_, _09059_);
  nor (_18546_, _18519_, _18545_);
  nor (_18547_, _18546_, _03710_);
  or (_18548_, _18547_, _07390_);
  nor (_18549_, _18548_, _18544_);
  and (_18550_, _18526_, _07390_);
  or (_18551_, _18550_, _04481_);
  nor (_18552_, _18551_, _18549_);
  or (_18554_, _18552_, _18504_);
  and (_18555_, _18554_, _03589_);
  nor (_18556_, _12313_, _09021_);
  nor (_18557_, _18556_, _18501_);
  nor (_18558_, _18557_, _03589_);
  nor (_18559_, _18558_, _18555_);
  nor (_18560_, _18559_, _08828_);
  not (_18561_, _18505_);
  nor (_18562_, _12327_, _09021_);
  nor (_18563_, _18562_, _07766_);
  and (_18565_, _05229_, _04303_);
  nor (_18566_, _18565_, _05886_);
  or (_18567_, _18566_, _18563_);
  and (_18568_, _18567_, _18561_);
  nor (_18569_, _18568_, _18560_);
  nor (_18570_, _18569_, _03780_);
  nor (_18571_, _12333_, _09021_);
  nor (_18572_, _18571_, _07778_);
  and (_18573_, _18572_, _18561_);
  nor (_18574_, _18573_, _18570_);
  nor (_18576_, _18574_, _03622_);
  nor (_18577_, _12207_, _09021_);
  nor (_18578_, _18577_, _07777_);
  and (_18579_, _18578_, _18561_);
  nor (_18580_, _18579_, _18576_);
  nor (_18581_, _18580_, _03790_);
  nor (_18582_, _18501_, _05618_);
  nor (_18583_, _18582_, _06828_);
  and (_18584_, _18583_, _18507_);
  nor (_18585_, _18584_, _18581_);
  or (_18587_, _18585_, _18499_);
  and (_18588_, _18565_, _05617_);
  nor (_18589_, _18588_, _07795_);
  and (_18590_, _18589_, _18561_);
  and (_18591_, _18506_, _05617_);
  or (_18592_, _18505_, _07793_);
  nor (_18593_, _18592_, _18591_);
  or (_18594_, _18593_, _03815_);
  nor (_18595_, _18594_, _18590_);
  and (_18596_, _18595_, _18587_);
  nor (_18598_, _18514_, _04246_);
  or (_18599_, _18598_, _03453_);
  nor (_18600_, _18599_, _18596_);
  nor (_18601_, _18535_, _03823_);
  or (_18602_, _18601_, _03447_);
  nor (_18603_, _18602_, _18600_);
  or (_18604_, _18501_, _03514_);
  nor (_18605_, _18604_, _18513_);
  nor (_18606_, _18605_, _18603_);
  or (_18607_, _18606_, _43004_);
  or (_18609_, _43000_, \oc8051_golden_model_1.IE [1]);
  and (_18610_, _18609_, _41806_);
  and (_43517_, _18610_, _18607_);
  not (_18611_, \oc8051_golden_model_1.IE [2]);
  nor (_18612_, _05229_, _18611_);
  and (_18613_, _05229_, _06332_);
  nor (_18614_, _18613_, _18612_);
  and (_18615_, _18614_, _03601_);
  nor (_18616_, _09021_, _04875_);
  nor (_18617_, _18616_, _18612_);
  and (_18619_, _18617_, _07390_);
  and (_18620_, _05229_, \oc8051_golden_model_1.ACC [2]);
  nor (_18621_, _18620_, _18612_);
  nor (_18622_, _18621_, _09029_);
  nor (_18623_, _04409_, _18611_);
  or (_18624_, _18623_, _18622_);
  and (_18625_, _18624_, _04081_);
  nor (_18626_, _12416_, _09021_);
  nor (_18627_, _18626_, _18612_);
  nor (_18628_, _18627_, _04081_);
  or (_18630_, _18628_, _18625_);
  and (_18631_, _18630_, _04055_);
  nor (_18632_, _05924_, _18611_);
  and (_18633_, _12411_, _05924_);
  nor (_18634_, _18633_, _18632_);
  nor (_18635_, _18634_, _04055_);
  or (_18636_, _18635_, _18631_);
  and (_18637_, _18636_, _03996_);
  nor (_18638_, _18617_, _03996_);
  or (_18639_, _18638_, _18637_);
  and (_18641_, _18639_, _03737_);
  nor (_18642_, _18621_, _03737_);
  or (_18643_, _18642_, _18641_);
  and (_18644_, _18643_, _03736_);
  and (_18645_, _12409_, _05924_);
  nor (_18646_, _18645_, _18632_);
  nor (_18647_, _18646_, _03736_);
  or (_18648_, _18647_, _03719_);
  or (_18649_, _18648_, _18644_);
  and (_18650_, _18633_, _12443_);
  or (_18652_, _18632_, _06840_);
  or (_18653_, _18652_, _18650_);
  and (_18654_, _18653_, _03710_);
  and (_18655_, _18654_, _18649_);
  nor (_18656_, _12461_, _09059_);
  nor (_18657_, _18656_, _18632_);
  nor (_18658_, _18657_, _03710_);
  nor (_18659_, _18658_, _07390_);
  not (_18660_, _18659_);
  nor (_18661_, _18660_, _18655_);
  nor (_18663_, _18661_, _18619_);
  nor (_18664_, _18663_, _04481_);
  and (_18665_, _06637_, _05229_);
  nor (_18666_, _18612_, _07400_);
  not (_18667_, _18666_);
  nor (_18668_, _18667_, _18665_);
  or (_18669_, _18668_, _03222_);
  nor (_18670_, _18669_, _18664_);
  nor (_18671_, _12519_, _09021_);
  nor (_18672_, _18612_, _18671_);
  nor (_18674_, _18672_, _03589_);
  or (_18675_, _18674_, _03601_);
  nor (_18676_, _18675_, _18670_);
  nor (_18677_, _18676_, _18615_);
  or (_18678_, _18677_, _03600_);
  and (_18679_, _12533_, _05229_);
  or (_18680_, _18679_, _18612_);
  or (_18681_, _18680_, _07766_);
  and (_18682_, _18681_, _07778_);
  and (_18683_, _18682_, _18678_);
  and (_18685_, _12539_, _05229_);
  nor (_18686_, _18685_, _18612_);
  nor (_18687_, _18686_, _07778_);
  nor (_18688_, _18687_, _18683_);
  nor (_18689_, _18688_, _03622_);
  nor (_18690_, _18612_, _05718_);
  not (_18691_, _18690_);
  nor (_18692_, _18614_, _07777_);
  and (_18693_, _18692_, _18691_);
  nor (_18694_, _18693_, _18689_);
  nor (_18696_, _18694_, _03790_);
  nor (_18697_, _18621_, _06828_);
  and (_18698_, _18697_, _18691_);
  or (_18699_, _18698_, _18696_);
  and (_18700_, _18699_, _07795_);
  nor (_18701_, _12532_, _09021_);
  nor (_18702_, _18701_, _18612_);
  nor (_18703_, _18702_, _07795_);
  or (_18704_, _18703_, _18700_);
  and (_18705_, _18704_, _07793_);
  nor (_18707_, _12538_, _09021_);
  nor (_18708_, _18707_, _18612_);
  nor (_18709_, _18708_, _07793_);
  or (_18710_, _18709_, _18705_);
  and (_18711_, _18710_, _04246_);
  nor (_18712_, _18627_, _04246_);
  or (_18713_, _18712_, _18711_);
  and (_18714_, _18713_, _03823_);
  nor (_18715_, _18646_, _03823_);
  or (_18716_, _18715_, _18714_);
  and (_18718_, _18716_, _03514_);
  and (_18719_, _12592_, _05229_);
  nor (_18720_, _18719_, _18612_);
  nor (_18721_, _18720_, _03514_);
  or (_18722_, _18721_, _18718_);
  or (_18723_, _18722_, _43004_);
  or (_18724_, _43000_, \oc8051_golden_model_1.IE [2]);
  and (_18725_, _18724_, _41806_);
  and (_43518_, _18725_, _18723_);
  not (_18726_, \oc8051_golden_model_1.IE [3]);
  nor (_18728_, _05229_, _18726_);
  and (_18729_, _05229_, _06276_);
  nor (_18730_, _18729_, _18728_);
  and (_18731_, _18730_, _03601_);
  nor (_18732_, _09021_, _05005_);
  nor (_18733_, _18732_, _18728_);
  and (_18734_, _18733_, _07390_);
  and (_18735_, _05229_, \oc8051_golden_model_1.ACC [3]);
  nor (_18736_, _18735_, _18728_);
  nor (_18737_, _18736_, _09029_);
  nor (_18739_, _04409_, _18726_);
  or (_18740_, _18739_, _18737_);
  and (_18741_, _18740_, _04081_);
  nor (_18742_, _12627_, _09021_);
  nor (_18743_, _18742_, _18728_);
  nor (_18744_, _18743_, _04081_);
  or (_18745_, _18744_, _18741_);
  and (_18746_, _18745_, _04055_);
  nor (_18747_, _05924_, _18726_);
  and (_18748_, _12631_, _05924_);
  nor (_18750_, _18748_, _18747_);
  nor (_18751_, _18750_, _04055_);
  or (_18752_, _18751_, _03723_);
  or (_18753_, _18752_, _18746_);
  nand (_18754_, _18733_, _03723_);
  and (_18755_, _18754_, _18753_);
  and (_18756_, _18755_, _03737_);
  nor (_18757_, _18736_, _03737_);
  or (_18758_, _18757_, _18756_);
  and (_18759_, _18758_, _03736_);
  and (_18761_, _12641_, _05924_);
  nor (_18762_, _18761_, _18747_);
  nor (_18763_, _18762_, _03736_);
  or (_18764_, _18763_, _03719_);
  or (_18765_, _18764_, _18759_);
  nor (_18766_, _18747_, _12648_);
  nor (_18767_, _18766_, _18750_);
  or (_18768_, _18767_, _06840_);
  and (_18769_, _18768_, _03710_);
  and (_18770_, _18769_, _18765_);
  nor (_18772_, _12612_, _09059_);
  nor (_18773_, _18772_, _18747_);
  nor (_18774_, _18773_, _03710_);
  nor (_18775_, _18774_, _07390_);
  not (_18776_, _18775_);
  nor (_18777_, _18776_, _18770_);
  nor (_18778_, _18777_, _18734_);
  nor (_18779_, _18778_, _04481_);
  and (_18780_, _06592_, _05229_);
  nor (_18781_, _18728_, _07400_);
  not (_18783_, _18781_);
  nor (_18784_, _18783_, _18780_);
  or (_18785_, _18784_, _03222_);
  nor (_18786_, _18785_, _18779_);
  nor (_18787_, _12718_, _09021_);
  nor (_18788_, _18728_, _18787_);
  nor (_18789_, _18788_, _03589_);
  or (_18790_, _18789_, _03601_);
  nor (_18791_, _18790_, _18786_);
  nor (_18792_, _18791_, _18731_);
  or (_18794_, _18792_, _03600_);
  and (_18795_, _12733_, _05229_);
  or (_18796_, _18795_, _18728_);
  or (_18797_, _18796_, _07766_);
  and (_18798_, _18797_, _07778_);
  and (_18799_, _18798_, _18794_);
  and (_18800_, _12739_, _05229_);
  nor (_18801_, _18800_, _18728_);
  nor (_18802_, _18801_, _07778_);
  nor (_18803_, _18802_, _18799_);
  nor (_18805_, _18803_, _03622_);
  nor (_18806_, _18728_, _05567_);
  not (_18807_, _18806_);
  nor (_18808_, _18730_, _07777_);
  and (_18809_, _18808_, _18807_);
  nor (_18810_, _18809_, _18805_);
  nor (_18811_, _18810_, _03790_);
  nor (_18812_, _18736_, _06828_);
  and (_18813_, _18812_, _18807_);
  nor (_18814_, _18813_, _03624_);
  not (_18816_, _18814_);
  nor (_18817_, _18816_, _18811_);
  nor (_18818_, _12732_, _09021_);
  or (_18819_, _18728_, _07795_);
  nor (_18820_, _18819_, _18818_);
  or (_18821_, _18820_, _03785_);
  nor (_18822_, _18821_, _18817_);
  nor (_18823_, _12738_, _09021_);
  nor (_18824_, _18823_, _18728_);
  nor (_18825_, _18824_, _07793_);
  or (_18827_, _18825_, _18822_);
  and (_18828_, _18827_, _04246_);
  nor (_18829_, _18743_, _04246_);
  or (_18830_, _18829_, _18828_);
  and (_18831_, _18830_, _03823_);
  nor (_18832_, _18762_, _03823_);
  or (_18833_, _18832_, _18831_);
  and (_18834_, _18833_, _03514_);
  and (_18835_, _12794_, _05229_);
  nor (_18836_, _18835_, _18728_);
  nor (_18838_, _18836_, _03514_);
  or (_18839_, _18838_, _18834_);
  or (_18840_, _18839_, _43004_);
  or (_18841_, _43000_, \oc8051_golden_model_1.IE [3]);
  and (_18842_, _18841_, _41806_);
  and (_43519_, _18842_, _18840_);
  not (_18843_, \oc8051_golden_model_1.IE [4]);
  nor (_18844_, _05229_, _18843_);
  nor (_18845_, _05777_, _09021_);
  nor (_18846_, _18845_, _18844_);
  and (_18848_, _18846_, _07390_);
  nor (_18849_, _05924_, _18843_);
  and (_18850_, _12827_, _05924_);
  nor (_18851_, _18850_, _18849_);
  nor (_18852_, _18851_, _03736_);
  and (_18853_, _05229_, \oc8051_golden_model_1.ACC [4]);
  nor (_18854_, _18853_, _18844_);
  nor (_18855_, _18854_, _09029_);
  nor (_18856_, _04409_, _18843_);
  or (_18857_, _18856_, _18855_);
  and (_18859_, _18857_, _04081_);
  nor (_18860_, _12841_, _09021_);
  nor (_18861_, _18860_, _18844_);
  nor (_18862_, _18861_, _04081_);
  or (_18863_, _18862_, _18859_);
  and (_18864_, _18863_, _04055_);
  and (_18865_, _12845_, _05924_);
  nor (_18866_, _18865_, _18849_);
  nor (_18867_, _18866_, _04055_);
  or (_18868_, _18867_, _03723_);
  or (_18870_, _18868_, _18864_);
  nand (_18871_, _18846_, _03723_);
  and (_18872_, _18871_, _18870_);
  and (_18873_, _18872_, _03737_);
  nor (_18874_, _18854_, _03737_);
  or (_18875_, _18874_, _18873_);
  and (_18876_, _18875_, _03736_);
  nor (_18877_, _18876_, _18852_);
  nor (_18878_, _18877_, _03719_);
  and (_18879_, _12861_, _05924_);
  nor (_18881_, _18879_, _18849_);
  nor (_18882_, _18881_, _06840_);
  nor (_18883_, _18882_, _18878_);
  nor (_18884_, _18883_, _03505_);
  nor (_18885_, _12825_, _09059_);
  nor (_18886_, _18885_, _18849_);
  nor (_18887_, _18886_, _03710_);
  nor (_18888_, _18887_, _07390_);
  not (_18889_, _18888_);
  nor (_18890_, _18889_, _18884_);
  nor (_18892_, _18890_, _18848_);
  nor (_18893_, _18892_, _04481_);
  and (_18894_, _06730_, _05229_);
  nor (_18895_, _18844_, _07400_);
  not (_18896_, _18895_);
  nor (_18897_, _18896_, _18894_);
  nor (_18898_, _18897_, _03222_);
  not (_18899_, _18898_);
  nor (_18900_, _18899_, _18893_);
  nor (_18901_, _12933_, _09021_);
  nor (_18903_, _18901_, _18844_);
  nor (_18904_, _18903_, _03589_);
  or (_18905_, _18904_, _08828_);
  or (_18906_, _18905_, _18900_);
  and (_18907_, _12821_, _05229_);
  or (_18908_, _18844_, _07766_);
  or (_18909_, _18908_, _18907_);
  and (_18910_, _06298_, _05229_);
  nor (_18911_, _18910_, _18844_);
  and (_18912_, _18911_, _03601_);
  nor (_18914_, _18912_, _03780_);
  and (_18915_, _18914_, _18909_);
  and (_18916_, _18915_, _18906_);
  and (_18917_, _12817_, _05229_);
  nor (_18918_, _18917_, _18844_);
  nor (_18919_, _18918_, _07778_);
  nor (_18920_, _18919_, _18916_);
  nor (_18921_, _18920_, _03622_);
  nor (_18922_, _18844_, _05825_);
  not (_18923_, _18922_);
  nor (_18925_, _18911_, _07777_);
  and (_18926_, _18925_, _18923_);
  nor (_18927_, _18926_, _18921_);
  nor (_18928_, _18927_, _03790_);
  nor (_18929_, _18854_, _06828_);
  and (_18930_, _18929_, _18923_);
  or (_18931_, _18930_, _18928_);
  and (_18932_, _18931_, _07795_);
  nor (_18933_, _12819_, _09021_);
  nor (_18934_, _18933_, _18844_);
  nor (_18936_, _18934_, _07795_);
  or (_18937_, _18936_, _18932_);
  and (_18938_, _18937_, _07793_);
  nor (_18939_, _12816_, _09021_);
  nor (_18940_, _18939_, _18844_);
  nor (_18941_, _18940_, _07793_);
  or (_18942_, _18941_, _18938_);
  and (_18943_, _18942_, _04246_);
  nor (_18944_, _18861_, _04246_);
  or (_18945_, _18944_, _18943_);
  and (_18947_, _18945_, _03823_);
  nor (_18948_, _18851_, _03823_);
  or (_18949_, _18948_, _18947_);
  and (_18950_, _18949_, _03514_);
  and (_18951_, _13003_, _05229_);
  nor (_18952_, _18951_, _18844_);
  nor (_18953_, _18952_, _03514_);
  or (_18954_, _18953_, _18950_);
  or (_18955_, _18954_, _43004_);
  or (_18956_, _43000_, \oc8051_golden_model_1.IE [4]);
  and (_18958_, _18956_, _41806_);
  and (_43520_, _18958_, _18955_);
  not (_18959_, \oc8051_golden_model_1.IE [5]);
  nor (_18960_, _05229_, _18959_);
  and (_18961_, _06684_, _05229_);
  or (_18962_, _18961_, _18960_);
  and (_18963_, _18962_, _04481_);
  and (_18964_, _05229_, \oc8051_golden_model_1.ACC [5]);
  nor (_18965_, _18964_, _18960_);
  nor (_18966_, _18965_, _09029_);
  nor (_18968_, _04409_, _18959_);
  or (_18969_, _18968_, _18966_);
  and (_18970_, _18969_, _04081_);
  nor (_18971_, _13014_, _09021_);
  nor (_18972_, _18971_, _18960_);
  nor (_18973_, _18972_, _04081_);
  or (_18974_, _18973_, _18970_);
  and (_18975_, _18974_, _04055_);
  nor (_18976_, _05924_, _18959_);
  and (_18977_, _13037_, _05924_);
  nor (_18979_, _18977_, _18976_);
  nor (_18980_, _18979_, _04055_);
  or (_18981_, _18980_, _03723_);
  or (_18982_, _18981_, _18975_);
  nor (_18983_, _05469_, _09021_);
  nor (_18984_, _18983_, _18960_);
  nand (_18985_, _18984_, _03723_);
  and (_18986_, _18985_, _18982_);
  and (_18987_, _18986_, _03737_);
  nor (_18988_, _18965_, _03737_);
  or (_18990_, _18988_, _18987_);
  and (_18991_, _18990_, _03736_);
  and (_18992_, _13047_, _05924_);
  nor (_18993_, _18992_, _18976_);
  nor (_18994_, _18993_, _03736_);
  or (_18995_, _18994_, _03719_);
  or (_18996_, _18995_, _18991_);
  nor (_18997_, _18976_, _13054_);
  nor (_18998_, _18997_, _18979_);
  or (_18999_, _18998_, _06840_);
  and (_19001_, _18999_, _03710_);
  and (_19002_, _19001_, _18996_);
  nor (_19003_, _13020_, _09059_);
  nor (_19004_, _19003_, _18976_);
  nor (_19005_, _19004_, _03710_);
  nor (_19006_, _19005_, _07390_);
  not (_19007_, _19006_);
  nor (_19008_, _19007_, _19002_);
  and (_19009_, _18984_, _07390_);
  or (_19010_, _19009_, _04481_);
  nor (_19012_, _19010_, _19008_);
  or (_19013_, _19012_, _18963_);
  and (_19014_, _19013_, _03589_);
  nor (_19015_, _13127_, _09021_);
  nor (_19016_, _19015_, _18960_);
  nor (_19017_, _19016_, _03589_);
  or (_19018_, _19017_, _08828_);
  or (_19019_, _19018_, _19014_);
  and (_19020_, _13141_, _05229_);
  or (_19021_, _18960_, _07766_);
  or (_19023_, _19021_, _19020_);
  and (_19024_, _06306_, _05229_);
  nor (_19025_, _19024_, _18960_);
  and (_19026_, _19025_, _03601_);
  nor (_19027_, _19026_, _03780_);
  and (_19028_, _19027_, _19023_);
  and (_19029_, _19028_, _19019_);
  and (_19030_, _13147_, _05229_);
  nor (_19031_, _19030_, _18960_);
  nor (_19032_, _19031_, _07778_);
  nor (_19034_, _19032_, _19029_);
  nor (_19035_, _19034_, _03622_);
  nor (_19036_, _18960_, _05518_);
  not (_19037_, _19036_);
  nor (_19038_, _19025_, _07777_);
  and (_19039_, _19038_, _19037_);
  nor (_19040_, _19039_, _19035_);
  nor (_19041_, _19040_, _03790_);
  nor (_19042_, _18965_, _06828_);
  and (_19043_, _19042_, _19037_);
  or (_19045_, _19043_, _19041_);
  and (_19046_, _19045_, _07795_);
  nor (_19047_, _13140_, _09021_);
  nor (_19048_, _19047_, _18960_);
  nor (_19049_, _19048_, _07795_);
  or (_19050_, _19049_, _19046_);
  and (_19051_, _19050_, _07793_);
  nor (_19052_, _13146_, _09021_);
  nor (_19053_, _19052_, _18960_);
  nor (_19054_, _19053_, _07793_);
  or (_19056_, _19054_, _19051_);
  and (_19057_, _19056_, _04246_);
  nor (_19058_, _18972_, _04246_);
  or (_19059_, _19058_, _19057_);
  and (_19060_, _19059_, _03823_);
  nor (_19061_, _18993_, _03823_);
  or (_19062_, _19061_, _19060_);
  and (_19063_, _19062_, _03514_);
  and (_19064_, _13199_, _05229_);
  nor (_19065_, _19064_, _18960_);
  nor (_19067_, _19065_, _03514_);
  or (_19068_, _19067_, _19063_);
  or (_19069_, _19068_, _43004_);
  or (_19070_, _43000_, \oc8051_golden_model_1.IE [5]);
  and (_19071_, _19070_, _41806_);
  and (_43521_, _19071_, _19069_);
  not (_19072_, \oc8051_golden_model_1.IE [6]);
  nor (_19073_, _05229_, _19072_);
  and (_19074_, _06455_, _05229_);
  or (_19075_, _19074_, _19073_);
  and (_19077_, _19075_, _04481_);
  and (_19078_, _05229_, \oc8051_golden_model_1.ACC [6]);
  nor (_19079_, _19078_, _19073_);
  nor (_19080_, _19079_, _09029_);
  nor (_19081_, _04409_, _19072_);
  or (_19082_, _19081_, _19080_);
  and (_19083_, _19082_, _04081_);
  nor (_19084_, _13242_, _09021_);
  nor (_19085_, _19084_, _19073_);
  nor (_19086_, _19085_, _04081_);
  or (_19088_, _19086_, _19083_);
  and (_19089_, _19088_, _04055_);
  nor (_19090_, _05924_, _19072_);
  and (_19091_, _13229_, _05924_);
  nor (_19092_, _19091_, _19090_);
  nor (_19093_, _19092_, _04055_);
  or (_19094_, _19093_, _03723_);
  or (_19095_, _19094_, _19089_);
  nor (_19096_, _05363_, _09021_);
  nor (_19097_, _19096_, _19073_);
  nand (_19099_, _19097_, _03723_);
  and (_19100_, _19099_, _19095_);
  and (_19101_, _19100_, _03737_);
  nor (_19102_, _19079_, _03737_);
  or (_19103_, _19102_, _19101_);
  and (_19104_, _19103_, _03736_);
  and (_19105_, _13253_, _05924_);
  nor (_19106_, _19105_, _19090_);
  nor (_19107_, _19106_, _03736_);
  or (_19108_, _19107_, _19104_);
  and (_19110_, _19108_, _06840_);
  nor (_19111_, _19090_, _13260_);
  nor (_19112_, _19111_, _19092_);
  and (_19113_, _19112_, _03719_);
  or (_19114_, _19113_, _19110_);
  and (_19115_, _19114_, _03710_);
  nor (_19116_, _13226_, _09059_);
  nor (_19117_, _19116_, _19090_);
  nor (_19118_, _19117_, _03710_);
  nor (_19119_, _19118_, _07390_);
  not (_19121_, _19119_);
  nor (_19122_, _19121_, _19115_);
  and (_19123_, _19097_, _07390_);
  or (_19124_, _19123_, _04481_);
  nor (_19125_, _19124_, _19122_);
  or (_19126_, _19125_, _19077_);
  and (_19127_, _19126_, _03589_);
  nor (_19128_, _13332_, _09021_);
  nor (_19129_, _19128_, _19073_);
  nor (_19130_, _19129_, _03589_);
  or (_19132_, _19130_, _08828_);
  or (_19133_, _19132_, _19127_);
  and (_19134_, _13347_, _05229_);
  or (_19135_, _19073_, _07766_);
  or (_19136_, _19135_, _19134_);
  and (_19137_, _13339_, _05229_);
  nor (_19138_, _19137_, _19073_);
  and (_19139_, _19138_, _03601_);
  nor (_19140_, _19139_, _03780_);
  and (_19141_, _19140_, _19136_);
  and (_19143_, _19141_, _19133_);
  and (_19144_, _13353_, _05229_);
  nor (_19145_, _19144_, _19073_);
  nor (_19146_, _19145_, _07778_);
  nor (_19147_, _19146_, _19143_);
  nor (_19148_, _19147_, _03622_);
  nor (_19149_, _19073_, _05412_);
  not (_19150_, _19149_);
  nor (_19151_, _19138_, _07777_);
  and (_19152_, _19151_, _19150_);
  nor (_19154_, _19152_, _19148_);
  nor (_19155_, _19154_, _03790_);
  nor (_19156_, _19079_, _06828_);
  and (_19157_, _19156_, _19150_);
  nor (_19158_, _19157_, _03624_);
  not (_19159_, _19158_);
  nor (_19160_, _19159_, _19155_);
  nor (_19161_, _13346_, _09021_);
  or (_19162_, _19073_, _07795_);
  nor (_19163_, _19162_, _19161_);
  or (_19165_, _19163_, _03785_);
  nor (_19166_, _19165_, _19160_);
  nor (_19167_, _13352_, _09021_);
  nor (_19168_, _19167_, _19073_);
  nor (_19169_, _19168_, _07793_);
  or (_19170_, _19169_, _19166_);
  and (_19171_, _19170_, _04246_);
  nor (_19172_, _19085_, _04246_);
  or (_19173_, _19172_, _19171_);
  and (_19174_, _19173_, _03823_);
  nor (_19176_, _19106_, _03823_);
  or (_19177_, _19176_, _19174_);
  and (_19178_, _19177_, _03514_);
  and (_19179_, _13402_, _05229_);
  nor (_19180_, _19179_, _19073_);
  nor (_19181_, _19180_, _03514_);
  or (_19182_, _19181_, _19178_);
  or (_19183_, _19182_, _43004_);
  or (_19184_, _43000_, \oc8051_golden_model_1.IE [6]);
  and (_19185_, _19184_, _41806_);
  and (_43522_, _19185_, _19183_);
  not (_19187_, \oc8051_golden_model_1.IP [0]);
  nor (_19188_, _05251_, _19187_);
  and (_19189_, _12128_, _05251_);
  nor (_19190_, _19189_, _19188_);
  nor (_19191_, _19190_, _07778_);
  and (_19192_, _05251_, _06274_);
  nor (_19193_, _19192_, _19188_);
  and (_19194_, _19193_, _03601_);
  and (_19195_, _05251_, _04620_);
  nor (_19197_, _19195_, _19188_);
  and (_19198_, _19197_, _07390_);
  nor (_19199_, _05666_, _09129_);
  nor (_19200_, _19199_, _19188_);
  nor (_19201_, _19200_, _04081_);
  nor (_19202_, _04409_, _19187_);
  and (_19203_, _05251_, \oc8051_golden_model_1.ACC [0]);
  nor (_19204_, _19203_, _19188_);
  nor (_19205_, _19204_, _09029_);
  nor (_19206_, _19205_, _19202_);
  nor (_19208_, _19206_, _03610_);
  or (_19209_, _19208_, _03715_);
  nor (_19210_, _19209_, _19201_);
  and (_19211_, _12021_, _05908_);
  nor (_19212_, _05908_, _19187_);
  or (_19213_, _19212_, _04055_);
  nor (_19214_, _19213_, _19211_);
  or (_19215_, _19214_, _03723_);
  nor (_19216_, _19215_, _19210_);
  nor (_19217_, _19197_, _03996_);
  or (_19219_, _19217_, _19216_);
  and (_19220_, _19219_, _03737_);
  nor (_19221_, _19204_, _03737_);
  or (_19222_, _19221_, _19220_);
  and (_19223_, _19222_, _03736_);
  and (_19224_, _19188_, _03714_);
  or (_19225_, _19224_, _19223_);
  and (_19226_, _19225_, _06840_);
  nor (_19227_, _19200_, _06840_);
  or (_19228_, _19227_, _19226_);
  and (_19230_, _19228_, _03710_);
  nor (_19231_, _12052_, _09166_);
  nor (_19232_, _19231_, _19212_);
  nor (_19233_, _19232_, _03710_);
  or (_19234_, _19233_, _07390_);
  nor (_19235_, _19234_, _19230_);
  nor (_19236_, _19235_, _19198_);
  nor (_19237_, _19236_, _04481_);
  and (_19238_, _06546_, _05251_);
  nor (_19239_, _19188_, _07400_);
  not (_19241_, _19239_);
  nor (_19242_, _19241_, _19238_);
  or (_19243_, _19242_, _03222_);
  nor (_19244_, _19243_, _19237_);
  nor (_19245_, _12109_, _09129_);
  nor (_19246_, _19245_, _19188_);
  nor (_19247_, _19246_, _03589_);
  or (_19248_, _19247_, _03601_);
  nor (_19249_, _19248_, _19244_);
  nor (_19250_, _19249_, _19194_);
  or (_19252_, _19250_, _03600_);
  and (_19253_, _12124_, _05251_);
  or (_19254_, _19253_, _19188_);
  or (_19255_, _19254_, _07766_);
  and (_19256_, _19255_, _07778_);
  and (_19257_, _19256_, _19252_);
  nor (_19258_, _19257_, _19191_);
  nor (_19259_, _19258_, _03622_);
  or (_19260_, _19193_, _07777_);
  nor (_19261_, _19260_, _19199_);
  nor (_19263_, _19261_, _19259_);
  nor (_19264_, _19263_, _03790_);
  and (_19265_, _12005_, _05251_);
  or (_19266_, _19265_, _19188_);
  and (_19267_, _19266_, _03790_);
  or (_19268_, _19267_, _19264_);
  and (_19269_, _19268_, _07795_);
  nor (_19270_, _12122_, _09129_);
  nor (_19271_, _19270_, _19188_);
  nor (_19272_, _19271_, _07795_);
  or (_19274_, _19272_, _19269_);
  and (_19275_, _19274_, _07793_);
  nor (_19276_, _12003_, _09129_);
  nor (_19277_, _19276_, _19188_);
  nor (_19278_, _19277_, _07793_);
  or (_19279_, _19278_, _19275_);
  and (_19280_, _19279_, _04246_);
  nor (_19281_, _19200_, _04246_);
  or (_19282_, _19281_, _19280_);
  and (_19283_, _19282_, _03823_);
  and (_19285_, _19188_, _03453_);
  or (_19286_, _19285_, _19283_);
  and (_19287_, _19286_, _03514_);
  nor (_19288_, _19200_, _03514_);
  or (_19289_, _19288_, _19287_);
  or (_19290_, _19289_, _43004_);
  or (_19291_, _43000_, \oc8051_golden_model_1.IP [0]);
  and (_19292_, _19291_, _41806_);
  and (_43525_, _19292_, _19290_);
  not (_19293_, \oc8051_golden_model_1.IP [1]);
  nor (_19295_, _05251_, _19293_);
  and (_19296_, _06501_, _05251_);
  or (_19297_, _19296_, _19295_);
  and (_19298_, _19297_, _04481_);
  nor (_19299_, _05251_, \oc8051_golden_model_1.IP [1]);
  and (_19300_, _05251_, _03274_);
  nor (_19301_, _19300_, _19299_);
  and (_19302_, _19301_, _04409_);
  nor (_19303_, _04409_, _19293_);
  or (_19304_, _19303_, _19302_);
  and (_19306_, _19304_, _04081_);
  and (_19307_, _12213_, _05251_);
  nor (_19308_, _19307_, _19299_);
  and (_19309_, _19308_, _03610_);
  or (_19310_, _19309_, _19306_);
  and (_19311_, _19310_, _04055_);
  and (_19312_, _12224_, _05908_);
  nor (_19313_, _05908_, _19293_);
  or (_19314_, _19313_, _03723_);
  or (_19315_, _19314_, _19312_);
  and (_19317_, _19315_, _14265_);
  nor (_19318_, _19317_, _19311_);
  and (_19319_, _05251_, _06764_);
  nor (_19320_, _19319_, _19295_);
  and (_19321_, _19320_, _03723_);
  nor (_19322_, _19321_, _19318_);
  and (_19323_, _19322_, _03737_);
  and (_19324_, _19301_, _03729_);
  or (_19325_, _19324_, _19323_);
  and (_19326_, _19325_, _03736_);
  and (_19328_, _12211_, _05908_);
  nor (_19329_, _19328_, _19313_);
  nor (_19330_, _19329_, _03736_);
  or (_19331_, _19330_, _19326_);
  and (_19332_, _19331_, _06840_);
  and (_19333_, _19312_, _12239_);
  or (_19334_, _19333_, _19313_);
  and (_19335_, _19334_, _03719_);
  or (_19336_, _19335_, _19332_);
  and (_19337_, _19336_, _03710_);
  nor (_19339_, _12256_, _09166_);
  nor (_19340_, _19313_, _19339_);
  nor (_19341_, _19340_, _03710_);
  or (_19342_, _19341_, _07390_);
  nor (_19343_, _19342_, _19337_);
  and (_19344_, _19320_, _07390_);
  or (_19345_, _19344_, _04481_);
  nor (_19346_, _19345_, _19343_);
  or (_19347_, _19346_, _19298_);
  and (_19348_, _19347_, _03589_);
  nor (_19350_, _12313_, _09129_);
  nor (_19351_, _19350_, _19295_);
  nor (_19352_, _19351_, _03589_);
  nor (_19353_, _19352_, _19348_);
  nor (_19354_, _19353_, _08828_);
  nor (_19355_, _12327_, _09129_);
  nor (_19356_, _19355_, _07766_);
  and (_19357_, _05251_, _04303_);
  nor (_19358_, _19357_, _05886_);
  nor (_19359_, _19358_, _19356_);
  nor (_19361_, _19359_, _19299_);
  nor (_19362_, _19361_, _19354_);
  nor (_19363_, _19362_, _03780_);
  not (_19364_, _19299_);
  nor (_19365_, _12333_, _09129_);
  nor (_19366_, _19365_, _07778_);
  and (_19367_, _19366_, _19364_);
  nor (_19368_, _19367_, _19363_);
  nor (_19369_, _19368_, _03622_);
  nor (_19370_, _12207_, _09129_);
  nor (_19372_, _19370_, _07777_);
  and (_19373_, _19372_, _19364_);
  nor (_19374_, _19373_, _19369_);
  nor (_19375_, _19374_, _03790_);
  nor (_19376_, _19295_, _05618_);
  nor (_19377_, _19376_, _06828_);
  and (_19378_, _19377_, _19301_);
  nor (_19379_, _19378_, _19375_);
  or (_19380_, _19379_, _18499_);
  and (_19381_, _19357_, _05617_);
  or (_19383_, _19299_, _07795_);
  or (_19384_, _19383_, _19381_);
  and (_19385_, _19300_, _05617_);
  or (_19386_, _19299_, _07793_);
  or (_19387_, _19386_, _19385_);
  and (_19388_, _19387_, _04246_);
  and (_19389_, _19388_, _19384_);
  and (_19390_, _19389_, _19380_);
  nor (_19391_, _19308_, _04246_);
  or (_19392_, _19391_, _03453_);
  nor (_19394_, _19392_, _19390_);
  nor (_19395_, _19329_, _03823_);
  or (_19396_, _19395_, _03447_);
  nor (_19397_, _19396_, _19394_);
  or (_19398_, _19295_, _03514_);
  nor (_19399_, _19398_, _19307_);
  nor (_19400_, _19399_, _19397_);
  or (_19401_, _19400_, _43004_);
  or (_19402_, _43000_, \oc8051_golden_model_1.IP [1]);
  and (_19403_, _19402_, _41806_);
  and (_43526_, _19403_, _19401_);
  not (_19405_, \oc8051_golden_model_1.IP [2]);
  nor (_19406_, _05251_, _19405_);
  and (_19407_, _05251_, _06332_);
  nor (_19408_, _19407_, _19406_);
  and (_19409_, _19408_, _03601_);
  nor (_19410_, _09129_, _04875_);
  nor (_19411_, _19410_, _19406_);
  and (_19412_, _19411_, _07390_);
  and (_19413_, _05251_, \oc8051_golden_model_1.ACC [2]);
  nor (_19415_, _19413_, _19406_);
  nor (_19416_, _19415_, _09029_);
  nor (_19417_, _04409_, _19405_);
  or (_19418_, _19417_, _19416_);
  and (_19419_, _19418_, _04081_);
  nor (_19420_, _12416_, _09129_);
  nor (_19421_, _19420_, _19406_);
  nor (_19422_, _19421_, _04081_);
  or (_19423_, _19422_, _19419_);
  and (_19424_, _19423_, _04055_);
  nor (_19426_, _05908_, _19405_);
  and (_19427_, _12411_, _05908_);
  nor (_19428_, _19427_, _19426_);
  nor (_19429_, _19428_, _04055_);
  or (_19430_, _19429_, _19424_);
  and (_19431_, _19430_, _03996_);
  nor (_19432_, _19411_, _03996_);
  or (_19433_, _19432_, _19431_);
  and (_19434_, _19433_, _03737_);
  nor (_19435_, _19415_, _03737_);
  or (_19437_, _19435_, _19434_);
  and (_19438_, _19437_, _03736_);
  and (_19439_, _12409_, _05908_);
  nor (_19440_, _19439_, _19426_);
  nor (_19441_, _19440_, _03736_);
  or (_19442_, _19441_, _03719_);
  or (_19443_, _19442_, _19438_);
  and (_19444_, _19427_, _12443_);
  or (_19445_, _19426_, _06840_);
  or (_19446_, _19445_, _19444_);
  and (_19448_, _19446_, _03710_);
  and (_19449_, _19448_, _19443_);
  nor (_19450_, _12461_, _09166_);
  nor (_19451_, _19450_, _19426_);
  nor (_19452_, _19451_, _03710_);
  nor (_19453_, _19452_, _07390_);
  not (_19454_, _19453_);
  nor (_19455_, _19454_, _19449_);
  nor (_19456_, _19455_, _19412_);
  nor (_19457_, _19456_, _04481_);
  and (_19459_, _06637_, _05251_);
  nor (_19460_, _19406_, _07400_);
  not (_19461_, _19460_);
  nor (_19462_, _19461_, _19459_);
  or (_19463_, _19462_, _03222_);
  nor (_19464_, _19463_, _19457_);
  nor (_19465_, _12519_, _09129_);
  nor (_19466_, _19406_, _19465_);
  nor (_19467_, _19466_, _03589_);
  or (_19468_, _19467_, _03601_);
  nor (_19470_, _19468_, _19464_);
  nor (_19471_, _19470_, _19409_);
  or (_19472_, _19471_, _03600_);
  and (_19473_, _12533_, _05251_);
  or (_19474_, _19473_, _19406_);
  or (_19475_, _19474_, _07766_);
  and (_19476_, _19475_, _07778_);
  and (_19477_, _19476_, _19472_);
  and (_19478_, _12539_, _05251_);
  nor (_19479_, _19478_, _19406_);
  nor (_19481_, _19479_, _07778_);
  nor (_19482_, _19481_, _19477_);
  nor (_19483_, _19482_, _03622_);
  nor (_19484_, _19406_, _05718_);
  not (_19485_, _19484_);
  nor (_19486_, _19408_, _07777_);
  and (_19487_, _19486_, _19485_);
  nor (_19488_, _19487_, _19483_);
  nor (_19489_, _19488_, _03790_);
  nor (_19490_, _19415_, _06828_);
  and (_19492_, _19490_, _19485_);
  nor (_19493_, _19492_, _03624_);
  not (_19494_, _19493_);
  nor (_19495_, _19494_, _19489_);
  nor (_19496_, _12532_, _09129_);
  or (_19497_, _19406_, _07795_);
  nor (_19498_, _19497_, _19496_);
  or (_19499_, _19498_, _03785_);
  nor (_19500_, _19499_, _19495_);
  nor (_19501_, _12538_, _09129_);
  nor (_19503_, _19501_, _19406_);
  nor (_19504_, _19503_, _07793_);
  or (_19505_, _19504_, _19500_);
  and (_19506_, _19505_, _04246_);
  nor (_19507_, _19421_, _04246_);
  or (_19508_, _19507_, _19506_);
  and (_19509_, _19508_, _03823_);
  nor (_19510_, _19440_, _03823_);
  or (_19511_, _19510_, _19509_);
  and (_19512_, _19511_, _03514_);
  and (_19514_, _12592_, _05251_);
  nor (_19515_, _19514_, _19406_);
  nor (_19516_, _19515_, _03514_);
  or (_19517_, _19516_, _19512_);
  or (_19518_, _19517_, _43004_);
  or (_19519_, _43000_, \oc8051_golden_model_1.IP [2]);
  and (_19520_, _19519_, _41806_);
  and (_43527_, _19520_, _19518_);
  not (_19521_, \oc8051_golden_model_1.IP [3]);
  nor (_19522_, _05251_, _19521_);
  and (_19524_, _05251_, _06276_);
  nor (_19525_, _19524_, _19522_);
  and (_19526_, _19525_, _03601_);
  nor (_19527_, _09129_, _05005_);
  nor (_19528_, _19527_, _19522_);
  and (_19529_, _19528_, _07390_);
  and (_19530_, _05251_, \oc8051_golden_model_1.ACC [3]);
  nor (_19531_, _19530_, _19522_);
  nor (_19532_, _19531_, _09029_);
  nor (_19533_, _04409_, _19521_);
  or (_19535_, _19533_, _19532_);
  and (_19536_, _19535_, _04081_);
  nor (_19537_, _12627_, _09129_);
  nor (_19538_, _19537_, _19522_);
  nor (_19539_, _19538_, _04081_);
  or (_19540_, _19539_, _19536_);
  and (_19541_, _19540_, _04055_);
  nor (_19542_, _05908_, _19521_);
  and (_19543_, _12631_, _05908_);
  nor (_19544_, _19543_, _19542_);
  nor (_19546_, _19544_, _04055_);
  or (_19547_, _19546_, _03723_);
  or (_19548_, _19547_, _19541_);
  nand (_19549_, _19528_, _03723_);
  and (_19550_, _19549_, _19548_);
  and (_19551_, _19550_, _03737_);
  nor (_19552_, _19531_, _03737_);
  or (_19553_, _19552_, _19551_);
  and (_19554_, _19553_, _03736_);
  and (_19555_, _12641_, _05908_);
  nor (_19557_, _19555_, _19542_);
  nor (_19558_, _19557_, _03736_);
  or (_19559_, _19558_, _19554_);
  and (_19560_, _19559_, _06840_);
  nor (_19561_, _19542_, _12648_);
  nor (_19562_, _19561_, _19544_);
  and (_19563_, _19562_, _03719_);
  or (_19564_, _19563_, _19560_);
  and (_19565_, _19564_, _03710_);
  nor (_19566_, _12612_, _09166_);
  nor (_19568_, _19566_, _19542_);
  nor (_19569_, _19568_, _03710_);
  nor (_19570_, _19569_, _07390_);
  not (_19571_, _19570_);
  nor (_19572_, _19571_, _19565_);
  nor (_19573_, _19572_, _19529_);
  nor (_19574_, _19573_, _04481_);
  and (_19575_, _06592_, _05251_);
  nor (_19576_, _19522_, _07400_);
  not (_19577_, _19576_);
  nor (_19579_, _19577_, _19575_);
  or (_19580_, _19579_, _03222_);
  nor (_19581_, _19580_, _19574_);
  nor (_19582_, _12718_, _09129_);
  nor (_19583_, _19522_, _19582_);
  nor (_19584_, _19583_, _03589_);
  or (_19585_, _19584_, _03601_);
  nor (_19586_, _19585_, _19581_);
  nor (_19587_, _19586_, _19526_);
  or (_19588_, _19587_, _03600_);
  and (_19590_, _12733_, _05251_);
  or (_19591_, _19590_, _19522_);
  or (_19592_, _19591_, _07766_);
  and (_19593_, _19592_, _07778_);
  and (_19594_, _19593_, _19588_);
  and (_19595_, _12739_, _05251_);
  nor (_19596_, _19595_, _19522_);
  nor (_19597_, _19596_, _07778_);
  nor (_19598_, _19597_, _19594_);
  nor (_19599_, _19598_, _03622_);
  nor (_19601_, _19522_, _05567_);
  not (_19602_, _19601_);
  nor (_19603_, _19525_, _07777_);
  and (_19604_, _19603_, _19602_);
  nor (_19605_, _19604_, _19599_);
  nor (_19606_, _19605_, _03790_);
  nor (_19607_, _19531_, _06828_);
  and (_19608_, _19607_, _19602_);
  nor (_19609_, _19608_, _03624_);
  not (_19610_, _19609_);
  nor (_19612_, _19610_, _19606_);
  nor (_19613_, _12732_, _09129_);
  or (_19614_, _19522_, _07795_);
  nor (_19615_, _19614_, _19613_);
  or (_19616_, _19615_, _03785_);
  nor (_19617_, _19616_, _19612_);
  nor (_19618_, _12738_, _09129_);
  nor (_19619_, _19618_, _19522_);
  nor (_19620_, _19619_, _07793_);
  or (_19621_, _19620_, _19617_);
  and (_19623_, _19621_, _04246_);
  nor (_19624_, _19538_, _04246_);
  or (_19625_, _19624_, _19623_);
  and (_19626_, _19625_, _03823_);
  nor (_19627_, _19557_, _03823_);
  or (_19628_, _19627_, _19626_);
  and (_19629_, _19628_, _03514_);
  and (_19630_, _12794_, _05251_);
  nor (_19631_, _19630_, _19522_);
  nor (_19632_, _19631_, _03514_);
  or (_19634_, _19632_, _19629_);
  or (_19635_, _19634_, _43004_);
  or (_19636_, _43000_, \oc8051_golden_model_1.IP [3]);
  and (_19637_, _19636_, _41806_);
  and (_43530_, _19637_, _19635_);
  not (_19638_, \oc8051_golden_model_1.IP [4]);
  nor (_19639_, _05251_, _19638_);
  nor (_19640_, _05777_, _09129_);
  nor (_19641_, _19640_, _19639_);
  and (_19642_, _19641_, _07390_);
  nor (_19644_, _05908_, _19638_);
  and (_19645_, _12827_, _05908_);
  nor (_19646_, _19645_, _19644_);
  nor (_19647_, _19646_, _03736_);
  and (_19648_, _05251_, \oc8051_golden_model_1.ACC [4]);
  nor (_19649_, _19648_, _19639_);
  nor (_19650_, _19649_, _09029_);
  nor (_19651_, _04409_, _19638_);
  or (_19652_, _19651_, _19650_);
  and (_19653_, _19652_, _04081_);
  nor (_19655_, _12841_, _09129_);
  nor (_19656_, _19655_, _19639_);
  nor (_19657_, _19656_, _04081_);
  or (_19658_, _19657_, _19653_);
  and (_19659_, _19658_, _04055_);
  and (_19660_, _12845_, _05908_);
  nor (_19661_, _19660_, _19644_);
  nor (_19662_, _19661_, _04055_);
  or (_19663_, _19662_, _03723_);
  or (_19664_, _19663_, _19659_);
  nand (_19666_, _19641_, _03723_);
  and (_19667_, _19666_, _19664_);
  and (_19668_, _19667_, _03737_);
  nor (_19669_, _19649_, _03737_);
  or (_19670_, _19669_, _19668_);
  and (_19671_, _19670_, _03736_);
  nor (_19672_, _19671_, _19647_);
  nor (_19673_, _19672_, _03719_);
  nor (_19674_, _19644_, _12860_);
  or (_19675_, _19661_, _06840_);
  nor (_19677_, _19675_, _19674_);
  nor (_19678_, _19677_, _19673_);
  nor (_19679_, _19678_, _03505_);
  nor (_19680_, _12825_, _09166_);
  nor (_19681_, _19680_, _19644_);
  nor (_19682_, _19681_, _03710_);
  nor (_19683_, _19682_, _07390_);
  not (_19684_, _19683_);
  nor (_19685_, _19684_, _19679_);
  nor (_19686_, _19685_, _19642_);
  nor (_19688_, _19686_, _04481_);
  and (_19689_, _06730_, _05251_);
  nor (_19690_, _19639_, _07400_);
  not (_19691_, _19690_);
  nor (_19692_, _19691_, _19689_);
  nor (_19693_, _19692_, _03222_);
  not (_19694_, _19693_);
  nor (_19695_, _19694_, _19688_);
  nor (_19696_, _12933_, _09129_);
  nor (_19697_, _19696_, _19639_);
  nor (_19699_, _19697_, _03589_);
  or (_19700_, _19699_, _08828_);
  or (_19701_, _19700_, _19695_);
  and (_19702_, _12821_, _05251_);
  or (_19703_, _19639_, _07766_);
  or (_19704_, _19703_, _19702_);
  and (_19705_, _06298_, _05251_);
  nor (_19706_, _19705_, _19639_);
  and (_19707_, _19706_, _03601_);
  nor (_19708_, _19707_, _03780_);
  and (_19710_, _19708_, _19704_);
  and (_19711_, _19710_, _19701_);
  and (_19712_, _12817_, _05251_);
  nor (_19713_, _19712_, _19639_);
  nor (_19714_, _19713_, _07778_);
  nor (_19715_, _19714_, _19711_);
  nor (_19716_, _19715_, _03622_);
  nor (_19717_, _19639_, _05825_);
  not (_19718_, _19717_);
  nor (_19719_, _19706_, _07777_);
  and (_19721_, _19719_, _19718_);
  nor (_19722_, _19721_, _19716_);
  nor (_19723_, _19722_, _03790_);
  nor (_19724_, _19649_, _06828_);
  and (_19725_, _19724_, _19718_);
  or (_19726_, _19725_, _19723_);
  and (_19727_, _19726_, _07795_);
  nor (_19728_, _12819_, _09129_);
  nor (_19729_, _19728_, _19639_);
  nor (_19730_, _19729_, _07795_);
  or (_19732_, _19730_, _19727_);
  and (_19733_, _19732_, _07793_);
  nor (_19734_, _12816_, _09129_);
  nor (_19735_, _19734_, _19639_);
  nor (_19736_, _19735_, _07793_);
  or (_19737_, _19736_, _19733_);
  and (_19738_, _19737_, _04246_);
  nor (_19739_, _19656_, _04246_);
  or (_19740_, _19739_, _19738_);
  and (_19741_, _19740_, _03823_);
  nor (_19743_, _19646_, _03823_);
  or (_19744_, _19743_, _19741_);
  and (_19745_, _19744_, _03514_);
  and (_19746_, _13003_, _05251_);
  nor (_19747_, _19746_, _19639_);
  nor (_19748_, _19747_, _03514_);
  or (_19749_, _19748_, _19745_);
  or (_19750_, _19749_, _43004_);
  or (_19751_, _43000_, \oc8051_golden_model_1.IP [4]);
  and (_19752_, _19751_, _41806_);
  and (_43531_, _19752_, _19750_);
  not (_19754_, \oc8051_golden_model_1.IP [5]);
  nor (_19755_, _05251_, _19754_);
  and (_19756_, _06684_, _05251_);
  or (_19757_, _19756_, _19755_);
  and (_19758_, _19757_, _04481_);
  and (_19759_, _05251_, \oc8051_golden_model_1.ACC [5]);
  nor (_19760_, _19759_, _19755_);
  nor (_19761_, _19760_, _09029_);
  nor (_19762_, _04409_, _19754_);
  or (_19764_, _19762_, _19761_);
  and (_19765_, _19764_, _04081_);
  nor (_19766_, _13014_, _09129_);
  nor (_19767_, _19766_, _19755_);
  nor (_19768_, _19767_, _04081_);
  or (_19769_, _19768_, _19765_);
  and (_19770_, _19769_, _04055_);
  nor (_19771_, _05908_, _19754_);
  and (_19772_, _13037_, _05908_);
  nor (_19773_, _19772_, _19771_);
  nor (_19775_, _19773_, _04055_);
  or (_19776_, _19775_, _03723_);
  or (_19777_, _19776_, _19770_);
  nor (_19778_, _05469_, _09129_);
  nor (_19779_, _19778_, _19755_);
  nand (_19780_, _19779_, _03723_);
  and (_19781_, _19780_, _19777_);
  and (_19782_, _19781_, _03737_);
  nor (_19783_, _19760_, _03737_);
  or (_19784_, _19783_, _19782_);
  and (_19786_, _19784_, _03736_);
  and (_19787_, _13047_, _05908_);
  nor (_19788_, _19787_, _19771_);
  nor (_19789_, _19788_, _03736_);
  or (_19790_, _19789_, _19786_);
  and (_19791_, _19790_, _06840_);
  nor (_19792_, _19771_, _13054_);
  nor (_19793_, _19792_, _19773_);
  and (_19794_, _19793_, _03719_);
  or (_19795_, _19794_, _19791_);
  and (_19797_, _19795_, _03710_);
  nor (_19798_, _13020_, _09166_);
  nor (_19799_, _19798_, _19771_);
  nor (_19800_, _19799_, _03710_);
  nor (_19801_, _19800_, _07390_);
  not (_19802_, _19801_);
  nor (_19803_, _19802_, _19797_);
  and (_19804_, _19779_, _07390_);
  or (_19805_, _19804_, _04481_);
  nor (_19806_, _19805_, _19803_);
  or (_19808_, _19806_, _19758_);
  and (_19809_, _19808_, _03589_);
  nor (_19810_, _13127_, _09129_);
  nor (_19811_, _19810_, _19755_);
  nor (_19812_, _19811_, _03589_);
  or (_19813_, _19812_, _08828_);
  or (_19814_, _19813_, _19809_);
  and (_19815_, _13141_, _05251_);
  or (_19816_, _19755_, _07766_);
  or (_19817_, _19816_, _19815_);
  and (_19819_, _06306_, _05251_);
  nor (_19820_, _19819_, _19755_);
  and (_19821_, _19820_, _03601_);
  nor (_19822_, _19821_, _03780_);
  and (_19823_, _19822_, _19817_);
  and (_19824_, _19823_, _19814_);
  and (_19825_, _13147_, _05251_);
  nor (_19826_, _19825_, _19755_);
  nor (_19827_, _19826_, _07778_);
  nor (_19828_, _19827_, _19824_);
  nor (_19830_, _19828_, _03622_);
  nor (_19831_, _19755_, _05518_);
  not (_19832_, _19831_);
  nor (_19833_, _19820_, _07777_);
  and (_19834_, _19833_, _19832_);
  nor (_19835_, _19834_, _19830_);
  nor (_19836_, _19835_, _03790_);
  nor (_19837_, _19760_, _06828_);
  and (_19838_, _19837_, _19832_);
  or (_19839_, _19838_, _19836_);
  and (_19841_, _19839_, _07795_);
  nor (_19842_, _13140_, _09129_);
  nor (_19843_, _19842_, _19755_);
  nor (_19844_, _19843_, _07795_);
  or (_19845_, _19844_, _19841_);
  and (_19846_, _19845_, _07793_);
  nor (_19847_, _13146_, _09129_);
  nor (_19848_, _19847_, _19755_);
  nor (_19849_, _19848_, _07793_);
  or (_19850_, _19849_, _19846_);
  and (_19852_, _19850_, _04246_);
  nor (_19853_, _19767_, _04246_);
  or (_19854_, _19853_, _19852_);
  and (_19855_, _19854_, _03823_);
  nor (_19856_, _19788_, _03823_);
  or (_19857_, _19856_, _19855_);
  and (_19858_, _19857_, _03514_);
  and (_19859_, _13199_, _05251_);
  nor (_19860_, _19859_, _19755_);
  nor (_19861_, _19860_, _03514_);
  or (_19863_, _19861_, _19858_);
  or (_19864_, _19863_, _43004_);
  or (_19865_, _43000_, \oc8051_golden_model_1.IP [5]);
  and (_19866_, _19865_, _41806_);
  and (_43532_, _19866_, _19864_);
  not (_19867_, \oc8051_golden_model_1.IP [6]);
  nor (_19868_, _05251_, _19867_);
  and (_19869_, _06455_, _05251_);
  or (_19870_, _19869_, _19868_);
  and (_19871_, _19870_, _04481_);
  and (_19873_, _05251_, \oc8051_golden_model_1.ACC [6]);
  nor (_19874_, _19873_, _19868_);
  nor (_19875_, _19874_, _09029_);
  nor (_19876_, _04409_, _19867_);
  or (_19877_, _19876_, _19875_);
  and (_19878_, _19877_, _04081_);
  nor (_19879_, _13242_, _09129_);
  nor (_19880_, _19879_, _19868_);
  nor (_19881_, _19880_, _04081_);
  or (_19882_, _19881_, _19878_);
  and (_19884_, _19882_, _04055_);
  nor (_19885_, _05908_, _19867_);
  and (_19886_, _13229_, _05908_);
  nor (_19887_, _19886_, _19885_);
  nor (_19888_, _19887_, _04055_);
  or (_19889_, _19888_, _03723_);
  or (_19890_, _19889_, _19884_);
  nor (_19891_, _05363_, _09129_);
  nor (_19892_, _19891_, _19868_);
  nand (_19893_, _19892_, _03723_);
  and (_19895_, _19893_, _19890_);
  and (_19896_, _19895_, _03737_);
  nor (_19897_, _19874_, _03737_);
  or (_19898_, _19897_, _19896_);
  and (_19899_, _19898_, _03736_);
  and (_19900_, _13253_, _05908_);
  nor (_19901_, _19900_, _19885_);
  nor (_19902_, _19901_, _03736_);
  or (_19903_, _19902_, _03719_);
  or (_19904_, _19903_, _19899_);
  nor (_19906_, _19885_, _13260_);
  nor (_19907_, _19906_, _19887_);
  or (_19908_, _19907_, _06840_);
  and (_19909_, _19908_, _03710_);
  and (_19910_, _19909_, _19904_);
  nor (_19911_, _13226_, _09166_);
  nor (_19912_, _19911_, _19885_);
  nor (_19913_, _19912_, _03710_);
  nor (_19914_, _19913_, _07390_);
  not (_19915_, _19914_);
  nor (_19917_, _19915_, _19910_);
  and (_19918_, _19892_, _07390_);
  or (_19919_, _19918_, _04481_);
  nor (_19920_, _19919_, _19917_);
  or (_19921_, _19920_, _19871_);
  and (_19922_, _19921_, _03589_);
  nor (_19923_, _13332_, _09129_);
  nor (_19924_, _19923_, _19868_);
  nor (_19925_, _19924_, _03589_);
  or (_19926_, _19925_, _08828_);
  or (_19928_, _19926_, _19922_);
  and (_19929_, _13347_, _05251_);
  or (_19930_, _19868_, _07766_);
  or (_19931_, _19930_, _19929_);
  and (_19932_, _13339_, _05251_);
  nor (_19933_, _19932_, _19868_);
  and (_19934_, _19933_, _03601_);
  nor (_19935_, _19934_, _03780_);
  and (_19936_, _19935_, _19931_);
  and (_19937_, _19936_, _19928_);
  and (_19939_, _13353_, _05251_);
  nor (_19940_, _19939_, _19868_);
  nor (_19941_, _19940_, _07778_);
  nor (_19942_, _19941_, _19937_);
  nor (_19943_, _19942_, _03622_);
  nor (_19944_, _19868_, _05412_);
  not (_19945_, _19944_);
  nor (_19946_, _19933_, _07777_);
  and (_19947_, _19946_, _19945_);
  nor (_19948_, _19947_, _19943_);
  nor (_19950_, _19948_, _03790_);
  nor (_19951_, _19874_, _06828_);
  and (_19952_, _19951_, _19945_);
  or (_19953_, _19952_, _19950_);
  and (_19954_, _19953_, _07795_);
  nor (_19955_, _13346_, _09129_);
  nor (_19956_, _19955_, _19868_);
  nor (_19957_, _19956_, _07795_);
  or (_19958_, _19957_, _19954_);
  and (_19959_, _19958_, _07793_);
  nor (_19961_, _13352_, _09129_);
  nor (_19962_, _19961_, _19868_);
  nor (_19963_, _19962_, _07793_);
  or (_19964_, _19963_, _19959_);
  and (_19965_, _19964_, _04246_);
  nor (_19966_, _19880_, _04246_);
  or (_19967_, _19966_, _19965_);
  and (_19968_, _19967_, _03823_);
  nor (_19969_, _19901_, _03823_);
  or (_19970_, _19969_, _19968_);
  and (_19972_, _19970_, _03514_);
  and (_19973_, _13402_, _05251_);
  nor (_19974_, _19973_, _19868_);
  nor (_19975_, _19974_, _03514_);
  or (_19976_, _19975_, _19972_);
  or (_19977_, _19976_, _43004_);
  or (_19978_, _43000_, \oc8051_golden_model_1.IP [6]);
  and (_19979_, _19978_, _41806_);
  and (_43533_, _19979_, _19977_);
  not (_19980_, \oc8051_golden_model_1.P0 [0]);
  nor (_19982_, _43000_, _19980_);
  or (_19983_, _19982_, rst);
  nor (_19984_, _05293_, _19980_);
  and (_19985_, _12128_, _05293_);
  or (_19986_, _19985_, _19984_);
  and (_19987_, _19986_, _03780_);
  and (_19988_, _05293_, _04620_);
  or (_19989_, _19988_, _19984_);
  or (_19990_, _19989_, _06838_);
  nor (_19991_, _05666_, _09236_);
  or (_19993_, _19991_, _19984_);
  and (_19994_, _19993_, _03610_);
  nor (_19995_, _04409_, _19980_);
  and (_19996_, _05293_, \oc8051_golden_model_1.ACC [0]);
  or (_19997_, _19996_, _19984_);
  and (_19998_, _19997_, _04409_);
  or (_19999_, _19998_, _19995_);
  and (_20000_, _19999_, _04081_);
  or (_20001_, _20000_, _03715_);
  or (_20002_, _20001_, _19994_);
  and (_20004_, _12021_, _05209_);
  nor (_20005_, _05209_, _19980_);
  or (_20006_, _20005_, _04055_);
  or (_20007_, _20006_, _20004_);
  and (_20008_, _20007_, _03996_);
  and (_20009_, _20008_, _20002_);
  and (_20010_, _19989_, _03723_);
  or (_20011_, _20010_, _03729_);
  or (_20012_, _20011_, _20009_);
  or (_20013_, _19997_, _03737_);
  and (_20015_, _20013_, _03736_);
  and (_20016_, _20015_, _20012_);
  and (_20017_, _19984_, _03714_);
  or (_20018_, _20017_, _03719_);
  or (_20019_, _20018_, _20016_);
  or (_20020_, _19993_, _06840_);
  and (_20021_, _20020_, _03710_);
  and (_20022_, _20021_, _20019_);
  or (_20023_, _12051_, _12009_);
  and (_20024_, _20023_, _05209_);
  or (_20026_, _20024_, _20005_);
  and (_20027_, _20026_, _03505_);
  or (_20028_, _20027_, _07390_);
  or (_20029_, _20028_, _20022_);
  and (_20030_, _20029_, _19990_);
  or (_20031_, _20030_, _04481_);
  and (_20032_, _06546_, _05293_);
  or (_20033_, _19984_, _07400_);
  or (_20034_, _20033_, _20032_);
  and (_20035_, _20034_, _03589_);
  and (_20037_, _20035_, _20031_);
  and (_20038_, _06340_, \oc8051_golden_model_1.P1 [0]);
  and (_20039_, _06343_, \oc8051_golden_model_1.P0 [0]);
  and (_20040_, _06346_, \oc8051_golden_model_1.P2 [0]);
  and (_20041_, _06348_, \oc8051_golden_model_1.P3 [0]);
  or (_20042_, _20041_, _20040_);
  or (_20043_, _20042_, _20039_);
  nor (_20044_, _20043_, _20038_);
  and (_20045_, _20044_, _12076_);
  and (_20046_, _20045_, _12090_);
  nand (_20048_, _20046_, _12106_);
  or (_20049_, _20048_, _12064_);
  and (_20050_, _20049_, _05293_);
  or (_20051_, _20050_, _19984_);
  and (_20052_, _20051_, _03222_);
  or (_20053_, _20052_, _20037_);
  or (_20054_, _20053_, _08828_);
  and (_20055_, _12124_, _05293_);
  or (_20056_, _19984_, _07766_);
  or (_20057_, _20056_, _20055_);
  and (_20059_, _05293_, _06274_);
  or (_20060_, _20059_, _19984_);
  or (_20061_, _20060_, _05886_);
  and (_20062_, _20061_, _07778_);
  and (_20063_, _20062_, _20057_);
  and (_20064_, _20063_, _20054_);
  or (_20065_, _20064_, _19987_);
  and (_20066_, _20065_, _07777_);
  nand (_20067_, _20060_, _03622_);
  nor (_20068_, _20067_, _19991_);
  or (_20070_, _20068_, _20066_);
  and (_20071_, _20070_, _06828_);
  or (_20072_, _19984_, _05666_);
  and (_20073_, _19997_, _03790_);
  and (_20074_, _20073_, _20072_);
  or (_20075_, _20074_, _03624_);
  or (_20076_, _20075_, _20071_);
  nor (_20077_, _12122_, _09236_);
  or (_20078_, _19984_, _07795_);
  or (_20079_, _20078_, _20077_);
  and (_20081_, _20079_, _07793_);
  and (_20082_, _20081_, _20076_);
  nor (_20083_, _12003_, _09236_);
  or (_20084_, _20083_, _19984_);
  and (_20085_, _20084_, _03785_);
  or (_20086_, _20085_, _03815_);
  or (_20087_, _20086_, _20082_);
  or (_20088_, _19993_, _04246_);
  and (_20089_, _20088_, _03823_);
  and (_20090_, _20089_, _20087_);
  and (_20092_, _19984_, _03453_);
  or (_20093_, _20092_, _03447_);
  or (_20094_, _20093_, _20090_);
  or (_20095_, _19993_, _03514_);
  and (_20096_, _20095_, _43000_);
  and (_20097_, _20096_, _20094_);
  or (_43534_, _20097_, _19983_);
  or (_20098_, _05293_, \oc8051_golden_model_1.P0 [1]);
  and (_20099_, _12213_, _05293_);
  not (_20100_, _20099_);
  and (_20102_, _20100_, _20098_);
  or (_20103_, _20102_, _04081_);
  nand (_20104_, _05293_, _03274_);
  and (_20105_, _20104_, _20098_);
  and (_20106_, _20105_, _04409_);
  not (_20107_, \oc8051_golden_model_1.P0 [1]);
  nor (_20108_, _04409_, _20107_);
  or (_20109_, _20108_, _03610_);
  or (_20110_, _20109_, _20106_);
  and (_20111_, _20110_, _04055_);
  and (_20113_, _20111_, _20103_);
  and (_20114_, _12224_, _05209_);
  nor (_20115_, _05209_, _20107_);
  or (_20116_, _20115_, _03723_);
  or (_20117_, _20116_, _20114_);
  and (_20118_, _20117_, _14265_);
  or (_20119_, _20118_, _20113_);
  nor (_20120_, _05293_, _20107_);
  and (_20121_, _05293_, _06764_);
  or (_20122_, _20121_, _20120_);
  or (_20124_, _20122_, _03996_);
  and (_20125_, _20124_, _20119_);
  or (_20126_, _20125_, _03729_);
  or (_20127_, _20105_, _03737_);
  and (_20128_, _20127_, _03736_);
  and (_20129_, _20128_, _20126_);
  and (_20130_, _12211_, _05209_);
  or (_20131_, _20130_, _20115_);
  and (_20132_, _20131_, _03714_);
  or (_20133_, _20132_, _03719_);
  or (_20135_, _20133_, _20129_);
  and (_20136_, _20114_, _12239_);
  or (_20137_, _20115_, _06840_);
  or (_20138_, _20137_, _20136_);
  and (_20139_, _20138_, _20135_);
  and (_20140_, _20139_, _03710_);
  or (_20141_, _12255_, _12211_);
  and (_20142_, _20141_, _05209_);
  or (_20143_, _20115_, _20142_);
  and (_20144_, _20143_, _03505_);
  or (_20146_, _20144_, _07390_);
  or (_20147_, _20146_, _20140_);
  or (_20148_, _20122_, _06838_);
  and (_20149_, _20148_, _20147_);
  or (_20150_, _20149_, _04481_);
  and (_20151_, _06501_, _05293_);
  or (_20152_, _20120_, _07400_);
  or (_20153_, _20152_, _20151_);
  and (_20154_, _20153_, _03589_);
  and (_20155_, _20154_, _20150_);
  and (_20157_, _06340_, \oc8051_golden_model_1.P1 [1]);
  and (_20158_, _06343_, \oc8051_golden_model_1.P0 [1]);
  and (_20159_, _06346_, \oc8051_golden_model_1.P2 [1]);
  and (_20160_, _06348_, \oc8051_golden_model_1.P3 [1]);
  or (_20161_, _20160_, _20159_);
  or (_20162_, _20161_, _20158_);
  nor (_20163_, _20162_, _20157_);
  and (_20164_, _20163_, _12280_);
  and (_20165_, _20164_, _12294_);
  nand (_20166_, _20165_, _12310_);
  or (_20168_, _20166_, _12268_);
  and (_20169_, _20168_, _05293_);
  or (_20170_, _20169_, _20120_);
  and (_20171_, _20170_, _03222_);
  or (_20172_, _20171_, _20155_);
  and (_20173_, _20172_, _03602_);
  or (_20174_, _12327_, _09236_);
  and (_20175_, _20174_, _03600_);
  nand (_20176_, _05293_, _04303_);
  and (_20177_, _20176_, _03601_);
  or (_20179_, _20177_, _20175_);
  and (_20180_, _20179_, _20098_);
  or (_20181_, _20180_, _20173_);
  and (_20182_, _20181_, _07778_);
  or (_20183_, _12333_, _09236_);
  and (_20184_, _20098_, _03780_);
  and (_20185_, _20184_, _20183_);
  or (_20186_, _20185_, _20182_);
  and (_20187_, _20186_, _07777_);
  or (_20188_, _12207_, _09236_);
  and (_20190_, _20098_, _03622_);
  and (_20191_, _20190_, _20188_);
  or (_20192_, _20191_, _20187_);
  and (_20193_, _20192_, _06828_);
  or (_20194_, _20120_, _05618_);
  and (_20195_, _20105_, _03790_);
  and (_20196_, _20195_, _20194_);
  or (_20197_, _20196_, _20193_);
  and (_20198_, _20197_, _03786_);
  or (_20199_, _20176_, _05618_);
  and (_20201_, _20098_, _03624_);
  and (_20202_, _20201_, _20199_);
  or (_20203_, _20104_, _05618_);
  and (_20204_, _20098_, _03785_);
  and (_20205_, _20204_, _20203_);
  or (_20206_, _20205_, _03815_);
  or (_20207_, _20206_, _20202_);
  or (_20208_, _20207_, _20198_);
  or (_20209_, _20102_, _04246_);
  and (_20210_, _20209_, _03823_);
  and (_20212_, _20210_, _20208_);
  and (_20213_, _20131_, _03453_);
  or (_20214_, _20213_, _03447_);
  or (_20215_, _20214_, _20212_);
  or (_20216_, _20120_, _03514_);
  or (_20217_, _20216_, _20099_);
  and (_20218_, _20217_, _43000_);
  and (_20219_, _20218_, _20215_);
  nor (_20220_, _43000_, _20107_);
  or (_20221_, _20220_, rst);
  or (_43535_, _20221_, _20219_);
  not (_20223_, \oc8051_golden_model_1.P0 [2]);
  nor (_20224_, _05293_, _20223_);
  nor (_20225_, _09236_, _04875_);
  or (_20226_, _20225_, _20224_);
  or (_20227_, _20226_, _06838_);
  and (_20228_, _20226_, _03723_);
  nor (_20229_, _05209_, _20223_);
  and (_20230_, _12411_, _05209_);
  or (_20231_, _20230_, _20229_);
  or (_20233_, _20231_, _04055_);
  nor (_20234_, _12416_, _09236_);
  or (_20235_, _20234_, _20224_);
  and (_20236_, _20235_, _03610_);
  nor (_20237_, _04409_, _20223_);
  and (_20238_, _05293_, \oc8051_golden_model_1.ACC [2]);
  or (_20239_, _20238_, _20224_);
  and (_20240_, _20239_, _04409_);
  or (_20241_, _20240_, _20237_);
  and (_20242_, _20241_, _04081_);
  or (_20244_, _20242_, _03715_);
  or (_20245_, _20244_, _20236_);
  and (_20246_, _20245_, _20233_);
  and (_20247_, _20246_, _03996_);
  or (_20248_, _20247_, _20228_);
  or (_20249_, _20248_, _03729_);
  or (_20250_, _20239_, _03737_);
  and (_20251_, _20250_, _03736_);
  and (_20252_, _20251_, _20249_);
  and (_20253_, _12409_, _05209_);
  or (_20255_, _20253_, _20229_);
  and (_20256_, _20255_, _03714_);
  or (_20257_, _20256_, _03719_);
  or (_20258_, _20257_, _20252_);
  or (_20259_, _20229_, _12443_);
  and (_20260_, _20259_, _20231_);
  or (_20261_, _20260_, _06840_);
  and (_20262_, _20261_, _03710_);
  and (_20263_, _20262_, _20258_);
  or (_20264_, _12460_, _12409_);
  and (_20266_, _20264_, _05209_);
  or (_20267_, _20266_, _20229_);
  and (_20268_, _20267_, _03505_);
  or (_20269_, _20268_, _07390_);
  or (_20270_, _20269_, _20263_);
  and (_20271_, _20270_, _20227_);
  or (_20272_, _20271_, _04481_);
  and (_20273_, _06637_, _05293_);
  or (_20274_, _20224_, _07400_);
  or (_20275_, _20274_, _20273_);
  and (_20277_, _20275_, _03589_);
  and (_20278_, _20277_, _20272_);
  and (_20279_, _06340_, \oc8051_golden_model_1.P1 [2]);
  and (_20280_, _06343_, \oc8051_golden_model_1.P0 [2]);
  and (_20281_, _06346_, \oc8051_golden_model_1.P2 [2]);
  and (_20282_, _06348_, \oc8051_golden_model_1.P3 [2]);
  or (_20283_, _20282_, _20281_);
  or (_20284_, _20283_, _20280_);
  nor (_20285_, _20284_, _20279_);
  and (_20286_, _20285_, _12486_);
  and (_20288_, _20286_, _12496_);
  nand (_20289_, _20288_, _12516_);
  or (_20290_, _20289_, _12474_);
  and (_20291_, _20290_, _05293_);
  or (_20292_, _20224_, _20291_);
  and (_20293_, _20292_, _03222_);
  or (_20294_, _20293_, _20278_);
  or (_20295_, _20294_, _08828_);
  and (_20296_, _12533_, _05293_);
  or (_20297_, _20224_, _07766_);
  or (_20299_, _20297_, _20296_);
  and (_20300_, _05293_, _06332_);
  or (_20301_, _20300_, _20224_);
  or (_20302_, _20301_, _05886_);
  and (_20303_, _20302_, _07778_);
  and (_20304_, _20303_, _20299_);
  and (_20305_, _20304_, _20295_);
  and (_20306_, _12539_, _05293_);
  or (_20307_, _20306_, _20224_);
  and (_20308_, _20307_, _03780_);
  or (_20310_, _20308_, _20305_);
  and (_20311_, _20310_, _07777_);
  or (_20312_, _20224_, _05718_);
  and (_20313_, _20301_, _03622_);
  and (_20314_, _20313_, _20312_);
  or (_20315_, _20314_, _20311_);
  and (_20316_, _20315_, _06828_);
  and (_20317_, _20239_, _03790_);
  and (_20318_, _20317_, _20312_);
  or (_20319_, _20318_, _03624_);
  or (_20321_, _20319_, _20316_);
  nor (_20322_, _12532_, _09236_);
  or (_20323_, _20224_, _07795_);
  or (_20324_, _20323_, _20322_);
  and (_20325_, _20324_, _07793_);
  and (_20326_, _20325_, _20321_);
  nor (_20327_, _12538_, _09236_);
  or (_20328_, _20327_, _20224_);
  and (_20329_, _20328_, _03785_);
  or (_20330_, _20329_, _03815_);
  or (_20332_, _20330_, _20326_);
  or (_20333_, _20235_, _04246_);
  and (_20334_, _20333_, _03823_);
  and (_20335_, _20334_, _20332_);
  and (_20336_, _20255_, _03453_);
  or (_20337_, _20336_, _03447_);
  or (_20338_, _20337_, _20335_);
  and (_20339_, _12592_, _05293_);
  or (_20340_, _20224_, _03514_);
  or (_20341_, _20340_, _20339_);
  and (_20343_, _20341_, _43000_);
  and (_20344_, _20343_, _20338_);
  nor (_20345_, _43000_, _20223_);
  or (_20346_, _20345_, rst);
  or (_43536_, _20346_, _20344_);
  not (_20347_, \oc8051_golden_model_1.P0 [3]);
  nor (_20348_, _43000_, _20347_);
  or (_20349_, _20348_, rst);
  nor (_20350_, _05293_, _20347_);
  nor (_20351_, _09236_, _05005_);
  or (_20353_, _20351_, _20350_);
  or (_20354_, _20353_, _06838_);
  nor (_20355_, _12627_, _09236_);
  or (_20356_, _20355_, _20350_);
  or (_20357_, _20356_, _04081_);
  and (_20358_, _05293_, \oc8051_golden_model_1.ACC [3]);
  or (_20359_, _20358_, _20350_);
  and (_20360_, _20359_, _04409_);
  nor (_20361_, _04409_, _20347_);
  or (_20362_, _20361_, _03610_);
  or (_20364_, _20362_, _20360_);
  and (_20365_, _20364_, _04055_);
  and (_20366_, _20365_, _20357_);
  nor (_20367_, _05209_, _20347_);
  and (_20368_, _12631_, _05209_);
  or (_20369_, _20368_, _20367_);
  and (_20370_, _20369_, _03715_);
  or (_20371_, _20370_, _03723_);
  or (_20372_, _20371_, _20366_);
  or (_20373_, _20353_, _03996_);
  and (_20375_, _20373_, _20372_);
  or (_20376_, _20375_, _03729_);
  or (_20377_, _20359_, _03737_);
  and (_20378_, _20377_, _03736_);
  and (_20379_, _20378_, _20376_);
  and (_20380_, _12641_, _05209_);
  or (_20381_, _20380_, _20367_);
  and (_20382_, _20381_, _03714_);
  or (_20383_, _20382_, _03719_);
  or (_20384_, _20383_, _20379_);
  or (_20386_, _20367_, _12648_);
  and (_20387_, _20386_, _20369_);
  or (_20388_, _20387_, _06840_);
  and (_20389_, _20388_, _03710_);
  and (_20390_, _20389_, _20384_);
  or (_20391_, _12641_, _12610_);
  and (_20392_, _20391_, _05209_);
  or (_20393_, _20392_, _20367_);
  and (_20394_, _20393_, _03505_);
  or (_20395_, _20394_, _07390_);
  or (_20397_, _20395_, _20390_);
  and (_20398_, _20397_, _20354_);
  or (_20399_, _20398_, _04481_);
  and (_20400_, _06592_, _05293_);
  or (_20401_, _20350_, _07400_);
  or (_20402_, _20401_, _20400_);
  and (_20403_, _20402_, _03589_);
  and (_20404_, _20403_, _20399_);
  and (_20405_, _06343_, \oc8051_golden_model_1.P0 [3]);
  and (_20406_, _06340_, \oc8051_golden_model_1.P1 [3]);
  and (_20408_, _06346_, \oc8051_golden_model_1.P2 [3]);
  and (_20409_, _06348_, \oc8051_golden_model_1.P3 [3]);
  or (_20410_, _20409_, _20408_);
  or (_20411_, _20410_, _20406_);
  nor (_20412_, _20411_, _20405_);
  and (_20413_, _20412_, _12713_);
  and (_20414_, _20413_, _12700_);
  nand (_20415_, _20414_, _12693_);
  or (_20416_, _20415_, _12672_);
  and (_20417_, _20416_, _05293_);
  or (_20419_, _20350_, _20417_);
  and (_20420_, _20419_, _03222_);
  or (_20421_, _20420_, _20404_);
  or (_20422_, _20421_, _08828_);
  and (_20423_, _12733_, _05293_);
  or (_20424_, _20350_, _07766_);
  or (_20425_, _20424_, _20423_);
  and (_20426_, _05293_, _06276_);
  or (_20427_, _20426_, _20350_);
  or (_20428_, _20427_, _05886_);
  and (_20430_, _20428_, _07778_);
  and (_20431_, _20430_, _20425_);
  and (_20432_, _20431_, _20422_);
  and (_20433_, _12739_, _05293_);
  or (_20434_, _20433_, _20350_);
  and (_20435_, _20434_, _03780_);
  or (_20436_, _20435_, _20432_);
  and (_20437_, _20436_, _07777_);
  or (_20438_, _20350_, _05567_);
  and (_20439_, _20427_, _03622_);
  and (_20441_, _20439_, _20438_);
  or (_20442_, _20441_, _20437_);
  and (_20443_, _20442_, _06828_);
  and (_20444_, _20359_, _03790_);
  and (_20445_, _20444_, _20438_);
  or (_20446_, _20445_, _03624_);
  or (_20447_, _20446_, _20443_);
  nor (_20448_, _12732_, _09236_);
  or (_20449_, _20350_, _07795_);
  or (_20450_, _20449_, _20448_);
  and (_20452_, _20450_, _07793_);
  and (_20453_, _20452_, _20447_);
  nor (_20454_, _12738_, _09236_);
  or (_20455_, _20454_, _20350_);
  and (_20456_, _20455_, _03785_);
  or (_20457_, _20456_, _03815_);
  or (_20458_, _20457_, _20453_);
  or (_20459_, _20356_, _04246_);
  and (_20460_, _20459_, _03823_);
  and (_20461_, _20460_, _20458_);
  and (_20462_, _20381_, _03453_);
  or (_20463_, _20462_, _03447_);
  or (_20464_, _20463_, _20461_);
  and (_20465_, _12794_, _05293_);
  or (_20466_, _20350_, _03514_);
  or (_20467_, _20466_, _20465_);
  and (_20468_, _20467_, _43000_);
  and (_20469_, _20468_, _20464_);
  or (_43537_, _20469_, _20349_);
  and (_20470_, _09236_, \oc8051_golden_model_1.P0 [4]);
  nor (_20472_, _05777_, _09236_);
  or (_20473_, _20472_, _20470_);
  or (_20474_, _20473_, _06838_);
  not (_20475_, \oc8051_golden_model_1.P0 [4]);
  nor (_20476_, _05209_, _20475_);
  and (_20477_, _12827_, _05209_);
  or (_20478_, _20477_, _20476_);
  and (_20479_, _20478_, _03714_);
  nor (_20480_, _12841_, _09236_);
  or (_20481_, _20480_, _20470_);
  or (_20483_, _20481_, _04081_);
  and (_20484_, _05293_, \oc8051_golden_model_1.ACC [4]);
  or (_20485_, _20484_, _20470_);
  and (_20486_, _20485_, _04409_);
  nor (_20487_, _04409_, _20475_);
  or (_20488_, _20487_, _03610_);
  or (_20489_, _20488_, _20486_);
  and (_20490_, _20489_, _04055_);
  and (_20491_, _20490_, _20483_);
  and (_20492_, _12845_, _05209_);
  or (_20494_, _20492_, _20476_);
  and (_20495_, _20494_, _03715_);
  or (_20496_, _20495_, _03723_);
  or (_20497_, _20496_, _20491_);
  or (_20498_, _20473_, _03996_);
  and (_20499_, _20498_, _20497_);
  or (_20500_, _20499_, _03729_);
  or (_20501_, _20485_, _03737_);
  and (_20502_, _20501_, _03736_);
  and (_20503_, _20502_, _20500_);
  or (_20504_, _20503_, _20479_);
  and (_20505_, _20504_, _06840_);
  and (_20506_, _12861_, _05209_);
  or (_20507_, _20506_, _20476_);
  and (_20508_, _20507_, _03719_);
  or (_20509_, _20508_, _20505_);
  and (_20510_, _20509_, _03710_);
  or (_20511_, _12827_, _12824_);
  and (_20512_, _20511_, _05209_);
  or (_20513_, _20512_, _20476_);
  and (_20515_, _20513_, _03505_);
  or (_20516_, _20515_, _07390_);
  or (_20517_, _20516_, _20510_);
  and (_20518_, _20517_, _20474_);
  or (_20519_, _20518_, _04481_);
  and (_20520_, _06730_, _05293_);
  or (_20521_, _20470_, _07400_);
  or (_20522_, _20521_, _20520_);
  and (_20523_, _20522_, _03589_);
  and (_20524_, _20523_, _20519_);
  and (_20526_, _06343_, \oc8051_golden_model_1.P0 [4]);
  and (_20527_, _06340_, \oc8051_golden_model_1.P1 [4]);
  and (_20528_, _06346_, \oc8051_golden_model_1.P2 [4]);
  and (_20529_, _06348_, \oc8051_golden_model_1.P3 [4]);
  or (_20530_, _20529_, _20528_);
  or (_20531_, _20530_, _20527_);
  nor (_20532_, _20531_, _20526_);
  and (_20533_, _20532_, _12899_);
  and (_20534_, _20533_, _12913_);
  nand (_20535_, _20534_, _12930_);
  or (_20536_, _20535_, _12887_);
  and (_20537_, _20536_, _05293_);
  or (_20538_, _20537_, _20470_);
  and (_20539_, _20538_, _03222_);
  or (_20540_, _20539_, _08828_);
  or (_20541_, _20540_, _20524_);
  and (_20542_, _12821_, _05293_);
  or (_20543_, _20470_, _07766_);
  or (_20544_, _20543_, _20542_);
  and (_20545_, _06298_, _05293_);
  or (_20547_, _20545_, _20470_);
  or (_20548_, _20547_, _05886_);
  and (_20549_, _20548_, _07778_);
  and (_20550_, _20549_, _20544_);
  and (_20551_, _20550_, _20541_);
  and (_20552_, _12817_, _05293_);
  or (_20553_, _20552_, _20470_);
  and (_20554_, _20553_, _03780_);
  or (_20555_, _20554_, _20551_);
  and (_20556_, _20555_, _07777_);
  or (_20558_, _20470_, _05825_);
  and (_20559_, _20547_, _03622_);
  and (_20560_, _20559_, _20558_);
  or (_20561_, _20560_, _20556_);
  and (_20562_, _20561_, _06828_);
  and (_20563_, _20485_, _03790_);
  and (_20564_, _20563_, _20558_);
  or (_20565_, _20564_, _03624_);
  or (_20566_, _20565_, _20562_);
  nor (_20567_, _12819_, _09236_);
  or (_20568_, _20470_, _07795_);
  or (_20569_, _20568_, _20567_);
  and (_20570_, _20569_, _07793_);
  and (_20571_, _20570_, _20566_);
  nor (_20572_, _12816_, _09236_);
  or (_20573_, _20572_, _20470_);
  and (_20574_, _20573_, _03785_);
  or (_20575_, _20574_, _03815_);
  or (_20576_, _20575_, _20571_);
  or (_20577_, _20481_, _04246_);
  and (_20579_, _20577_, _03823_);
  and (_20580_, _20579_, _20576_);
  and (_20581_, _20478_, _03453_);
  or (_20582_, _20581_, _03447_);
  or (_20583_, _20582_, _20580_);
  and (_20584_, _13003_, _05293_);
  or (_20585_, _20470_, _03514_);
  or (_20586_, _20585_, _20584_);
  and (_20587_, _20586_, _43000_);
  and (_20588_, _20587_, _20583_);
  nor (_20590_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_20591_, _20590_, _04794_);
  or (_43538_, _20591_, _20588_);
  not (_20592_, \oc8051_golden_model_1.P0 [5]);
  nor (_20593_, _43000_, _20592_);
  or (_20594_, _20593_, rst);
  nor (_20595_, _05293_, _20592_);
  nor (_20596_, _13014_, _09236_);
  or (_20597_, _20596_, _20595_);
  or (_20598_, _20597_, _04081_);
  and (_20599_, _05293_, \oc8051_golden_model_1.ACC [5]);
  or (_20600_, _20599_, _20595_);
  and (_20601_, _20600_, _04409_);
  nor (_20602_, _04409_, _20592_);
  or (_20603_, _20602_, _03610_);
  or (_20604_, _20603_, _20601_);
  and (_20605_, _20604_, _04055_);
  and (_20606_, _20605_, _20598_);
  nor (_20607_, _05209_, _20592_);
  and (_20608_, _13037_, _05209_);
  or (_20610_, _20608_, _20607_);
  and (_20611_, _20610_, _03715_);
  or (_20612_, _20611_, _03723_);
  or (_20613_, _20612_, _20606_);
  nor (_20614_, _05469_, _09236_);
  or (_20615_, _20614_, _20595_);
  or (_20616_, _20615_, _03996_);
  and (_20617_, _20616_, _20613_);
  or (_20618_, _20617_, _03729_);
  or (_20619_, _20600_, _03737_);
  and (_20621_, _20619_, _03736_);
  and (_20622_, _20621_, _20618_);
  and (_20623_, _13047_, _05209_);
  or (_20624_, _20623_, _20607_);
  and (_20625_, _20624_, _03714_);
  or (_20626_, _20625_, _03719_);
  or (_20627_, _20626_, _20622_);
  or (_20628_, _20607_, _13054_);
  and (_20629_, _20628_, _20610_);
  or (_20630_, _20629_, _06840_);
  and (_20631_, _20630_, _03710_);
  and (_20632_, _20631_, _20627_);
  or (_20633_, _13047_, _13019_);
  and (_20634_, _20633_, _05209_);
  or (_20635_, _20634_, _20607_);
  and (_20636_, _20635_, _03505_);
  or (_20637_, _20636_, _07390_);
  or (_20638_, _20637_, _20632_);
  or (_20639_, _20615_, _06838_);
  and (_20640_, _20639_, _20638_);
  or (_20642_, _20640_, _04481_);
  and (_20643_, _06684_, _05293_);
  or (_20644_, _20595_, _07400_);
  or (_20645_, _20644_, _20643_);
  and (_20646_, _20645_, _03589_);
  and (_20647_, _20646_, _20642_);
  and (_20648_, _06340_, \oc8051_golden_model_1.P1 [5]);
  and (_20649_, _06343_, \oc8051_golden_model_1.P0 [5]);
  and (_20650_, _06346_, \oc8051_golden_model_1.P2 [5]);
  and (_20651_, _06348_, \oc8051_golden_model_1.P3 [5]);
  or (_20653_, _20651_, _20650_);
  or (_20654_, _20653_, _20649_);
  or (_20655_, _20654_, _20648_);
  nor (_20656_, _20655_, _13103_);
  and (_20657_, _20656_, _13122_);
  and (_20658_, _20657_, _13102_);
  nand (_20659_, _20658_, _13095_);
  or (_20660_, _20659_, _13081_);
  and (_20661_, _20660_, _05293_);
  or (_20662_, _20661_, _20595_);
  and (_20663_, _20662_, _03222_);
  or (_20664_, _20663_, _08828_);
  or (_20665_, _20664_, _20647_);
  and (_20666_, _13141_, _05293_);
  or (_20667_, _20595_, _07766_);
  or (_20668_, _20667_, _20666_);
  and (_20669_, _06306_, _05293_);
  or (_20670_, _20669_, _20595_);
  or (_20671_, _20670_, _05886_);
  and (_20672_, _20671_, _07778_);
  and (_20674_, _20672_, _20668_);
  and (_20675_, _20674_, _20665_);
  and (_20676_, _13147_, _05293_);
  or (_20677_, _20676_, _20595_);
  and (_20678_, _20677_, _03780_);
  or (_20679_, _20678_, _20675_);
  and (_20680_, _20679_, _07777_);
  or (_20681_, _20595_, _05518_);
  and (_20682_, _20670_, _03622_);
  and (_20683_, _20682_, _20681_);
  or (_20685_, _20683_, _20680_);
  and (_20686_, _20685_, _06828_);
  and (_20687_, _20600_, _03790_);
  and (_20688_, _20687_, _20681_);
  or (_20689_, _20688_, _03624_);
  or (_20690_, _20689_, _20686_);
  nor (_20691_, _13140_, _09236_);
  or (_20692_, _20595_, _07795_);
  or (_20693_, _20692_, _20691_);
  and (_20694_, _20693_, _07793_);
  and (_20695_, _20694_, _20690_);
  nor (_20696_, _13146_, _09236_);
  or (_20697_, _20696_, _20595_);
  and (_20698_, _20697_, _03785_);
  or (_20699_, _20698_, _03815_);
  or (_20700_, _20699_, _20695_);
  or (_20701_, _20597_, _04246_);
  and (_20702_, _20701_, _03823_);
  and (_20703_, _20702_, _20700_);
  and (_20704_, _20624_, _03453_);
  or (_20706_, _20704_, _03447_);
  or (_20707_, _20706_, _20703_);
  and (_20708_, _13199_, _05293_);
  or (_20709_, _20595_, _03514_);
  or (_20710_, _20709_, _20708_);
  and (_20711_, _20710_, _43000_);
  and (_20712_, _20711_, _20707_);
  or (_43539_, _20712_, _20594_);
  not (_20713_, \oc8051_golden_model_1.P0 [6]);
  nor (_20714_, _05293_, _20713_);
  nor (_20716_, _13242_, _09236_);
  or (_20717_, _20716_, _20714_);
  or (_20718_, _20717_, _04081_);
  and (_20719_, _05293_, \oc8051_golden_model_1.ACC [6]);
  or (_20720_, _20719_, _20714_);
  and (_20721_, _20720_, _04409_);
  nor (_20722_, _04409_, _20713_);
  or (_20723_, _20722_, _03610_);
  or (_20724_, _20723_, _20721_);
  and (_20725_, _20724_, _04055_);
  and (_20726_, _20725_, _20718_);
  nor (_20727_, _05209_, _20713_);
  and (_20728_, _13229_, _05209_);
  or (_20729_, _20728_, _20727_);
  and (_20730_, _20729_, _03715_);
  or (_20731_, _20730_, _03723_);
  or (_20732_, _20731_, _20726_);
  nor (_20733_, _05363_, _09236_);
  or (_20734_, _20733_, _20714_);
  or (_20735_, _20734_, _03996_);
  and (_20737_, _20735_, _20732_);
  or (_20738_, _20737_, _03729_);
  or (_20739_, _20720_, _03737_);
  and (_20740_, _20739_, _03736_);
  and (_20741_, _20740_, _20738_);
  and (_20742_, _13253_, _05209_);
  or (_20743_, _20742_, _20727_);
  and (_20744_, _20743_, _03714_);
  or (_20745_, _20744_, _03719_);
  or (_20746_, _20745_, _20741_);
  or (_20748_, _20727_, _13260_);
  and (_20749_, _20748_, _20729_);
  or (_20750_, _20749_, _06840_);
  and (_20751_, _20750_, _03710_);
  and (_20752_, _20751_, _20746_);
  or (_20753_, _13253_, _13225_);
  and (_20754_, _20753_, _05209_);
  or (_20755_, _20754_, _20727_);
  and (_20756_, _20755_, _03505_);
  or (_20757_, _20756_, _07390_);
  or (_20758_, _20757_, _20752_);
  or (_20759_, _20734_, _06838_);
  and (_20760_, _20759_, _20758_);
  or (_20761_, _20760_, _04481_);
  and (_20762_, _06455_, _05293_);
  or (_20763_, _20714_, _07400_);
  or (_20764_, _20763_, _20762_);
  and (_20765_, _20764_, _03589_);
  and (_20766_, _20765_, _20761_);
  and (_20767_, _06340_, \oc8051_golden_model_1.P1 [6]);
  and (_20769_, _06343_, \oc8051_golden_model_1.P0 [6]);
  and (_20770_, _06346_, \oc8051_golden_model_1.P2 [6]);
  and (_20771_, _06348_, \oc8051_golden_model_1.P3 [6]);
  or (_20772_, _20771_, _20770_);
  or (_20773_, _20772_, _20769_);
  nor (_20774_, _20773_, _20767_);
  and (_20775_, _20774_, _13290_);
  and (_20776_, _20775_, _13313_);
  nand (_20777_, _20776_, _13329_);
  or (_20778_, _20777_, _13287_);
  and (_20780_, _20778_, _05293_);
  or (_20781_, _20780_, _20714_);
  and (_20782_, _20781_, _03222_);
  or (_20783_, _20782_, _08828_);
  or (_20784_, _20783_, _20766_);
  and (_20785_, _13347_, _05293_);
  or (_20786_, _20714_, _07766_);
  or (_20787_, _20786_, _20785_);
  and (_20788_, _13339_, _05293_);
  or (_20789_, _20788_, _20714_);
  or (_20790_, _20789_, _05886_);
  and (_20791_, _20790_, _07778_);
  and (_20792_, _20791_, _20787_);
  and (_20793_, _20792_, _20784_);
  and (_20794_, _13353_, _05293_);
  or (_20795_, _20794_, _20714_);
  and (_20796_, _20795_, _03780_);
  or (_20797_, _20796_, _20793_);
  and (_20798_, _20797_, _07777_);
  or (_20799_, _20714_, _05412_);
  and (_20801_, _20789_, _03622_);
  and (_20802_, _20801_, _20799_);
  or (_20803_, _20802_, _20798_);
  and (_20804_, _20803_, _06828_);
  and (_20805_, _20720_, _03790_);
  and (_20806_, _20805_, _20799_);
  or (_20807_, _20806_, _03624_);
  or (_20808_, _20807_, _20804_);
  nor (_20809_, _13346_, _09236_);
  or (_20810_, _20714_, _07795_);
  or (_20812_, _20810_, _20809_);
  and (_20813_, _20812_, _07793_);
  and (_20814_, _20813_, _20808_);
  nor (_20815_, _13352_, _09236_);
  or (_20816_, _20815_, _20714_);
  and (_20817_, _20816_, _03785_);
  or (_20818_, _20817_, _03815_);
  or (_20819_, _20818_, _20814_);
  or (_20820_, _20717_, _04246_);
  and (_20821_, _20820_, _03823_);
  and (_20822_, _20821_, _20819_);
  and (_20823_, _20743_, _03453_);
  or (_20824_, _20823_, _03447_);
  or (_20825_, _20824_, _20822_);
  and (_20826_, _13402_, _05293_);
  or (_20827_, _20714_, _03514_);
  or (_20828_, _20827_, _20826_);
  and (_20829_, _20828_, _43000_);
  and (_20830_, _20829_, _20825_);
  nor (_20831_, _43000_, _20713_);
  or (_20833_, _20831_, rst);
  or (_43540_, _20833_, _20830_);
  not (_20834_, \oc8051_golden_model_1.P1 [0]);
  nor (_20835_, _43000_, _20834_);
  or (_20836_, _20835_, rst);
  nor (_20837_, _05266_, _20834_);
  and (_20838_, _12128_, _05266_);
  or (_20839_, _20838_, _20837_);
  and (_20840_, _20839_, _03780_);
  and (_20841_, _05266_, _04620_);
  or (_20843_, _20841_, _20837_);
  or (_20844_, _20843_, _06838_);
  nor (_20845_, _05666_, _09352_);
  or (_20846_, _20845_, _20837_);
  and (_20847_, _20846_, _03610_);
  nor (_20848_, _04409_, _20834_);
  and (_20849_, _05266_, \oc8051_golden_model_1.ACC [0]);
  or (_20850_, _20849_, _20837_);
  and (_20851_, _20850_, _04409_);
  or (_20852_, _20851_, _20848_);
  and (_20853_, _20852_, _04081_);
  or (_20854_, _20853_, _03715_);
  or (_20855_, _20854_, _20847_);
  and (_20856_, _12021_, _05916_);
  nor (_20857_, _05916_, _20834_);
  or (_20858_, _20857_, _04055_);
  or (_20859_, _20858_, _20856_);
  and (_20860_, _20859_, _03996_);
  and (_20861_, _20860_, _20855_);
  and (_20862_, _20843_, _03723_);
  or (_20864_, _20862_, _03729_);
  or (_20865_, _20864_, _20861_);
  or (_20866_, _20850_, _03737_);
  and (_20867_, _20866_, _03736_);
  and (_20868_, _20867_, _20865_);
  and (_20869_, _20837_, _03714_);
  or (_20870_, _20869_, _03719_);
  or (_20871_, _20870_, _20868_);
  or (_20872_, _20846_, _06840_);
  and (_20873_, _20872_, _03710_);
  and (_20875_, _20873_, _20871_);
  and (_20876_, _20023_, _05916_);
  or (_20877_, _20876_, _20857_);
  and (_20878_, _20877_, _03505_);
  or (_20879_, _20878_, _07390_);
  or (_20880_, _20879_, _20875_);
  and (_20881_, _20880_, _20844_);
  or (_20882_, _20881_, _04481_);
  and (_20883_, _06546_, _05266_);
  or (_20884_, _20837_, _07400_);
  or (_20886_, _20884_, _20883_);
  and (_20887_, _20886_, _03589_);
  and (_20888_, _20887_, _20882_);
  and (_20889_, _20049_, _05266_);
  or (_20890_, _20889_, _20837_);
  and (_20891_, _20890_, _03222_);
  or (_20892_, _20891_, _20888_);
  or (_20893_, _20892_, _08828_);
  and (_20894_, _12124_, _05266_);
  or (_20895_, _20837_, _07766_);
  or (_20896_, _20895_, _20894_);
  and (_20897_, _05266_, _06274_);
  or (_20898_, _20897_, _20837_);
  or (_20899_, _20898_, _05886_);
  and (_20900_, _20899_, _07778_);
  and (_20901_, _20900_, _20896_);
  and (_20902_, _20901_, _20893_);
  or (_20903_, _20902_, _20840_);
  and (_20904_, _20903_, _07777_);
  nand (_20905_, _20898_, _03622_);
  nor (_20907_, _20905_, _20845_);
  or (_20908_, _20907_, _20904_);
  and (_20909_, _20908_, _06828_);
  or (_20910_, _20837_, _05666_);
  and (_20911_, _20850_, _03790_);
  and (_20912_, _20911_, _20910_);
  or (_20913_, _20912_, _03624_);
  or (_20914_, _20913_, _20909_);
  nor (_20915_, _12122_, _09352_);
  or (_20916_, _20837_, _07795_);
  or (_20918_, _20916_, _20915_);
  and (_20919_, _20918_, _07793_);
  and (_20920_, _20919_, _20914_);
  nor (_20921_, _12003_, _09352_);
  or (_20922_, _20921_, _20837_);
  and (_20923_, _20922_, _03785_);
  or (_20924_, _20923_, _03815_);
  or (_20925_, _20924_, _20920_);
  or (_20926_, _20846_, _04246_);
  and (_20927_, _20926_, _03823_);
  and (_20928_, _20927_, _20925_);
  and (_20929_, _20837_, _03453_);
  or (_20930_, _20929_, _03447_);
  or (_20931_, _20930_, _20928_);
  or (_20932_, _20846_, _03514_);
  and (_20933_, _20932_, _43000_);
  and (_20934_, _20933_, _20931_);
  or (_43543_, _20934_, _20836_);
  or (_20935_, _05266_, \oc8051_golden_model_1.P1 [1]);
  and (_20936_, _12213_, _05266_);
  not (_20938_, _20936_);
  and (_20939_, _20938_, _20935_);
  or (_20940_, _20939_, _04081_);
  nand (_20941_, _05266_, _03274_);
  and (_20942_, _20941_, _20935_);
  and (_20943_, _20942_, _04409_);
  not (_20944_, \oc8051_golden_model_1.P1 [1]);
  nor (_20945_, _04409_, _20944_);
  or (_20946_, _20945_, _03610_);
  or (_20947_, _20946_, _20943_);
  and (_20949_, _20947_, _04055_);
  and (_20950_, _20949_, _20940_);
  and (_20951_, _12224_, _05916_);
  nor (_20952_, _05916_, _20944_);
  or (_20953_, _20952_, _03723_);
  or (_20954_, _20953_, _20951_);
  and (_20955_, _20954_, _14265_);
  or (_20956_, _20955_, _20950_);
  nor (_20957_, _05266_, _20944_);
  and (_20958_, _05266_, _06764_);
  or (_20960_, _20958_, _20957_);
  or (_20961_, _20960_, _03996_);
  and (_20962_, _20961_, _20956_);
  or (_20963_, _20962_, _03729_);
  or (_20964_, _20942_, _03737_);
  and (_20965_, _20964_, _03736_);
  and (_20966_, _20965_, _20963_);
  and (_20967_, _12211_, _05916_);
  or (_20968_, _20967_, _20952_);
  and (_20969_, _20968_, _03714_);
  or (_20970_, _20969_, _03719_);
  or (_20971_, _20970_, _20966_);
  and (_20972_, _20951_, _12239_);
  or (_20973_, _20952_, _06840_);
  or (_20974_, _20973_, _20972_);
  and (_20975_, _20974_, _20971_);
  and (_20976_, _20975_, _03710_);
  and (_20977_, _20141_, _05916_);
  or (_20978_, _20952_, _20977_);
  and (_20979_, _20978_, _03505_);
  or (_20981_, _20979_, _07390_);
  or (_20982_, _20981_, _20976_);
  or (_20983_, _20960_, _06838_);
  and (_20984_, _20983_, _20982_);
  or (_20985_, _20984_, _04481_);
  and (_20986_, _06501_, _05266_);
  or (_20987_, _20957_, _07400_);
  or (_20988_, _20987_, _20986_);
  and (_20989_, _20988_, _03589_);
  and (_20990_, _20989_, _20985_);
  and (_20992_, _20168_, _05266_);
  or (_20993_, _20992_, _20957_);
  and (_20994_, _20993_, _03222_);
  or (_20995_, _20994_, _20990_);
  and (_20996_, _20995_, _03602_);
  or (_20997_, _12327_, _09352_);
  and (_20998_, _20997_, _03600_);
  nand (_20999_, _05266_, _04303_);
  and (_21000_, _20999_, _03601_);
  or (_21001_, _21000_, _20998_);
  and (_21002_, _21001_, _20935_);
  or (_21003_, _21002_, _20996_);
  and (_21004_, _21003_, _07778_);
  or (_21005_, _12333_, _09352_);
  and (_21006_, _20935_, _03780_);
  and (_21007_, _21006_, _21005_);
  or (_21008_, _21007_, _21004_);
  and (_21009_, _21008_, _07777_);
  or (_21010_, _12207_, _09352_);
  and (_21011_, _20935_, _03622_);
  and (_21013_, _21011_, _21010_);
  or (_21014_, _21013_, _21009_);
  and (_21015_, _21014_, _06828_);
  or (_21016_, _20957_, _05618_);
  and (_21017_, _20942_, _03790_);
  and (_21018_, _21017_, _21016_);
  or (_21019_, _21018_, _21015_);
  and (_21020_, _21019_, _03786_);
  or (_21021_, _20999_, _05618_);
  and (_21022_, _20935_, _03624_);
  and (_21024_, _21022_, _21021_);
  or (_21025_, _20941_, _05618_);
  and (_21026_, _20935_, _03785_);
  and (_21027_, _21026_, _21025_);
  or (_21028_, _21027_, _03815_);
  or (_21029_, _21028_, _21024_);
  or (_21030_, _21029_, _21020_);
  or (_21031_, _20939_, _04246_);
  and (_21032_, _21031_, _03823_);
  and (_21033_, _21032_, _21030_);
  and (_21035_, _20968_, _03453_);
  or (_21036_, _21035_, _03447_);
  or (_21037_, _21036_, _21033_);
  or (_21038_, _20957_, _03514_);
  or (_21039_, _21038_, _20936_);
  and (_21040_, _21039_, _43000_);
  and (_21041_, _21040_, _21037_);
  nor (_21042_, _43000_, _20944_);
  or (_21043_, _21042_, rst);
  or (_43544_, _21043_, _21041_);
  not (_21045_, \oc8051_golden_model_1.P1 [2]);
  nor (_21046_, _43000_, _21045_);
  or (_21047_, _21046_, rst);
  nor (_21048_, _05266_, _21045_);
  nor (_21049_, _09352_, _04875_);
  or (_21050_, _21049_, _21048_);
  or (_21051_, _21050_, _06838_);
  or (_21052_, _21050_, _03996_);
  nor (_21053_, _12416_, _09352_);
  or (_21054_, _21053_, _21048_);
  or (_21056_, _21054_, _04081_);
  and (_21057_, _05266_, \oc8051_golden_model_1.ACC [2]);
  or (_21058_, _21057_, _21048_);
  and (_21059_, _21058_, _04409_);
  nor (_21060_, _04409_, _21045_);
  or (_21061_, _21060_, _03610_);
  or (_21062_, _21061_, _21059_);
  and (_21063_, _21062_, _04055_);
  and (_21064_, _21063_, _21056_);
  nor (_21065_, _05916_, _21045_);
  and (_21067_, _12411_, _05916_);
  or (_21068_, _21067_, _21065_);
  and (_21069_, _21068_, _03715_);
  or (_21070_, _21069_, _03723_);
  or (_21071_, _21070_, _21064_);
  and (_21072_, _21071_, _21052_);
  or (_21073_, _21072_, _03729_);
  or (_21074_, _21058_, _03737_);
  and (_21075_, _21074_, _03736_);
  and (_21076_, _21075_, _21073_);
  and (_21078_, _12409_, _05916_);
  or (_21079_, _21078_, _21065_);
  and (_21080_, _21079_, _03714_);
  or (_21081_, _21080_, _03719_);
  or (_21082_, _21081_, _21076_);
  and (_21083_, _21067_, _12443_);
  or (_21084_, _21065_, _06840_);
  or (_21085_, _21084_, _21083_);
  and (_21086_, _21085_, _03710_);
  and (_21087_, _21086_, _21082_);
  and (_21089_, _20264_, _05916_);
  or (_21090_, _21089_, _21065_);
  and (_21091_, _21090_, _03505_);
  or (_21092_, _21091_, _07390_);
  or (_21093_, _21092_, _21087_);
  and (_21094_, _21093_, _21051_);
  or (_21095_, _21094_, _04481_);
  and (_21096_, _06637_, _05266_);
  or (_21097_, _21048_, _07400_);
  or (_21098_, _21097_, _21096_);
  and (_21100_, _21098_, _03589_);
  and (_21101_, _21100_, _21095_);
  and (_21102_, _20290_, _05266_);
  or (_21103_, _21048_, _21102_);
  and (_21104_, _21103_, _03222_);
  or (_21105_, _21104_, _21101_);
  or (_21106_, _21105_, _08828_);
  and (_21107_, _12533_, _05266_);
  or (_21108_, _21048_, _07766_);
  or (_21109_, _21108_, _21107_);
  and (_21110_, _05266_, _06332_);
  or (_21111_, _21110_, _21048_);
  or (_21112_, _21111_, _05886_);
  and (_21113_, _21112_, _07778_);
  and (_21114_, _21113_, _21109_);
  and (_21115_, _21114_, _21106_);
  and (_21116_, _12539_, _05266_);
  or (_21117_, _21116_, _21048_);
  and (_21118_, _21117_, _03780_);
  or (_21119_, _21118_, _21115_);
  and (_21120_, _21119_, _07777_);
  or (_21121_, _21048_, _05718_);
  and (_21122_, _21111_, _03622_);
  and (_21123_, _21122_, _21121_);
  or (_21124_, _21123_, _21120_);
  and (_21125_, _21124_, _06828_);
  and (_21126_, _21058_, _03790_);
  and (_21127_, _21126_, _21121_);
  or (_21128_, _21127_, _03624_);
  or (_21129_, _21128_, _21125_);
  nor (_21131_, _12532_, _09352_);
  or (_21132_, _21048_, _07795_);
  or (_21133_, _21132_, _21131_);
  and (_21134_, _21133_, _07793_);
  and (_21135_, _21134_, _21129_);
  nor (_21136_, _12538_, _09352_);
  or (_21137_, _21136_, _21048_);
  and (_21138_, _21137_, _03785_);
  or (_21139_, _21138_, _03815_);
  or (_21140_, _21139_, _21135_);
  or (_21142_, _21054_, _04246_);
  and (_21143_, _21142_, _03823_);
  and (_21144_, _21143_, _21140_);
  and (_21145_, _21079_, _03453_);
  or (_21146_, _21145_, _03447_);
  or (_21147_, _21146_, _21144_);
  and (_21148_, _12592_, _05266_);
  or (_21149_, _21048_, _03514_);
  or (_21150_, _21149_, _21148_);
  and (_21151_, _21150_, _43000_);
  and (_21153_, _21151_, _21147_);
  or (_43545_, _21153_, _21047_);
  and (_21154_, _09352_, \oc8051_golden_model_1.P1 [3]);
  nor (_21155_, _09352_, _05005_);
  or (_21156_, _21155_, _21154_);
  or (_21157_, _21156_, _06838_);
  nor (_21158_, _12627_, _09352_);
  or (_21159_, _21158_, _21154_);
  or (_21160_, _21159_, _04081_);
  and (_21161_, _05266_, \oc8051_golden_model_1.ACC [3]);
  or (_21163_, _21161_, _21154_);
  and (_21164_, _21163_, _04409_);
  and (_21165_, _09029_, \oc8051_golden_model_1.P1 [3]);
  or (_21166_, _21165_, _03610_);
  or (_21167_, _21166_, _21164_);
  and (_21168_, _21167_, _04055_);
  and (_21169_, _21168_, _21160_);
  not (_21170_, _05916_);
  and (_21171_, _21170_, \oc8051_golden_model_1.P1 [3]);
  and (_21172_, _12631_, _05916_);
  or (_21174_, _21172_, _21171_);
  and (_21175_, _21174_, _03715_);
  or (_21176_, _21175_, _03723_);
  or (_21177_, _21176_, _21169_);
  or (_21178_, _21156_, _03996_);
  and (_21179_, _21178_, _21177_);
  or (_21180_, _21179_, _03729_);
  or (_21181_, _21163_, _03737_);
  and (_21182_, _21181_, _03736_);
  and (_21183_, _21182_, _21180_);
  and (_21185_, _12641_, _05916_);
  or (_21186_, _21185_, _21171_);
  and (_21187_, _21186_, _03714_);
  or (_21188_, _21187_, _03719_);
  or (_21189_, _21188_, _21183_);
  or (_21190_, _21171_, _12648_);
  and (_21191_, _21190_, _21174_);
  or (_21192_, _21191_, _06840_);
  and (_21193_, _21192_, _03710_);
  and (_21194_, _21193_, _21189_);
  and (_21196_, _20391_, _05916_);
  or (_21197_, _21196_, _21171_);
  and (_21198_, _21197_, _03505_);
  or (_21199_, _21198_, _07390_);
  or (_21200_, _21199_, _21194_);
  and (_21201_, _21200_, _21157_);
  or (_21202_, _21201_, _04481_);
  and (_21203_, _06592_, _05266_);
  or (_21204_, _21154_, _07400_);
  or (_21205_, _21204_, _21203_);
  and (_21207_, _21205_, _03589_);
  and (_21208_, _21207_, _21202_);
  and (_21209_, _20416_, _05266_);
  or (_21210_, _21154_, _21209_);
  and (_21211_, _21210_, _03222_);
  or (_21212_, _21211_, _21208_);
  or (_21213_, _21212_, _08828_);
  and (_21214_, _12733_, _05266_);
  or (_21215_, _21154_, _07766_);
  or (_21216_, _21215_, _21214_);
  and (_21218_, _05266_, _06276_);
  or (_21219_, _21218_, _21154_);
  or (_21220_, _21219_, _05886_);
  and (_21221_, _21220_, _07778_);
  and (_21222_, _21221_, _21216_);
  and (_21223_, _21222_, _21213_);
  and (_21224_, _12739_, _05266_);
  or (_21225_, _21224_, _21154_);
  and (_21226_, _21225_, _03780_);
  or (_21227_, _21226_, _21223_);
  and (_21229_, _21227_, _07777_);
  or (_21230_, _21154_, _05567_);
  and (_21231_, _21219_, _03622_);
  and (_21232_, _21231_, _21230_);
  or (_21233_, _21232_, _21229_);
  and (_21234_, _21233_, _06828_);
  and (_21235_, _21163_, _03790_);
  and (_21236_, _21235_, _21230_);
  or (_21237_, _21236_, _03624_);
  or (_21238_, _21237_, _21234_);
  nor (_21240_, _12732_, _09352_);
  or (_21241_, _21154_, _07795_);
  or (_21242_, _21241_, _21240_);
  and (_21243_, _21242_, _07793_);
  and (_21244_, _21243_, _21238_);
  nor (_21245_, _12738_, _09352_);
  or (_21246_, _21245_, _21154_);
  and (_21247_, _21246_, _03785_);
  or (_21248_, _21247_, _03815_);
  or (_21249_, _21248_, _21244_);
  or (_21251_, _21159_, _04246_);
  and (_21252_, _21251_, _03823_);
  and (_21253_, _21252_, _21249_);
  and (_21254_, _21186_, _03453_);
  or (_21255_, _21254_, _03447_);
  or (_21256_, _21255_, _21253_);
  and (_21257_, _12794_, _05266_);
  or (_21258_, _21154_, _03514_);
  or (_21259_, _21258_, _21257_);
  and (_21260_, _21259_, _43000_);
  and (_21262_, _21260_, _21256_);
  nor (_21263_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_21264_, _21263_, _04794_);
  or (_43546_, _21264_, _21262_);
  nor (_21265_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_21266_, _21265_, _04794_);
  and (_21267_, _09352_, \oc8051_golden_model_1.P1 [4]);
  nor (_21268_, _05777_, _09352_);
  or (_21269_, _21268_, _21267_);
  or (_21270_, _21269_, _06838_);
  and (_21272_, _21170_, \oc8051_golden_model_1.P1 [4]);
  and (_21273_, _12827_, _05916_);
  or (_21274_, _21273_, _21272_);
  and (_21275_, _21274_, _03714_);
  nor (_21276_, _12841_, _09352_);
  or (_21277_, _21276_, _21267_);
  or (_21278_, _21277_, _04081_);
  and (_21279_, _05266_, \oc8051_golden_model_1.ACC [4]);
  or (_21280_, _21279_, _21267_);
  and (_21281_, _21280_, _04409_);
  and (_21283_, _09029_, \oc8051_golden_model_1.P1 [4]);
  or (_21284_, _21283_, _03610_);
  or (_21285_, _21284_, _21281_);
  and (_21286_, _21285_, _04055_);
  and (_21287_, _21286_, _21278_);
  and (_21288_, _12845_, _05916_);
  or (_21289_, _21288_, _21272_);
  and (_21290_, _21289_, _03715_);
  or (_21291_, _21290_, _03723_);
  or (_21292_, _21291_, _21287_);
  or (_21294_, _21269_, _03996_);
  and (_21295_, _21294_, _21292_);
  or (_21296_, _21295_, _03729_);
  or (_21297_, _21280_, _03737_);
  and (_21298_, _21297_, _03736_);
  and (_21299_, _21298_, _21296_);
  or (_21300_, _21299_, _21275_);
  and (_21301_, _21300_, _06840_);
  and (_21302_, _12861_, _05916_);
  or (_21303_, _21302_, _21272_);
  and (_21305_, _21303_, _03719_);
  or (_21306_, _21305_, _21301_);
  and (_21307_, _21306_, _03710_);
  and (_21308_, _20511_, _05916_);
  or (_21309_, _21308_, _21272_);
  and (_21310_, _21309_, _03505_);
  or (_21311_, _21310_, _07390_);
  or (_21312_, _21311_, _21307_);
  and (_21313_, _21312_, _21270_);
  or (_21314_, _21313_, _04481_);
  and (_21316_, _06730_, _05266_);
  or (_21317_, _21267_, _07400_);
  or (_21318_, _21317_, _21316_);
  and (_21319_, _21318_, _03589_);
  and (_21320_, _21319_, _21314_);
  and (_21321_, _20536_, _05266_);
  or (_21322_, _21321_, _21267_);
  and (_21323_, _21322_, _03222_);
  or (_21324_, _21323_, _08828_);
  or (_21325_, _21324_, _21320_);
  and (_21327_, _12821_, _05266_);
  or (_21328_, _21267_, _07766_);
  or (_21329_, _21328_, _21327_);
  and (_21330_, _06298_, _05266_);
  or (_21331_, _21330_, _21267_);
  or (_21332_, _21331_, _05886_);
  and (_21333_, _21332_, _07778_);
  and (_21334_, _21333_, _21329_);
  and (_21335_, _21334_, _21325_);
  and (_21336_, _12817_, _05266_);
  or (_21338_, _21336_, _21267_);
  and (_21339_, _21338_, _03780_);
  or (_21340_, _21339_, _21335_);
  and (_21341_, _21340_, _07777_);
  or (_21342_, _21267_, _05825_);
  and (_21343_, _21331_, _03622_);
  and (_21344_, _21343_, _21342_);
  or (_21345_, _21344_, _21341_);
  and (_21346_, _21345_, _06828_);
  and (_21347_, _21280_, _03790_);
  and (_21349_, _21347_, _21342_);
  or (_21350_, _21349_, _03624_);
  or (_21351_, _21350_, _21346_);
  nor (_21352_, _12819_, _09352_);
  or (_21353_, _21267_, _07795_);
  or (_21354_, _21353_, _21352_);
  and (_21355_, _21354_, _07793_);
  and (_21356_, _21355_, _21351_);
  nor (_21357_, _12816_, _09352_);
  or (_21358_, _21357_, _21267_);
  and (_21360_, _21358_, _03785_);
  or (_21361_, _21360_, _03815_);
  or (_21362_, _21361_, _21356_);
  or (_21363_, _21277_, _04246_);
  and (_21364_, _21363_, _03823_);
  and (_21365_, _21364_, _21362_);
  and (_21366_, _21274_, _03453_);
  or (_21367_, _21366_, _03447_);
  or (_21368_, _21367_, _21365_);
  and (_21369_, _13003_, _05266_);
  or (_21371_, _21267_, _03514_);
  or (_21372_, _21371_, _21369_);
  and (_21373_, _21372_, _43000_);
  and (_21374_, _21373_, _21368_);
  or (_43547_, _21374_, _21266_);
  nor (_21375_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_21376_, _21375_, _04794_);
  and (_21377_, _09352_, \oc8051_golden_model_1.P1 [5]);
  nor (_21378_, _13014_, _09352_);
  or (_21379_, _21378_, _21377_);
  or (_21381_, _21379_, _04081_);
  and (_21382_, _05266_, \oc8051_golden_model_1.ACC [5]);
  or (_21383_, _21382_, _21377_);
  and (_21384_, _21383_, _04409_);
  and (_21385_, _09029_, \oc8051_golden_model_1.P1 [5]);
  or (_21386_, _21385_, _03610_);
  or (_21387_, _21386_, _21384_);
  and (_21388_, _21387_, _04055_);
  and (_21389_, _21388_, _21381_);
  and (_21390_, _21170_, \oc8051_golden_model_1.P1 [5]);
  and (_21392_, _13037_, _05916_);
  or (_21393_, _21392_, _21390_);
  and (_21394_, _21393_, _03715_);
  or (_21395_, _21394_, _03723_);
  or (_21396_, _21395_, _21389_);
  nor (_21397_, _05469_, _09352_);
  or (_21398_, _21397_, _21377_);
  or (_21399_, _21398_, _03996_);
  and (_21400_, _21399_, _21396_);
  or (_21401_, _21400_, _03729_);
  or (_21403_, _21383_, _03737_);
  and (_21404_, _21403_, _03736_);
  and (_21405_, _21404_, _21401_);
  and (_21406_, _13047_, _05916_);
  or (_21407_, _21406_, _21390_);
  and (_21408_, _21407_, _03714_);
  or (_21409_, _21408_, _03719_);
  or (_21410_, _21409_, _21405_);
  or (_21411_, _21390_, _13054_);
  and (_21412_, _21411_, _21393_);
  or (_21414_, _21412_, _06840_);
  and (_21415_, _21414_, _03710_);
  and (_21416_, _21415_, _21410_);
  and (_21417_, _20633_, _05916_);
  or (_21418_, _21417_, _21390_);
  and (_21419_, _21418_, _03505_);
  or (_21420_, _21419_, _07390_);
  or (_21421_, _21420_, _21416_);
  or (_21422_, _21398_, _06838_);
  and (_21423_, _21422_, _21421_);
  or (_21425_, _21423_, _04481_);
  and (_21426_, _06684_, _05266_);
  or (_21427_, _21377_, _07400_);
  or (_21428_, _21427_, _21426_);
  and (_21429_, _21428_, _03589_);
  and (_21430_, _21429_, _21425_);
  and (_21431_, _20660_, _05266_);
  or (_21432_, _21431_, _21377_);
  and (_21433_, _21432_, _03222_);
  or (_21434_, _21433_, _08828_);
  or (_21436_, _21434_, _21430_);
  and (_21437_, _13141_, _05266_);
  or (_21438_, _21377_, _07766_);
  or (_21439_, _21438_, _21437_);
  and (_21440_, _06306_, _05266_);
  or (_21441_, _21440_, _21377_);
  or (_21442_, _21441_, _05886_);
  and (_21443_, _21442_, _07778_);
  and (_21444_, _21443_, _21439_);
  and (_21445_, _21444_, _21436_);
  and (_21447_, _13147_, _05266_);
  or (_21448_, _21447_, _21377_);
  and (_21449_, _21448_, _03780_);
  or (_21450_, _21449_, _21445_);
  and (_21451_, _21450_, _07777_);
  or (_21452_, _21377_, _05518_);
  and (_21453_, _21441_, _03622_);
  and (_21454_, _21453_, _21452_);
  or (_21455_, _21454_, _21451_);
  and (_21456_, _21455_, _06828_);
  and (_21458_, _21383_, _03790_);
  and (_21459_, _21458_, _21452_);
  or (_21460_, _21459_, _03624_);
  or (_21461_, _21460_, _21456_);
  nor (_21462_, _13140_, _09352_);
  or (_21463_, _21377_, _07795_);
  or (_21464_, _21463_, _21462_);
  and (_21465_, _21464_, _07793_);
  and (_21466_, _21465_, _21461_);
  nor (_21467_, _13146_, _09352_);
  or (_21469_, _21467_, _21377_);
  and (_21470_, _21469_, _03785_);
  or (_21471_, _21470_, _03815_);
  or (_21472_, _21471_, _21466_);
  or (_21473_, _21379_, _04246_);
  and (_21474_, _21473_, _03823_);
  and (_21475_, _21474_, _21472_);
  and (_21476_, _21407_, _03453_);
  or (_21477_, _21476_, _03447_);
  or (_21478_, _21477_, _21475_);
  and (_21480_, _13199_, _05266_);
  or (_21481_, _21377_, _03514_);
  or (_21482_, _21481_, _21480_);
  and (_21483_, _21482_, _43000_);
  and (_21484_, _21483_, _21478_);
  or (_43550_, _21484_, _21376_);
  not (_21485_, \oc8051_golden_model_1.P1 [6]);
  nor (_21486_, _05266_, _21485_);
  nor (_21487_, _13242_, _09352_);
  or (_21488_, _21487_, _21486_);
  or (_21491_, _21488_, _04081_);
  and (_21492_, _05266_, \oc8051_golden_model_1.ACC [6]);
  or (_21493_, _21492_, _21486_);
  and (_21494_, _21493_, _04409_);
  nor (_21495_, _04409_, _21485_);
  or (_21496_, _21495_, _03610_);
  or (_21497_, _21496_, _21494_);
  and (_21498_, _21497_, _04055_);
  and (_21499_, _21498_, _21491_);
  nor (_21500_, _05916_, _21485_);
  and (_21503_, _13229_, _05916_);
  or (_21504_, _21503_, _21500_);
  and (_21505_, _21504_, _03715_);
  or (_21506_, _21505_, _03723_);
  or (_21507_, _21506_, _21499_);
  nor (_21508_, _05363_, _09352_);
  or (_21509_, _21508_, _21486_);
  or (_21510_, _21509_, _03996_);
  and (_21511_, _21510_, _21507_);
  or (_21512_, _21511_, _03729_);
  or (_21515_, _21493_, _03737_);
  and (_21516_, _21515_, _03736_);
  and (_21517_, _21516_, _21512_);
  and (_21518_, _13253_, _05916_);
  or (_21519_, _21518_, _21500_);
  and (_21520_, _21519_, _03714_);
  or (_21521_, _21520_, _03719_);
  or (_21522_, _21521_, _21517_);
  or (_21523_, _21500_, _13260_);
  and (_21524_, _21523_, _21504_);
  or (_21527_, _21524_, _06840_);
  and (_21528_, _21527_, _03710_);
  and (_21529_, _21528_, _21522_);
  and (_21530_, _20753_, _05916_);
  or (_21531_, _21530_, _21500_);
  and (_21532_, _21531_, _03505_);
  or (_21533_, _21532_, _07390_);
  or (_21534_, _21533_, _21529_);
  or (_21535_, _21509_, _06838_);
  and (_21536_, _21535_, _21534_);
  or (_21539_, _21536_, _04481_);
  and (_21540_, _06455_, _05266_);
  or (_21541_, _21486_, _07400_);
  or (_21542_, _21541_, _21540_);
  and (_21543_, _21542_, _03589_);
  and (_21544_, _21543_, _21539_);
  and (_21545_, _20778_, _05266_);
  or (_21546_, _21545_, _21486_);
  and (_21547_, _21546_, _03222_);
  or (_21548_, _21547_, _08828_);
  or (_21551_, _21548_, _21544_);
  and (_21552_, _13347_, _05266_);
  or (_21553_, _21486_, _07766_);
  or (_21554_, _21553_, _21552_);
  and (_21555_, _13339_, _05266_);
  or (_21556_, _21555_, _21486_);
  or (_21557_, _21556_, _05886_);
  and (_21558_, _21557_, _07778_);
  and (_21559_, _21558_, _21554_);
  and (_21560_, _21559_, _21551_);
  and (_21562_, _13353_, _05266_);
  or (_21563_, _21562_, _21486_);
  and (_21564_, _21563_, _03780_);
  or (_21565_, _21564_, _21560_);
  and (_21566_, _21565_, _07777_);
  or (_21567_, _21486_, _05412_);
  and (_21568_, _21556_, _03622_);
  and (_21569_, _21568_, _21567_);
  or (_21570_, _21569_, _21566_);
  and (_21571_, _21570_, _06828_);
  and (_21573_, _21493_, _03790_);
  and (_21574_, _21573_, _21567_);
  or (_21575_, _21574_, _03624_);
  or (_21576_, _21575_, _21571_);
  nor (_21577_, _13346_, _09352_);
  or (_21578_, _21486_, _07795_);
  or (_21579_, _21578_, _21577_);
  and (_21580_, _21579_, _07793_);
  and (_21581_, _21580_, _21576_);
  nor (_21582_, _13352_, _09352_);
  or (_21584_, _21582_, _21486_);
  and (_21585_, _21584_, _03785_);
  or (_21586_, _21585_, _03815_);
  or (_21587_, _21586_, _21581_);
  or (_21588_, _21488_, _04246_);
  and (_21589_, _21588_, _03823_);
  and (_21590_, _21589_, _21587_);
  and (_21591_, _21519_, _03453_);
  or (_21592_, _21591_, _03447_);
  or (_21593_, _21592_, _21590_);
  and (_21595_, _13402_, _05266_);
  or (_21596_, _21486_, _03514_);
  or (_21597_, _21596_, _21595_);
  and (_21598_, _21597_, _43000_);
  and (_21599_, _21598_, _21593_);
  nor (_21600_, _43000_, _21485_);
  or (_21601_, _21600_, rst);
  or (_43551_, _21601_, _21599_);
  not (_21602_, \oc8051_golden_model_1.P2 [0]);
  nor (_21603_, _43000_, _21602_);
  or (_21605_, _21603_, rst);
  nor (_21606_, _05235_, _21602_);
  and (_21607_, _12128_, _05235_);
  or (_21608_, _21607_, _21606_);
  and (_21609_, _21608_, _03780_);
  and (_21610_, _05235_, _04620_);
  or (_21611_, _21610_, _21606_);
  or (_21612_, _21611_, _06838_);
  nor (_21613_, _05666_, _09454_);
  or (_21614_, _21613_, _21606_);
  and (_21616_, _21614_, _03610_);
  nor (_21617_, _04409_, _21602_);
  and (_21618_, _05235_, \oc8051_golden_model_1.ACC [0]);
  or (_21619_, _21618_, _21606_);
  and (_21620_, _21619_, _04409_);
  or (_21621_, _21620_, _21617_);
  and (_21622_, _21621_, _04081_);
  or (_21623_, _21622_, _03715_);
  or (_21624_, _21623_, _21616_);
  and (_21625_, _12021_, _05918_);
  nor (_21627_, _05918_, _21602_);
  or (_21628_, _21627_, _04055_);
  or (_21629_, _21628_, _21625_);
  and (_21630_, _21629_, _03996_);
  and (_21631_, _21630_, _21624_);
  and (_21632_, _21611_, _03723_);
  or (_21633_, _21632_, _03729_);
  or (_21634_, _21633_, _21631_);
  or (_21635_, _21619_, _03737_);
  and (_21636_, _21635_, _03736_);
  and (_21638_, _21636_, _21634_);
  and (_21639_, _21606_, _03714_);
  or (_21640_, _21639_, _03719_);
  or (_21641_, _21640_, _21638_);
  or (_21642_, _21614_, _06840_);
  and (_21643_, _21642_, _03710_);
  and (_21644_, _21643_, _21641_);
  and (_21645_, _20023_, _05918_);
  or (_21646_, _21645_, _21627_);
  and (_21647_, _21646_, _03505_);
  or (_21649_, _21647_, _07390_);
  or (_21650_, _21649_, _21644_);
  and (_21651_, _21650_, _21612_);
  or (_21652_, _21651_, _04481_);
  and (_21653_, _06546_, _05235_);
  or (_21654_, _21606_, _07400_);
  or (_21655_, _21654_, _21653_);
  and (_21656_, _21655_, _03589_);
  and (_21657_, _21656_, _21652_);
  and (_21658_, _20049_, _05235_);
  or (_21660_, _21658_, _21606_);
  and (_21661_, _21660_, _03222_);
  or (_21662_, _21661_, _21657_);
  or (_21663_, _21662_, _08828_);
  and (_21664_, _12124_, _05235_);
  or (_21665_, _21606_, _07766_);
  or (_21666_, _21665_, _21664_);
  and (_21667_, _05235_, _06274_);
  or (_21668_, _21667_, _21606_);
  or (_21669_, _21668_, _05886_);
  and (_21671_, _21669_, _07778_);
  and (_21672_, _21671_, _21666_);
  and (_21673_, _21672_, _21663_);
  or (_21674_, _21673_, _21609_);
  and (_21675_, _21674_, _07777_);
  nand (_21676_, _21668_, _03622_);
  nor (_21677_, _21676_, _21613_);
  or (_21678_, _21677_, _21675_);
  and (_21679_, _21678_, _06828_);
  or (_21680_, _21606_, _05666_);
  and (_21682_, _21619_, _03790_);
  and (_21683_, _21682_, _21680_);
  or (_21684_, _21683_, _03624_);
  or (_21685_, _21684_, _21679_);
  nor (_21686_, _12122_, _09454_);
  or (_21687_, _21606_, _07795_);
  or (_21688_, _21687_, _21686_);
  and (_21689_, _21688_, _07793_);
  and (_21690_, _21689_, _21685_);
  nor (_21691_, _12003_, _09454_);
  or (_21693_, _21691_, _21606_);
  and (_21694_, _21693_, _03785_);
  or (_21695_, _21694_, _03815_);
  or (_21696_, _21695_, _21690_);
  or (_21697_, _21614_, _04246_);
  and (_21698_, _21697_, _03823_);
  and (_21699_, _21698_, _21696_);
  and (_21700_, _21606_, _03453_);
  or (_21701_, _21700_, _03447_);
  or (_21702_, _21701_, _21699_);
  or (_21704_, _21614_, _03514_);
  and (_21705_, _21704_, _43000_);
  and (_21706_, _21705_, _21702_);
  or (_43552_, _21706_, _21605_);
  or (_21707_, _05235_, \oc8051_golden_model_1.P2 [1]);
  and (_21708_, _12213_, _05235_);
  not (_21709_, _21708_);
  and (_21710_, _21709_, _21707_);
  or (_21711_, _21710_, _04081_);
  nand (_21712_, _05235_, _03274_);
  and (_21714_, _21712_, _21707_);
  and (_21715_, _21714_, _04409_);
  not (_21716_, \oc8051_golden_model_1.P2 [1]);
  nor (_21717_, _04409_, _21716_);
  or (_21718_, _21717_, _03610_);
  or (_21719_, _21718_, _21715_);
  and (_21720_, _21719_, _04055_);
  and (_21721_, _21720_, _21711_);
  and (_21722_, _12224_, _05918_);
  nor (_21723_, _05918_, _21716_);
  or (_21725_, _21723_, _03723_);
  or (_21726_, _21725_, _21722_);
  and (_21727_, _21726_, _14265_);
  or (_21728_, _21727_, _21721_);
  nor (_21729_, _05235_, _21716_);
  and (_21730_, _05235_, _06764_);
  or (_21731_, _21730_, _21729_);
  or (_21732_, _21731_, _03996_);
  and (_21733_, _21732_, _21728_);
  or (_21734_, _21733_, _03729_);
  or (_21736_, _21714_, _03737_);
  and (_21737_, _21736_, _03736_);
  and (_21738_, _21737_, _21734_);
  and (_21739_, _12211_, _05918_);
  or (_21740_, _21739_, _21723_);
  and (_21741_, _21740_, _03714_);
  or (_21742_, _21741_, _03719_);
  or (_21743_, _21742_, _21738_);
  and (_21744_, _21722_, _12239_);
  or (_21745_, _21723_, _06840_);
  or (_21747_, _21745_, _21744_);
  and (_21748_, _21747_, _21743_);
  and (_21749_, _21748_, _03710_);
  and (_21750_, _20141_, _05918_);
  or (_21751_, _21723_, _21750_);
  and (_21752_, _21751_, _03505_);
  or (_21753_, _21752_, _07390_);
  or (_21754_, _21753_, _21749_);
  or (_21755_, _21731_, _06838_);
  and (_21756_, _21755_, _21754_);
  or (_21758_, _21756_, _04481_);
  and (_21759_, _06501_, _05235_);
  or (_21760_, _21729_, _07400_);
  or (_21761_, _21760_, _21759_);
  and (_21762_, _21761_, _03589_);
  and (_21763_, _21762_, _21758_);
  and (_21764_, _20168_, _05235_);
  or (_21765_, _21764_, _21729_);
  and (_21766_, _21765_, _03222_);
  or (_21767_, _21766_, _21763_);
  and (_21769_, _21767_, _03602_);
  or (_21770_, _12327_, _09454_);
  and (_21771_, _21770_, _03600_);
  nand (_21772_, _05235_, _04303_);
  and (_21773_, _21772_, _03601_);
  or (_21774_, _21773_, _21771_);
  and (_21775_, _21774_, _21707_);
  or (_21776_, _21775_, _21769_);
  and (_21777_, _21776_, _07778_);
  or (_21778_, _12333_, _09454_);
  and (_21780_, _21707_, _03780_);
  and (_21781_, _21780_, _21778_);
  or (_21782_, _21781_, _21777_);
  and (_21783_, _21782_, _07777_);
  or (_21784_, _12207_, _09454_);
  and (_21785_, _21707_, _03622_);
  and (_21786_, _21785_, _21784_);
  or (_21787_, _21786_, _21783_);
  and (_21788_, _21787_, _06828_);
  or (_21789_, _21729_, _05618_);
  and (_21791_, _21714_, _03790_);
  and (_21792_, _21791_, _21789_);
  or (_21793_, _21792_, _21788_);
  and (_21794_, _21793_, _03786_);
  or (_21795_, _21772_, _05618_);
  and (_21796_, _21707_, _03624_);
  and (_21797_, _21796_, _21795_);
  or (_21798_, _21712_, _05618_);
  and (_21799_, _21707_, _03785_);
  and (_21800_, _21799_, _21798_);
  or (_21802_, _21800_, _03815_);
  or (_21803_, _21802_, _21797_);
  or (_21804_, _21803_, _21794_);
  or (_21805_, _21710_, _04246_);
  and (_21806_, _21805_, _03823_);
  and (_21807_, _21806_, _21804_);
  and (_21808_, _21740_, _03453_);
  or (_21809_, _21808_, _03447_);
  or (_21810_, _21809_, _21807_);
  or (_21811_, _21729_, _03514_);
  or (_21813_, _21811_, _21708_);
  and (_21814_, _21813_, _43000_);
  and (_21815_, _21814_, _21810_);
  nor (_21816_, _43000_, _21716_);
  or (_21817_, _21816_, rst);
  or (_43553_, _21817_, _21815_);
  not (_21818_, \oc8051_golden_model_1.P2 [2]);
  nor (_21819_, _43000_, _21818_);
  or (_21820_, _21819_, rst);
  nor (_21821_, _05235_, _21818_);
  nor (_21823_, _09454_, _04875_);
  or (_21824_, _21823_, _21821_);
  or (_21825_, _21824_, _06838_);
  or (_21826_, _21824_, _03996_);
  nor (_21827_, _12416_, _09454_);
  or (_21828_, _21827_, _21821_);
  or (_21829_, _21828_, _04081_);
  and (_21830_, _05235_, \oc8051_golden_model_1.ACC [2]);
  or (_21831_, _21830_, _21821_);
  and (_21832_, _21831_, _04409_);
  nor (_21834_, _04409_, _21818_);
  or (_21835_, _21834_, _03610_);
  or (_21836_, _21835_, _21832_);
  and (_21837_, _21836_, _04055_);
  and (_21838_, _21837_, _21829_);
  nor (_21839_, _05918_, _21818_);
  and (_21840_, _12411_, _05918_);
  or (_21841_, _21840_, _21839_);
  and (_21842_, _21841_, _03715_);
  or (_21843_, _21842_, _03723_);
  or (_21845_, _21843_, _21838_);
  and (_21846_, _21845_, _21826_);
  or (_21847_, _21846_, _03729_);
  or (_21848_, _21831_, _03737_);
  and (_21849_, _21848_, _03736_);
  and (_21850_, _21849_, _21847_);
  and (_21851_, _12409_, _05918_);
  or (_21852_, _21851_, _21839_);
  and (_21853_, _21852_, _03714_);
  or (_21854_, _21853_, _03719_);
  or (_21856_, _21854_, _21850_);
  and (_21857_, _21840_, _12443_);
  or (_21858_, _21839_, _06840_);
  or (_21859_, _21858_, _21857_);
  and (_21860_, _21859_, _03710_);
  and (_21861_, _21860_, _21856_);
  and (_21862_, _20264_, _05918_);
  or (_21863_, _21862_, _21839_);
  and (_21864_, _21863_, _03505_);
  or (_21865_, _21864_, _07390_);
  or (_21867_, _21865_, _21861_);
  and (_21868_, _21867_, _21825_);
  or (_21869_, _21868_, _04481_);
  and (_21870_, _06637_, _05235_);
  or (_21871_, _21821_, _07400_);
  or (_21872_, _21871_, _21870_);
  and (_21873_, _21872_, _03589_);
  and (_21874_, _21873_, _21869_);
  and (_21875_, _20290_, _05235_);
  or (_21876_, _21821_, _21875_);
  and (_21878_, _21876_, _03222_);
  or (_21879_, _21878_, _21874_);
  or (_21880_, _21879_, _08828_);
  and (_21881_, _12533_, _05235_);
  or (_21882_, _21821_, _07766_);
  or (_21883_, _21882_, _21881_);
  and (_21884_, _05235_, _06332_);
  or (_21885_, _21884_, _21821_);
  or (_21886_, _21885_, _05886_);
  and (_21887_, _21886_, _07778_);
  and (_21889_, _21887_, _21883_);
  and (_21890_, _21889_, _21880_);
  and (_21891_, _12539_, _05235_);
  or (_21892_, _21891_, _21821_);
  and (_21893_, _21892_, _03780_);
  or (_21894_, _21893_, _21890_);
  and (_21895_, _21894_, _07777_);
  or (_21896_, _21821_, _05718_);
  and (_21897_, _21885_, _03622_);
  and (_21898_, _21897_, _21896_);
  or (_21900_, _21898_, _21895_);
  and (_21901_, _21900_, _06828_);
  and (_21902_, _21831_, _03790_);
  and (_21903_, _21902_, _21896_);
  or (_21904_, _21903_, _03624_);
  or (_21905_, _21904_, _21901_);
  nor (_21906_, _12532_, _09454_);
  or (_21907_, _21821_, _07795_);
  or (_21908_, _21907_, _21906_);
  and (_21909_, _21908_, _07793_);
  and (_21911_, _21909_, _21905_);
  nor (_21912_, _12538_, _09454_);
  or (_21913_, _21912_, _21821_);
  and (_21914_, _21913_, _03785_);
  or (_21915_, _21914_, _03815_);
  or (_21916_, _21915_, _21911_);
  or (_21917_, _21828_, _04246_);
  and (_21918_, _21917_, _03823_);
  and (_21919_, _21918_, _21916_);
  and (_21920_, _21852_, _03453_);
  or (_21922_, _21920_, _03447_);
  or (_21923_, _21922_, _21919_);
  and (_21924_, _12592_, _05235_);
  or (_21925_, _21821_, _03514_);
  or (_21926_, _21925_, _21924_);
  and (_21927_, _21926_, _43000_);
  and (_21928_, _21927_, _21923_);
  or (_43554_, _21928_, _21820_);
  and (_21929_, _09454_, \oc8051_golden_model_1.P2 [3]);
  nor (_21930_, _09454_, _05005_);
  or (_21932_, _21930_, _21929_);
  or (_21933_, _21932_, _06838_);
  nor (_21934_, _12627_, _09454_);
  or (_21935_, _21934_, _21929_);
  or (_21936_, _21935_, _04081_);
  and (_21937_, _05235_, \oc8051_golden_model_1.ACC [3]);
  or (_21938_, _21937_, _21929_);
  and (_21939_, _21938_, _04409_);
  and (_21940_, _09029_, \oc8051_golden_model_1.P2 [3]);
  or (_21941_, _21940_, _03610_);
  or (_21943_, _21941_, _21939_);
  and (_21944_, _21943_, _04055_);
  and (_21945_, _21944_, _21936_);
  not (_21946_, _05918_);
  and (_21947_, _21946_, \oc8051_golden_model_1.P2 [3]);
  and (_21948_, _12631_, _05918_);
  or (_21949_, _21948_, _21947_);
  and (_21950_, _21949_, _03715_);
  or (_21951_, _21950_, _03723_);
  or (_21952_, _21951_, _21945_);
  or (_21954_, _21932_, _03996_);
  and (_21955_, _21954_, _21952_);
  or (_21956_, _21955_, _03729_);
  or (_21957_, _21938_, _03737_);
  and (_21958_, _21957_, _03736_);
  and (_21959_, _21958_, _21956_);
  and (_21960_, _12641_, _05918_);
  or (_21961_, _21960_, _21947_);
  and (_21962_, _21961_, _03714_);
  or (_21963_, _21962_, _03719_);
  or (_21965_, _21963_, _21959_);
  or (_21966_, _21947_, _12648_);
  and (_21967_, _21966_, _21949_);
  or (_21968_, _21967_, _06840_);
  and (_21969_, _21968_, _03710_);
  and (_21970_, _21969_, _21965_);
  and (_21971_, _20391_, _05918_);
  or (_21972_, _21971_, _21947_);
  and (_21973_, _21972_, _03505_);
  or (_21974_, _21973_, _07390_);
  or (_21976_, _21974_, _21970_);
  and (_21977_, _21976_, _21933_);
  or (_21978_, _21977_, _04481_);
  and (_21979_, _06592_, _05235_);
  or (_21980_, _21929_, _07400_);
  or (_21981_, _21980_, _21979_);
  and (_21982_, _21981_, _03589_);
  and (_21983_, _21982_, _21978_);
  and (_21984_, _20416_, _05235_);
  or (_21985_, _21929_, _21984_);
  and (_21987_, _21985_, _03222_);
  or (_21988_, _21987_, _21983_);
  or (_21989_, _21988_, _08828_);
  and (_21990_, _12733_, _05235_);
  or (_21991_, _21929_, _07766_);
  or (_21992_, _21991_, _21990_);
  and (_21993_, _05235_, _06276_);
  or (_21994_, _21993_, _21929_);
  or (_21995_, _21994_, _05886_);
  and (_21996_, _21995_, _07778_);
  and (_21998_, _21996_, _21992_);
  and (_21999_, _21998_, _21989_);
  and (_22000_, _12739_, _05235_);
  or (_22001_, _22000_, _21929_);
  and (_22002_, _22001_, _03780_);
  or (_22003_, _22002_, _21999_);
  and (_22004_, _22003_, _07777_);
  or (_22005_, _21929_, _05567_);
  and (_22006_, _21994_, _03622_);
  and (_22007_, _22006_, _22005_);
  or (_22009_, _22007_, _22004_);
  and (_22010_, _22009_, _06828_);
  and (_22011_, _21938_, _03790_);
  and (_22012_, _22011_, _22005_);
  or (_22013_, _22012_, _03624_);
  or (_22014_, _22013_, _22010_);
  nor (_22015_, _12732_, _09454_);
  or (_22016_, _21929_, _07795_);
  or (_22017_, _22016_, _22015_);
  and (_22018_, _22017_, _07793_);
  and (_22020_, _22018_, _22014_);
  nor (_22021_, _12738_, _09454_);
  or (_22022_, _22021_, _21929_);
  and (_22023_, _22022_, _03785_);
  or (_22024_, _22023_, _03815_);
  or (_22025_, _22024_, _22020_);
  or (_22026_, _21935_, _04246_);
  and (_22027_, _22026_, _03823_);
  and (_22028_, _22027_, _22025_);
  and (_22029_, _21961_, _03453_);
  or (_22031_, _22029_, _03447_);
  or (_22032_, _22031_, _22028_);
  and (_22033_, _12794_, _05235_);
  or (_22034_, _21929_, _03514_);
  or (_22035_, _22034_, _22033_);
  and (_22036_, _22035_, _43000_);
  and (_22037_, _22036_, _22032_);
  nor (_22038_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_22039_, _22038_, _04794_);
  or (_43555_, _22039_, _22037_);
  nor (_22041_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_22042_, _22041_, _04794_);
  and (_22043_, _09454_, \oc8051_golden_model_1.P2 [4]);
  nor (_22044_, _05777_, _09454_);
  or (_22045_, _22044_, _22043_);
  or (_22046_, _22045_, _06838_);
  and (_22047_, _21946_, \oc8051_golden_model_1.P2 [4]);
  and (_22048_, _12827_, _05918_);
  or (_22049_, _22048_, _22047_);
  and (_22050_, _22049_, _03714_);
  nor (_22051_, _12841_, _09454_);
  or (_22052_, _22051_, _22043_);
  or (_22053_, _22052_, _04081_);
  and (_22054_, _05235_, \oc8051_golden_model_1.ACC [4]);
  or (_22055_, _22054_, _22043_);
  and (_22056_, _22055_, _04409_);
  and (_22057_, _09029_, \oc8051_golden_model_1.P2 [4]);
  or (_22058_, _22057_, _03610_);
  or (_22059_, _22058_, _22056_);
  and (_22060_, _22059_, _04055_);
  and (_22063_, _22060_, _22053_);
  and (_22064_, _12845_, _05918_);
  or (_22065_, _22064_, _22047_);
  and (_22066_, _22065_, _03715_);
  or (_22067_, _22066_, _03723_);
  or (_22068_, _22067_, _22063_);
  or (_22069_, _22045_, _03996_);
  and (_22070_, _22069_, _22068_);
  or (_22071_, _22070_, _03729_);
  or (_22072_, _22055_, _03737_);
  and (_22074_, _22072_, _03736_);
  and (_22075_, _22074_, _22071_);
  or (_22076_, _22075_, _22050_);
  and (_22077_, _22076_, _06840_);
  and (_22078_, _12861_, _05918_);
  or (_22079_, _22078_, _22047_);
  and (_22080_, _22079_, _03719_);
  or (_22081_, _22080_, _22077_);
  and (_22082_, _22081_, _03710_);
  and (_22083_, _20511_, _05918_);
  or (_22085_, _22083_, _22047_);
  and (_22086_, _22085_, _03505_);
  or (_22087_, _22086_, _07390_);
  or (_22088_, _22087_, _22082_);
  and (_22089_, _22088_, _22046_);
  or (_22090_, _22089_, _04481_);
  and (_22091_, _06730_, _05235_);
  or (_22092_, _22043_, _07400_);
  or (_22093_, _22092_, _22091_);
  and (_22094_, _22093_, _03589_);
  and (_22096_, _22094_, _22090_);
  and (_22097_, _20536_, _05235_);
  or (_22098_, _22097_, _22043_);
  and (_22099_, _22098_, _03222_);
  or (_22100_, _22099_, _08828_);
  or (_22101_, _22100_, _22096_);
  and (_22102_, _12821_, _05235_);
  or (_22103_, _22043_, _07766_);
  or (_22104_, _22103_, _22102_);
  and (_22105_, _06298_, _05235_);
  or (_22107_, _22105_, _22043_);
  or (_22108_, _22107_, _05886_);
  and (_22109_, _22108_, _07778_);
  and (_22110_, _22109_, _22104_);
  and (_22111_, _22110_, _22101_);
  and (_22112_, _12817_, _05235_);
  or (_22113_, _22112_, _22043_);
  and (_22114_, _22113_, _03780_);
  or (_22115_, _22114_, _22111_);
  and (_22116_, _22115_, _07777_);
  or (_22118_, _22043_, _05825_);
  and (_22119_, _22107_, _03622_);
  and (_22120_, _22119_, _22118_);
  or (_22121_, _22120_, _22116_);
  and (_22122_, _22121_, _06828_);
  and (_22123_, _22055_, _03790_);
  and (_22124_, _22123_, _22118_);
  or (_22125_, _22124_, _03624_);
  or (_22126_, _22125_, _22122_);
  nor (_22127_, _12819_, _09454_);
  or (_22129_, _22043_, _07795_);
  or (_22130_, _22129_, _22127_);
  and (_22131_, _22130_, _07793_);
  and (_22132_, _22131_, _22126_);
  nor (_22133_, _12816_, _09454_);
  or (_22134_, _22133_, _22043_);
  and (_22135_, _22134_, _03785_);
  or (_22136_, _22135_, _03815_);
  or (_22137_, _22136_, _22132_);
  or (_22138_, _22052_, _04246_);
  and (_22140_, _22138_, _03823_);
  and (_22141_, _22140_, _22137_);
  and (_22142_, _22049_, _03453_);
  or (_22143_, _22142_, _03447_);
  or (_22144_, _22143_, _22141_);
  and (_22145_, _13003_, _05235_);
  or (_22146_, _22043_, _03514_);
  or (_22147_, _22146_, _22145_);
  and (_22148_, _22147_, _43000_);
  and (_22149_, _22148_, _22144_);
  or (_43556_, _22149_, _22042_);
  and (_22151_, _09454_, \oc8051_golden_model_1.P2 [5]);
  nor (_22152_, _13014_, _09454_);
  or (_22153_, _22152_, _22151_);
  or (_22154_, _22153_, _04081_);
  and (_22155_, _05235_, \oc8051_golden_model_1.ACC [5]);
  or (_22156_, _22155_, _22151_);
  and (_22157_, _22156_, _04409_);
  and (_22158_, _09029_, \oc8051_golden_model_1.P2 [5]);
  or (_22159_, _22158_, _03610_);
  or (_22161_, _22159_, _22157_);
  and (_22162_, _22161_, _04055_);
  and (_22163_, _22162_, _22154_);
  and (_22164_, _21946_, \oc8051_golden_model_1.P2 [5]);
  and (_22165_, _13037_, _05918_);
  or (_22166_, _22165_, _22164_);
  and (_22167_, _22166_, _03715_);
  or (_22168_, _22167_, _03723_);
  or (_22169_, _22168_, _22163_);
  nor (_22170_, _05469_, _09454_);
  or (_22172_, _22170_, _22151_);
  or (_22173_, _22172_, _03996_);
  and (_22174_, _22173_, _22169_);
  or (_22175_, _22174_, _03729_);
  or (_22176_, _22156_, _03737_);
  and (_22177_, _22176_, _03736_);
  and (_22178_, _22177_, _22175_);
  and (_22179_, _13047_, _05918_);
  or (_22180_, _22179_, _22164_);
  and (_22181_, _22180_, _03714_);
  or (_22183_, _22181_, _03719_);
  or (_22184_, _22183_, _22178_);
  or (_22185_, _22164_, _13054_);
  and (_22186_, _22185_, _22166_);
  or (_22187_, _22186_, _06840_);
  and (_22188_, _22187_, _03710_);
  and (_22189_, _22188_, _22184_);
  and (_22190_, _20633_, _05918_);
  or (_22191_, _22190_, _22164_);
  and (_22192_, _22191_, _03505_);
  or (_22194_, _22192_, _07390_);
  or (_22195_, _22194_, _22189_);
  or (_22196_, _22172_, _06838_);
  and (_22197_, _22196_, _22195_);
  or (_22198_, _22197_, _04481_);
  and (_22199_, _06684_, _05235_);
  or (_22200_, _22151_, _07400_);
  or (_22201_, _22200_, _22199_);
  and (_22202_, _22201_, _03589_);
  and (_22203_, _22202_, _22198_);
  and (_22205_, _20660_, _05235_);
  or (_22206_, _22205_, _22151_);
  and (_22207_, _22206_, _03222_);
  or (_22208_, _22207_, _08828_);
  or (_22209_, _22208_, _22203_);
  and (_22210_, _13141_, _05235_);
  or (_22211_, _22151_, _07766_);
  or (_22212_, _22211_, _22210_);
  and (_22213_, _06306_, _05235_);
  or (_22214_, _22213_, _22151_);
  or (_22216_, _22214_, _05886_);
  and (_22217_, _22216_, _07778_);
  and (_22218_, _22217_, _22212_);
  and (_22219_, _22218_, _22209_);
  and (_22220_, _13147_, _05235_);
  or (_22221_, _22220_, _22151_);
  and (_22222_, _22221_, _03780_);
  or (_22223_, _22222_, _22219_);
  and (_22224_, _22223_, _07777_);
  or (_22225_, _22151_, _05518_);
  and (_22227_, _22214_, _03622_);
  and (_22228_, _22227_, _22225_);
  or (_22229_, _22228_, _22224_);
  and (_22230_, _22229_, _06828_);
  and (_22231_, _22156_, _03790_);
  and (_22232_, _22231_, _22225_);
  or (_22233_, _22232_, _03624_);
  or (_22234_, _22233_, _22230_);
  nor (_22235_, _13140_, _09454_);
  or (_22236_, _22151_, _07795_);
  or (_22238_, _22236_, _22235_);
  and (_22239_, _22238_, _07793_);
  and (_22240_, _22239_, _22234_);
  nor (_22241_, _13146_, _09454_);
  or (_22242_, _22241_, _22151_);
  and (_22243_, _22242_, _03785_);
  or (_22244_, _22243_, _03815_);
  or (_22245_, _22244_, _22240_);
  or (_22246_, _22153_, _04246_);
  and (_22247_, _22246_, _03823_);
  and (_22249_, _22247_, _22245_);
  and (_22250_, _22180_, _03453_);
  or (_22251_, _22250_, _03447_);
  or (_22252_, _22251_, _22249_);
  and (_22253_, _13199_, _05235_);
  or (_22254_, _22151_, _03514_);
  or (_22255_, _22254_, _22253_);
  and (_22256_, _22255_, _43000_);
  and (_22257_, _22256_, _22252_);
  nor (_22258_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_22260_, _22258_, _04794_);
  or (_43557_, _22260_, _22257_);
  not (_22261_, \oc8051_golden_model_1.P2 [6]);
  nor (_22262_, _43000_, _22261_);
  or (_22263_, _22262_, rst);
  nor (_22264_, _05235_, _22261_);
  nor (_22265_, _13242_, _09454_);
  or (_22266_, _22265_, _22264_);
  or (_22267_, _22266_, _04081_);
  and (_22268_, _05235_, \oc8051_golden_model_1.ACC [6]);
  or (_22270_, _22268_, _22264_);
  and (_22271_, _22270_, _04409_);
  nor (_22272_, _04409_, _22261_);
  or (_22273_, _22272_, _03610_);
  or (_22274_, _22273_, _22271_);
  and (_22275_, _22274_, _04055_);
  and (_22276_, _22275_, _22267_);
  nor (_22277_, _05918_, _22261_);
  and (_22278_, _13229_, _05918_);
  or (_22279_, _22278_, _22277_);
  and (_22281_, _22279_, _03715_);
  or (_22282_, _22281_, _03723_);
  or (_22283_, _22282_, _22276_);
  nor (_22284_, _05363_, _09454_);
  or (_22285_, _22284_, _22264_);
  or (_22286_, _22285_, _03996_);
  and (_22287_, _22286_, _22283_);
  or (_22288_, _22287_, _03729_);
  or (_22289_, _22270_, _03737_);
  and (_22290_, _22289_, _03736_);
  and (_22292_, _22290_, _22288_);
  and (_22293_, _13253_, _05918_);
  or (_22294_, _22293_, _22277_);
  and (_22295_, _22294_, _03714_);
  or (_22296_, _22295_, _03719_);
  or (_22297_, _22296_, _22292_);
  or (_22298_, _22277_, _13260_);
  and (_22299_, _22298_, _22279_);
  or (_22300_, _22299_, _06840_);
  and (_22301_, _22300_, _03710_);
  and (_22303_, _22301_, _22297_);
  and (_22304_, _20753_, _05918_);
  or (_22305_, _22304_, _22277_);
  and (_22306_, _22305_, _03505_);
  or (_22307_, _22306_, _07390_);
  or (_22308_, _22307_, _22303_);
  or (_22309_, _22285_, _06838_);
  and (_22310_, _22309_, _22308_);
  or (_22311_, _22310_, _04481_);
  and (_22312_, _06455_, _05235_);
  or (_22314_, _22264_, _07400_);
  or (_22315_, _22314_, _22312_);
  and (_22316_, _22315_, _03589_);
  and (_22317_, _22316_, _22311_);
  and (_22318_, _20778_, _05235_);
  or (_22319_, _22318_, _22264_);
  and (_22320_, _22319_, _03222_);
  or (_22321_, _22320_, _08828_);
  or (_22322_, _22321_, _22317_);
  and (_22323_, _13347_, _05235_);
  or (_22326_, _22264_, _07766_);
  or (_22327_, _22326_, _22323_);
  and (_22328_, _13339_, _05235_);
  or (_22329_, _22328_, _22264_);
  or (_22330_, _22329_, _05886_);
  and (_22331_, _22330_, _07778_);
  and (_22332_, _22331_, _22327_);
  and (_22333_, _22332_, _22322_);
  and (_22334_, _13353_, _05235_);
  or (_22335_, _22334_, _22264_);
  and (_22337_, _22335_, _03780_);
  or (_22338_, _22337_, _22333_);
  and (_22339_, _22338_, _07777_);
  or (_22340_, _22264_, _05412_);
  and (_22341_, _22329_, _03622_);
  and (_22342_, _22341_, _22340_);
  or (_22343_, _22342_, _22339_);
  and (_22344_, _22343_, _06828_);
  and (_22345_, _22270_, _03790_);
  and (_22346_, _22345_, _22340_);
  or (_22348_, _22346_, _03624_);
  or (_22349_, _22348_, _22344_);
  nor (_22350_, _13346_, _09454_);
  or (_22351_, _22264_, _07795_);
  or (_22352_, _22351_, _22350_);
  and (_22353_, _22352_, _07793_);
  and (_22354_, _22353_, _22349_);
  nor (_22355_, _13352_, _09454_);
  or (_22356_, _22355_, _22264_);
  and (_22357_, _22356_, _03785_);
  or (_22359_, _22357_, _03815_);
  or (_22360_, _22359_, _22354_);
  or (_22361_, _22266_, _04246_);
  and (_22362_, _22361_, _03823_);
  and (_22363_, _22362_, _22360_);
  and (_22364_, _22294_, _03453_);
  or (_22365_, _22364_, _03447_);
  or (_22366_, _22365_, _22363_);
  and (_22367_, _13402_, _05235_);
  or (_22368_, _22264_, _03514_);
  or (_22370_, _22368_, _22367_);
  and (_22371_, _22370_, _43000_);
  and (_22372_, _22371_, _22366_);
  or (_43558_, _22372_, _22263_);
  not (_22373_, \oc8051_golden_model_1.P3 [0]);
  nor (_22374_, _05239_, _22373_);
  and (_22375_, _12128_, _05239_);
  or (_22376_, _22375_, _22374_);
  and (_22377_, _22376_, _03780_);
  and (_22378_, _05239_, _04620_);
  or (_22380_, _22378_, _22374_);
  or (_22381_, _22380_, _06838_);
  nor (_22382_, _05666_, _09557_);
  or (_22383_, _22382_, _22374_);
  or (_22384_, _22383_, _04081_);
  and (_22385_, _05239_, \oc8051_golden_model_1.ACC [0]);
  or (_22386_, _22385_, _22374_);
  and (_22387_, _22386_, _04409_);
  nor (_22388_, _04409_, _22373_);
  or (_22389_, _22388_, _03610_);
  or (_22391_, _22389_, _22387_);
  and (_22392_, _22391_, _04055_);
  and (_22393_, _22392_, _22384_);
  nor (_22394_, _05929_, _22373_);
  and (_22395_, _12021_, _05929_);
  or (_22396_, _22395_, _22394_);
  and (_22397_, _22396_, _03715_);
  or (_22398_, _22397_, _22393_);
  and (_22399_, _22398_, _03996_);
  and (_22400_, _22380_, _03723_);
  or (_22402_, _22400_, _03729_);
  or (_22403_, _22402_, _22399_);
  or (_22404_, _22386_, _03737_);
  and (_22405_, _22404_, _03736_);
  and (_22406_, _22405_, _22403_);
  and (_22407_, _22374_, _03714_);
  or (_22408_, _22407_, _03719_);
  or (_22409_, _22408_, _22406_);
  or (_22410_, _22383_, _06840_);
  and (_22411_, _22410_, _03710_);
  and (_22413_, _22411_, _22409_);
  and (_22414_, _20023_, _05929_);
  or (_22415_, _22414_, _22394_);
  and (_22416_, _22415_, _03505_);
  or (_22417_, _22416_, _07390_);
  or (_22418_, _22417_, _22413_);
  and (_22419_, _22418_, _22381_);
  or (_22420_, _22419_, _04481_);
  and (_22421_, _06546_, _05239_);
  or (_22422_, _22374_, _07400_);
  or (_22424_, _22422_, _22421_);
  and (_22425_, _22424_, _03589_);
  and (_22426_, _22425_, _22420_);
  and (_22427_, _20049_, _05239_);
  or (_22428_, _22427_, _22374_);
  and (_22429_, _22428_, _03222_);
  or (_22430_, _22429_, _22426_);
  or (_22431_, _22430_, _08828_);
  and (_22432_, _12124_, _05239_);
  or (_22433_, _22374_, _07766_);
  or (_22436_, _22433_, _22432_);
  and (_22437_, _05239_, _06274_);
  or (_22438_, _22437_, _22374_);
  or (_22439_, _22438_, _05886_);
  and (_22440_, _22439_, _07778_);
  and (_22441_, _22440_, _22436_);
  and (_22442_, _22441_, _22431_);
  or (_22443_, _22442_, _22377_);
  and (_22444_, _22443_, _07777_);
  nand (_22445_, _22438_, _03622_);
  nor (_22447_, _22445_, _22382_);
  or (_22448_, _22447_, _22444_);
  and (_22449_, _22448_, _06828_);
  or (_22450_, _22374_, _05666_);
  and (_22451_, _22386_, _03790_);
  and (_22452_, _22451_, _22450_);
  or (_22453_, _22452_, _03624_);
  or (_22454_, _22453_, _22449_);
  nor (_22455_, _12122_, _09557_);
  or (_22456_, _22374_, _07795_);
  or (_22458_, _22456_, _22455_);
  and (_22459_, _22458_, _07793_);
  and (_22460_, _22459_, _22454_);
  nor (_22461_, _12003_, _09557_);
  or (_22462_, _22461_, _22374_);
  and (_22463_, _22462_, _03785_);
  or (_22464_, _22463_, _03815_);
  or (_22465_, _22464_, _22460_);
  or (_22466_, _22383_, _04246_);
  and (_22467_, _22466_, _03823_);
  and (_22469_, _22467_, _22465_);
  and (_22470_, _22374_, _03453_);
  or (_22471_, _22470_, _03447_);
  or (_22472_, _22471_, _22469_);
  or (_22473_, _22383_, _03514_);
  and (_22474_, _22473_, _43000_);
  and (_22475_, _22474_, _22472_);
  nor (_22476_, _43000_, _22373_);
  or (_22477_, _22476_, rst);
  or (_43561_, _22477_, _22475_);
  or (_22479_, _05239_, \oc8051_golden_model_1.P3 [1]);
  and (_22480_, _12213_, _05239_);
  not (_22481_, _22480_);
  and (_22482_, _22481_, _22479_);
  or (_22483_, _22482_, _04081_);
  nand (_22484_, _05239_, _03274_);
  and (_22485_, _22484_, _22479_);
  and (_22486_, _22485_, _04409_);
  not (_22487_, \oc8051_golden_model_1.P3 [1]);
  nor (_22488_, _04409_, _22487_);
  or (_22490_, _22488_, _03610_);
  or (_22491_, _22490_, _22486_);
  and (_22492_, _22491_, _04055_);
  and (_22493_, _22492_, _22483_);
  and (_22494_, _12224_, _05929_);
  nor (_22495_, _05929_, _22487_);
  or (_22496_, _22495_, _03723_);
  or (_22497_, _22496_, _22494_);
  and (_22498_, _22497_, _14265_);
  or (_22499_, _22498_, _22493_);
  nor (_22501_, _05239_, _22487_);
  and (_22502_, _05239_, _06764_);
  or (_22503_, _22502_, _22501_);
  or (_22504_, _22503_, _03996_);
  and (_22505_, _22504_, _22499_);
  or (_22506_, _22505_, _03729_);
  or (_22507_, _22485_, _03737_);
  and (_22508_, _22507_, _03736_);
  and (_22509_, _22508_, _22506_);
  and (_22510_, _12211_, _05929_);
  or (_22512_, _22510_, _22495_);
  and (_22513_, _22512_, _03714_);
  or (_22514_, _22513_, _03719_);
  or (_22515_, _22514_, _22509_);
  and (_22516_, _22494_, _12239_);
  or (_22517_, _22495_, _06840_);
  or (_22518_, _22517_, _22516_);
  and (_22519_, _22518_, _22515_);
  and (_22520_, _22519_, _03710_);
  and (_22521_, _20141_, _05929_);
  or (_22523_, _22495_, _22521_);
  and (_22524_, _22523_, _03505_);
  or (_22525_, _22524_, _07390_);
  or (_22526_, _22525_, _22520_);
  or (_22527_, _22503_, _06838_);
  and (_22528_, _22527_, _22526_);
  or (_22529_, _22528_, _04481_);
  and (_22530_, _06501_, _05239_);
  or (_22531_, _22501_, _07400_);
  or (_22532_, _22531_, _22530_);
  and (_22534_, _22532_, _03589_);
  and (_22535_, _22534_, _22529_);
  and (_22536_, _20168_, _05239_);
  or (_22537_, _22536_, _22501_);
  and (_22538_, _22537_, _03222_);
  or (_22539_, _22538_, _22535_);
  and (_22540_, _22539_, _03602_);
  or (_22541_, _12327_, _09557_);
  and (_22542_, _22541_, _03600_);
  nand (_22543_, _05239_, _04303_);
  and (_22545_, _22543_, _03601_);
  or (_22546_, _22545_, _22542_);
  and (_22547_, _22546_, _22479_);
  or (_22548_, _22547_, _22540_);
  and (_22549_, _22548_, _07778_);
  or (_22550_, _12333_, _09557_);
  and (_22551_, _22479_, _03780_);
  and (_22552_, _22551_, _22550_);
  or (_22553_, _22552_, _22549_);
  and (_22554_, _22553_, _07777_);
  or (_22556_, _12207_, _09557_);
  and (_22557_, _22479_, _03622_);
  and (_22558_, _22557_, _22556_);
  or (_22559_, _22558_, _22554_);
  and (_22560_, _22559_, _06828_);
  or (_22561_, _22501_, _05618_);
  and (_22562_, _22485_, _03790_);
  and (_22563_, _22562_, _22561_);
  or (_22564_, _22563_, _22560_);
  and (_22565_, _22564_, _03786_);
  or (_22567_, _22543_, _05618_);
  and (_22568_, _22479_, _03624_);
  and (_22569_, _22568_, _22567_);
  or (_22570_, _22484_, _05618_);
  and (_22571_, _22479_, _03785_);
  and (_22572_, _22571_, _22570_);
  or (_22573_, _22572_, _03815_);
  or (_22574_, _22573_, _22569_);
  or (_22575_, _22574_, _22565_);
  or (_22576_, _22482_, _04246_);
  and (_22578_, _22576_, _03823_);
  and (_22579_, _22578_, _22575_);
  and (_22580_, _22512_, _03453_);
  or (_22581_, _22580_, _03447_);
  or (_22582_, _22581_, _22579_);
  or (_22583_, _22501_, _03514_);
  or (_22584_, _22583_, _22480_);
  and (_22585_, _22584_, _43000_);
  and (_22586_, _22585_, _22582_);
  nor (_22587_, _43000_, _22487_);
  or (_22589_, _22587_, rst);
  or (_43562_, _22589_, _22586_);
  not (_22590_, \oc8051_golden_model_1.P3 [2]);
  nor (_22591_, _05239_, _22590_);
  nor (_22592_, _09557_, _04875_);
  or (_22593_, _22592_, _22591_);
  or (_22594_, _22593_, _06838_);
  and (_22595_, _22593_, _03723_);
  nor (_22596_, _05929_, _22590_);
  and (_22597_, _12411_, _05929_);
  or (_22599_, _22597_, _22596_);
  or (_22600_, _22599_, _04055_);
  nor (_22601_, _12416_, _09557_);
  or (_22602_, _22601_, _22591_);
  and (_22603_, _22602_, _03610_);
  nor (_22604_, _04409_, _22590_);
  and (_22605_, _05239_, \oc8051_golden_model_1.ACC [2]);
  or (_22606_, _22605_, _22591_);
  and (_22607_, _22606_, _04409_);
  or (_22608_, _22607_, _22604_);
  and (_22610_, _22608_, _04081_);
  or (_22611_, _22610_, _03715_);
  or (_22612_, _22611_, _22603_);
  and (_22613_, _22612_, _22600_);
  and (_22614_, _22613_, _03996_);
  or (_22615_, _22614_, _22595_);
  or (_22616_, _22615_, _03729_);
  or (_22617_, _22606_, _03737_);
  and (_22618_, _22617_, _03736_);
  and (_22619_, _22618_, _22616_);
  and (_22621_, _12409_, _05929_);
  or (_22622_, _22621_, _22596_);
  and (_22623_, _22622_, _03714_);
  or (_22624_, _22623_, _03719_);
  or (_22625_, _22624_, _22619_);
  or (_22626_, _22596_, _12443_);
  and (_22627_, _22626_, _22599_);
  or (_22628_, _22627_, _06840_);
  and (_22629_, _22628_, _03710_);
  and (_22630_, _22629_, _22625_);
  and (_22632_, _20264_, _05929_);
  or (_22633_, _22632_, _22596_);
  and (_22634_, _22633_, _03505_);
  or (_22635_, _22634_, _07390_);
  or (_22636_, _22635_, _22630_);
  and (_22637_, _22636_, _22594_);
  or (_22638_, _22637_, _04481_);
  and (_22639_, _06637_, _05239_);
  or (_22640_, _22591_, _07400_);
  or (_22641_, _22640_, _22639_);
  and (_22643_, _22641_, _03589_);
  and (_22644_, _22643_, _22638_);
  and (_22645_, _20290_, _05239_);
  or (_22646_, _22591_, _22645_);
  and (_22647_, _22646_, _03222_);
  or (_22648_, _22647_, _22644_);
  or (_22649_, _22648_, _08828_);
  and (_22650_, _12533_, _05239_);
  or (_22651_, _22591_, _07766_);
  or (_22652_, _22651_, _22650_);
  and (_22654_, _05239_, _06332_);
  or (_22655_, _22654_, _22591_);
  or (_22656_, _22655_, _05886_);
  and (_22657_, _22656_, _07778_);
  and (_22658_, _22657_, _22652_);
  and (_22659_, _22658_, _22649_);
  and (_22660_, _12539_, _05239_);
  or (_22661_, _22660_, _22591_);
  and (_22662_, _22661_, _03780_);
  or (_22663_, _22662_, _22659_);
  and (_22665_, _22663_, _07777_);
  or (_22666_, _22591_, _05718_);
  and (_22667_, _22655_, _03622_);
  and (_22668_, _22667_, _22666_);
  or (_22669_, _22668_, _22665_);
  and (_22670_, _22669_, _06828_);
  and (_22671_, _22606_, _03790_);
  and (_22672_, _22671_, _22666_);
  or (_22673_, _22672_, _03624_);
  or (_22674_, _22673_, _22670_);
  nor (_22676_, _12532_, _09557_);
  or (_22677_, _22591_, _07795_);
  or (_22678_, _22677_, _22676_);
  and (_22679_, _22678_, _07793_);
  and (_22680_, _22679_, _22674_);
  nor (_22681_, _12538_, _09557_);
  or (_22682_, _22681_, _22591_);
  and (_22683_, _22682_, _03785_);
  or (_22684_, _22683_, _03815_);
  or (_22685_, _22684_, _22680_);
  or (_22687_, _22602_, _04246_);
  and (_22688_, _22687_, _03823_);
  and (_22689_, _22688_, _22685_);
  and (_22690_, _22622_, _03453_);
  or (_22691_, _22690_, _03447_);
  or (_22692_, _22691_, _22689_);
  and (_22693_, _12592_, _05239_);
  or (_22694_, _22591_, _03514_);
  or (_22695_, _22694_, _22693_);
  and (_22696_, _22695_, _43000_);
  and (_22698_, _22696_, _22692_);
  nor (_22699_, _43000_, _22590_);
  or (_22700_, _22699_, rst);
  or (_43563_, _22700_, _22698_);
  and (_22701_, _09557_, \oc8051_golden_model_1.P3 [3]);
  nor (_22702_, _09557_, _05005_);
  or (_22703_, _22702_, _22701_);
  or (_22704_, _22703_, _06838_);
  nor (_22705_, _12627_, _09557_);
  or (_22706_, _22705_, _22701_);
  or (_22708_, _22706_, _04081_);
  and (_22709_, _05239_, \oc8051_golden_model_1.ACC [3]);
  or (_22710_, _22709_, _22701_);
  and (_22711_, _22710_, _04409_);
  and (_22712_, _09029_, \oc8051_golden_model_1.P3 [3]);
  or (_22713_, _22712_, _03610_);
  or (_22714_, _22713_, _22711_);
  and (_22715_, _22714_, _04055_);
  and (_22716_, _22715_, _22708_);
  not (_22717_, _05929_);
  and (_22719_, _22717_, \oc8051_golden_model_1.P3 [3]);
  and (_22720_, _12631_, _05929_);
  or (_22721_, _22720_, _22719_);
  and (_22722_, _22721_, _03715_);
  or (_22723_, _22722_, _03723_);
  or (_22724_, _22723_, _22716_);
  or (_22725_, _22703_, _03996_);
  and (_22726_, _22725_, _22724_);
  or (_22727_, _22726_, _03729_);
  or (_22728_, _22710_, _03737_);
  and (_22730_, _22728_, _03736_);
  and (_22731_, _22730_, _22727_);
  and (_22732_, _12641_, _05929_);
  or (_22733_, _22732_, _22719_);
  and (_22734_, _22733_, _03714_);
  or (_22735_, _22734_, _03719_);
  or (_22736_, _22735_, _22731_);
  or (_22737_, _22719_, _12648_);
  and (_22738_, _22737_, _22721_);
  or (_22739_, _22738_, _06840_);
  and (_22741_, _22739_, _03710_);
  and (_22742_, _22741_, _22736_);
  and (_22743_, _20391_, _05929_);
  or (_22744_, _22743_, _22719_);
  and (_22745_, _22744_, _03505_);
  or (_22746_, _22745_, _07390_);
  or (_22747_, _22746_, _22742_);
  and (_22748_, _22747_, _22704_);
  or (_22749_, _22748_, _04481_);
  and (_22750_, _06592_, _05239_);
  or (_22752_, _22701_, _07400_);
  or (_22753_, _22752_, _22750_);
  and (_22754_, _22753_, _03589_);
  and (_22755_, _22754_, _22749_);
  and (_22756_, _20416_, _05239_);
  or (_22757_, _22701_, _22756_);
  and (_22758_, _22757_, _03222_);
  or (_22759_, _22758_, _22755_);
  or (_22760_, _22759_, _08828_);
  and (_22761_, _12733_, _05239_);
  or (_22763_, _22701_, _07766_);
  or (_22764_, _22763_, _22761_);
  and (_22765_, _05239_, _06276_);
  or (_22766_, _22765_, _22701_);
  or (_22767_, _22766_, _05886_);
  and (_22768_, _22767_, _07778_);
  and (_22769_, _22768_, _22764_);
  and (_22770_, _22769_, _22760_);
  and (_22771_, _12739_, _05239_);
  or (_22772_, _22771_, _22701_);
  and (_22774_, _22772_, _03780_);
  or (_22775_, _22774_, _22770_);
  and (_22776_, _22775_, _07777_);
  or (_22777_, _22701_, _05567_);
  and (_22778_, _22766_, _03622_);
  and (_22779_, _22778_, _22777_);
  or (_22780_, _22779_, _22776_);
  and (_22781_, _22780_, _06828_);
  and (_22782_, _22710_, _03790_);
  and (_22783_, _22782_, _22777_);
  or (_22785_, _22783_, _03624_);
  or (_22786_, _22785_, _22781_);
  nor (_22787_, _12732_, _09557_);
  or (_22788_, _22701_, _07795_);
  or (_22789_, _22788_, _22787_);
  and (_22790_, _22789_, _07793_);
  and (_22791_, _22790_, _22786_);
  nor (_22792_, _12738_, _09557_);
  or (_22793_, _22792_, _22701_);
  and (_22794_, _22793_, _03785_);
  or (_22796_, _22794_, _03815_);
  or (_22797_, _22796_, _22791_);
  or (_22798_, _22706_, _04246_);
  and (_22799_, _22798_, _03823_);
  and (_22800_, _22799_, _22797_);
  and (_22801_, _22733_, _03453_);
  or (_22802_, _22801_, _03447_);
  or (_22803_, _22802_, _22800_);
  and (_22804_, _12794_, _05239_);
  or (_22805_, _22701_, _03514_);
  or (_22807_, _22805_, _22804_);
  and (_22808_, _22807_, _43000_);
  and (_22809_, _22808_, _22803_);
  nor (_22810_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_22811_, _22810_, _04794_);
  or (_43564_, _22811_, _22809_);
  and (_22812_, _09557_, \oc8051_golden_model_1.P3 [4]);
  nor (_22813_, _05777_, _09557_);
  or (_22814_, _22813_, _22812_);
  or (_22815_, _22814_, _06838_);
  and (_22817_, _22717_, \oc8051_golden_model_1.P3 [4]);
  and (_22818_, _12827_, _05929_);
  or (_22819_, _22818_, _22817_);
  and (_22820_, _22819_, _03714_);
  nor (_22821_, _12841_, _09557_);
  or (_22822_, _22821_, _22812_);
  or (_22823_, _22822_, _04081_);
  and (_22824_, _05239_, \oc8051_golden_model_1.ACC [4]);
  or (_22825_, _22824_, _22812_);
  and (_22826_, _22825_, _04409_);
  and (_22828_, _09029_, \oc8051_golden_model_1.P3 [4]);
  or (_22829_, _22828_, _03610_);
  or (_22830_, _22829_, _22826_);
  and (_22831_, _22830_, _04055_);
  and (_22832_, _22831_, _22823_);
  and (_22833_, _12845_, _05929_);
  or (_22834_, _22833_, _22817_);
  and (_22835_, _22834_, _03715_);
  or (_22836_, _22835_, _03723_);
  or (_22837_, _22836_, _22832_);
  or (_22839_, _22814_, _03996_);
  and (_22840_, _22839_, _22837_);
  or (_22841_, _22840_, _03729_);
  or (_22842_, _22825_, _03737_);
  and (_22843_, _22842_, _03736_);
  and (_22844_, _22843_, _22841_);
  or (_22845_, _22844_, _22820_);
  and (_22846_, _22845_, _06840_);
  or (_22847_, _22817_, _12860_);
  and (_22848_, _22847_, _03719_);
  and (_22850_, _22848_, _22834_);
  or (_22851_, _22850_, _22846_);
  and (_22852_, _22851_, _03710_);
  and (_22853_, _20511_, _05929_);
  or (_22854_, _22853_, _22817_);
  and (_22855_, _22854_, _03505_);
  or (_22856_, _22855_, _07390_);
  or (_22857_, _22856_, _22852_);
  and (_22858_, _22857_, _22815_);
  or (_22859_, _22858_, _04481_);
  and (_22861_, _06730_, _05239_);
  or (_22862_, _22812_, _07400_);
  or (_22863_, _22862_, _22861_);
  and (_22864_, _22863_, _03589_);
  and (_22865_, _22864_, _22859_);
  and (_22866_, _20536_, _05239_);
  or (_22867_, _22866_, _22812_);
  and (_22868_, _22867_, _03222_);
  or (_22869_, _22868_, _08828_);
  or (_22870_, _22869_, _22865_);
  and (_22872_, _12821_, _05239_);
  or (_22873_, _22812_, _07766_);
  or (_22874_, _22873_, _22872_);
  and (_22875_, _06298_, _05239_);
  or (_22876_, _22875_, _22812_);
  or (_22877_, _22876_, _05886_);
  and (_22878_, _22877_, _07778_);
  and (_22879_, _22878_, _22874_);
  and (_22880_, _22879_, _22870_);
  and (_22881_, _12817_, _05239_);
  or (_22883_, _22881_, _22812_);
  and (_22884_, _22883_, _03780_);
  or (_22885_, _22884_, _22880_);
  and (_22886_, _22885_, _07777_);
  or (_22887_, _22812_, _05825_);
  and (_22888_, _22876_, _03622_);
  and (_22889_, _22888_, _22887_);
  or (_22890_, _22889_, _22886_);
  and (_22891_, _22890_, _06828_);
  and (_22892_, _22825_, _03790_);
  and (_22894_, _22892_, _22887_);
  or (_22895_, _22894_, _03624_);
  or (_22896_, _22895_, _22891_);
  nor (_22897_, _12819_, _09557_);
  or (_22898_, _22812_, _07795_);
  or (_22899_, _22898_, _22897_);
  and (_22900_, _22899_, _07793_);
  and (_22901_, _22900_, _22896_);
  nor (_22902_, _12816_, _09557_);
  or (_22903_, _22902_, _22812_);
  and (_22905_, _22903_, _03785_);
  or (_22906_, _22905_, _03815_);
  or (_22907_, _22906_, _22901_);
  or (_22908_, _22822_, _04246_);
  and (_22909_, _22908_, _03823_);
  and (_22910_, _22909_, _22907_);
  and (_22911_, _22819_, _03453_);
  or (_22912_, _22911_, _03447_);
  or (_22913_, _22912_, _22910_);
  and (_22914_, _13003_, _05239_);
  or (_22916_, _22812_, _03514_);
  or (_22917_, _22916_, _22914_);
  and (_22918_, _22917_, _43000_);
  and (_22919_, _22918_, _22913_);
  nor (_22920_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_22921_, _22920_, _04794_);
  or (_43565_, _22921_, _22919_);
  nor (_22922_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_22923_, _22922_, _04794_);
  and (_22924_, _09557_, \oc8051_golden_model_1.P3 [5]);
  nor (_22926_, _13014_, _09557_);
  or (_22927_, _22926_, _22924_);
  or (_22928_, _22927_, _04081_);
  and (_22929_, _05239_, \oc8051_golden_model_1.ACC [5]);
  or (_22930_, _22929_, _22924_);
  and (_22931_, _22930_, _04409_);
  and (_22932_, _09029_, \oc8051_golden_model_1.P3 [5]);
  or (_22933_, _22932_, _03610_);
  or (_22934_, _22933_, _22931_);
  and (_22935_, _22934_, _04055_);
  and (_22937_, _22935_, _22928_);
  and (_22938_, _22717_, \oc8051_golden_model_1.P3 [5]);
  and (_22939_, _13037_, _05929_);
  or (_22940_, _22939_, _22938_);
  and (_22941_, _22940_, _03715_);
  or (_22942_, _22941_, _03723_);
  or (_22943_, _22942_, _22937_);
  nor (_22944_, _05469_, _09557_);
  or (_22945_, _22944_, _22924_);
  or (_22946_, _22945_, _03996_);
  and (_22948_, _22946_, _22943_);
  or (_22949_, _22948_, _03729_);
  or (_22950_, _22930_, _03737_);
  and (_22951_, _22950_, _03736_);
  and (_22952_, _22951_, _22949_);
  and (_22953_, _13047_, _05929_);
  or (_22954_, _22953_, _22938_);
  and (_22955_, _22954_, _03714_);
  or (_22956_, _22955_, _03719_);
  or (_22957_, _22956_, _22952_);
  or (_22959_, _22938_, _13054_);
  and (_22960_, _22959_, _22940_);
  or (_22961_, _22960_, _06840_);
  and (_22962_, _22961_, _03710_);
  and (_22963_, _22962_, _22957_);
  and (_22964_, _20633_, _05929_);
  or (_22965_, _22964_, _22938_);
  and (_22966_, _22965_, _03505_);
  or (_22967_, _22966_, _07390_);
  or (_22968_, _22967_, _22963_);
  or (_22970_, _22945_, _06838_);
  and (_22971_, _22970_, _22968_);
  or (_22972_, _22971_, _04481_);
  and (_22973_, _06684_, _05239_);
  or (_22974_, _22924_, _07400_);
  or (_22975_, _22974_, _22973_);
  and (_22976_, _22975_, _03589_);
  and (_22977_, _22976_, _22972_);
  and (_22978_, _20660_, _05239_);
  or (_22979_, _22978_, _22924_);
  and (_22981_, _22979_, _03222_);
  or (_22982_, _22981_, _08828_);
  or (_22983_, _22982_, _22977_);
  and (_22984_, _13141_, _05239_);
  or (_22985_, _22924_, _07766_);
  or (_22986_, _22985_, _22984_);
  and (_22987_, _06306_, _05239_);
  or (_22988_, _22987_, _22924_);
  or (_22989_, _22988_, _05886_);
  and (_22990_, _22989_, _07778_);
  and (_22991_, _22990_, _22986_);
  and (_22992_, _22991_, _22983_);
  and (_22993_, _13147_, _05239_);
  or (_22994_, _22993_, _22924_);
  and (_22995_, _22994_, _03780_);
  or (_22996_, _22995_, _22992_);
  and (_22997_, _22996_, _07777_);
  or (_22998_, _22924_, _05518_);
  and (_22999_, _22988_, _03622_);
  and (_23000_, _22999_, _22998_);
  or (_23003_, _23000_, _22997_);
  and (_23004_, _23003_, _06828_);
  and (_23005_, _22930_, _03790_);
  and (_23006_, _23005_, _22998_);
  or (_23007_, _23006_, _03624_);
  or (_23008_, _23007_, _23004_);
  nor (_23009_, _13140_, _09557_);
  or (_23010_, _22924_, _07795_);
  or (_23011_, _23010_, _23009_);
  and (_23012_, _23011_, _07793_);
  and (_23014_, _23012_, _23008_);
  nor (_23015_, _13146_, _09557_);
  or (_23016_, _23015_, _22924_);
  and (_23017_, _23016_, _03785_);
  or (_23018_, _23017_, _03815_);
  or (_23019_, _23018_, _23014_);
  or (_23020_, _22927_, _04246_);
  and (_23021_, _23020_, _03823_);
  and (_23022_, _23021_, _23019_);
  and (_23023_, _22954_, _03453_);
  or (_23024_, _23023_, _03447_);
  or (_23025_, _23024_, _23022_);
  and (_23026_, _13199_, _05239_);
  or (_23027_, _22924_, _03514_);
  or (_23028_, _23027_, _23026_);
  and (_23029_, _23028_, _43000_);
  and (_23030_, _23029_, _23025_);
  or (_43566_, _23030_, _22923_);
  not (_23031_, \oc8051_golden_model_1.P3 [6]);
  nor (_23032_, _05239_, _23031_);
  nor (_23035_, _13242_, _09557_);
  or (_23036_, _23035_, _23032_);
  or (_23037_, _23036_, _04081_);
  and (_23038_, _05239_, \oc8051_golden_model_1.ACC [6]);
  or (_23039_, _23038_, _23032_);
  and (_23040_, _23039_, _04409_);
  nor (_23041_, _04409_, _23031_);
  or (_23042_, _23041_, _03610_);
  or (_23043_, _23042_, _23040_);
  and (_23044_, _23043_, _04055_);
  and (_23046_, _23044_, _23037_);
  nor (_23047_, _05929_, _23031_);
  and (_23048_, _13229_, _05929_);
  or (_23049_, _23048_, _23047_);
  and (_23050_, _23049_, _03715_);
  or (_23051_, _23050_, _03723_);
  or (_23052_, _23051_, _23046_);
  nor (_23053_, _05363_, _09557_);
  or (_23054_, _23053_, _23032_);
  or (_23055_, _23054_, _03996_);
  and (_23056_, _23055_, _23052_);
  or (_23057_, _23056_, _03729_);
  or (_23058_, _23039_, _03737_);
  and (_23059_, _23058_, _03736_);
  and (_23060_, _23059_, _23057_);
  and (_23061_, _13253_, _05929_);
  or (_23062_, _23061_, _23047_);
  and (_23063_, _23062_, _03714_);
  or (_23064_, _23063_, _03719_);
  or (_23065_, _23064_, _23060_);
  or (_23068_, _23047_, _13260_);
  and (_23069_, _23068_, _23049_);
  or (_23070_, _23069_, _06840_);
  and (_23071_, _23070_, _03710_);
  and (_23072_, _23071_, _23065_);
  and (_23073_, _20753_, _05929_);
  or (_23074_, _23073_, _23047_);
  and (_23075_, _23074_, _03505_);
  or (_23076_, _23075_, _07390_);
  or (_23077_, _23076_, _23072_);
  or (_23079_, _23054_, _06838_);
  and (_23080_, _23079_, _23077_);
  or (_23081_, _23080_, _04481_);
  and (_23082_, _06455_, _05239_);
  or (_23083_, _23032_, _07400_);
  or (_23084_, _23083_, _23082_);
  and (_23085_, _23084_, _03589_);
  and (_23086_, _23085_, _23081_);
  and (_23087_, _20778_, _05239_);
  or (_23088_, _23087_, _23032_);
  and (_23089_, _23088_, _03222_);
  or (_23090_, _23089_, _08828_);
  or (_23091_, _23090_, _23086_);
  and (_23092_, _13347_, _05239_);
  or (_23093_, _23032_, _07766_);
  or (_23094_, _23093_, _23092_);
  and (_23095_, _13339_, _05239_);
  or (_23096_, _23095_, _23032_);
  or (_23097_, _23096_, _05886_);
  and (_23098_, _23097_, _07778_);
  and (_23101_, _23098_, _23094_);
  and (_23102_, _23101_, _23091_);
  and (_23103_, _13353_, _05239_);
  or (_23104_, _23103_, _23032_);
  and (_23105_, _23104_, _03780_);
  or (_23106_, _23105_, _23102_);
  and (_23107_, _23106_, _07777_);
  or (_23108_, _23032_, _05412_);
  and (_23109_, _23096_, _03622_);
  and (_23110_, _23109_, _23108_);
  or (_23112_, _23110_, _23107_);
  and (_23113_, _23112_, _06828_);
  and (_23114_, _23039_, _03790_);
  and (_23115_, _23114_, _23108_);
  or (_23116_, _23115_, _03624_);
  or (_23117_, _23116_, _23113_);
  nor (_23118_, _13346_, _09557_);
  or (_23119_, _23032_, _07795_);
  or (_23120_, _23119_, _23118_);
  and (_23121_, _23120_, _07793_);
  and (_23122_, _23121_, _23117_);
  nor (_23123_, _13352_, _09557_);
  or (_23124_, _23123_, _23032_);
  and (_23125_, _23124_, _03785_);
  or (_23126_, _23125_, _03815_);
  or (_23127_, _23126_, _23122_);
  or (_23128_, _23036_, _04246_);
  and (_23129_, _23128_, _03823_);
  and (_23130_, _23129_, _23127_);
  and (_23131_, _23062_, _03453_);
  or (_23134_, _23131_, _03447_);
  or (_23135_, _23134_, _23130_);
  and (_23136_, _13402_, _05239_);
  or (_23137_, _23032_, _03514_);
  or (_23138_, _23137_, _23136_);
  and (_23139_, _23138_, _43000_);
  and (_23140_, _23139_, _23135_);
  nor (_23141_, _43000_, _23031_);
  or (_23142_, _23141_, rst);
  or (_43567_, _23142_, _23140_);
  and (_23144_, _43004_, \oc8051_golden_model_1.PSW [0]);
  not (_23145_, _15783_);
  nor (_23146_, _16424_, _23145_);
  and (_23147_, _16424_, _23145_);
  nor (_23148_, _23147_, _23146_);
  nor (_23149_, _23148_, _17075_);
  and (_23150_, _23148_, _17075_);
  nor (_23151_, _23150_, _23149_);
  not (_23152_, _23151_);
  nor (_23153_, _15460_, _14988_);
  and (_23154_, _15460_, _14988_);
  nor (_23155_, _23154_, _23153_);
  and (_23156_, _23155_, _16105_);
  nor (_23157_, _23155_, _16105_);
  nor (_23158_, _23157_, _23156_);
  and (_23159_, _23158_, _16761_);
  nor (_23160_, _23158_, _16761_);
  or (_23161_, _23160_, _23159_);
  and (_23162_, _23161_, _08801_);
  nor (_23163_, _23161_, _08801_);
  or (_23166_, _23163_, _23162_);
  nand (_23167_, _23166_, _23152_);
  or (_23168_, _23166_, _23152_);
  and (_23169_, _23168_, _03447_);
  and (_23170_, _23169_, _23167_);
  not (_23171_, _15529_);
  nor (_23172_, _15263_, _14957_);
  and (_23173_, _15263_, _14957_);
  nor (_23174_, _23173_, _23172_);
  nor (_23175_, _23174_, _23171_);
  and (_23177_, _23174_, _23171_);
  or (_23178_, _23177_, _23175_);
  and (_23179_, _23178_, _15888_);
  nor (_23180_, _23178_, _15888_);
  or (_23181_, _23180_, _23179_);
  and (_23182_, _23181_, _16199_);
  nor (_23183_, _23181_, _16199_);
  or (_23184_, _23183_, _23182_);
  and (_23185_, _23184_, _16529_);
  nor (_23186_, _23184_, _16529_);
  or (_23187_, _23186_, _23185_);
  and (_23188_, _23187_, _16862_);
  nor (_23189_, _23187_, _16862_);
  or (_23190_, _23189_, _23188_);
  and (_23191_, _23190_, _08140_);
  nor (_23192_, _23190_, _08140_);
  or (_23193_, _23192_, _23191_);
  and (_23194_, _23193_, _03453_);
  nor (_23195_, _07525_, _07524_);
  nor (_23196_, _23195_, _07433_);
  and (_23199_, _23195_, _07433_);
  nor (_23200_, _23199_, _23196_);
  nor (_23201_, _07449_, _07448_);
  nor (_23202_, _23201_, _15450_);
  and (_23203_, _23201_, _15450_);
  nor (_23204_, _23203_, _23202_);
  and (_23205_, _23204_, _23200_);
  nor (_23206_, _23204_, _23200_);
  nor (_23207_, _23206_, _23205_);
  or (_23208_, _23207_, _06075_);
  nand (_23210_, _23207_, _06075_);
  and (_23211_, _23210_, _23208_);
  nor (_23212_, _03628_, _03203_);
  and (_23213_, _23212_, _08733_);
  nor (_23214_, _03972_, _03515_);
  and (_23215_, _23214_, _23213_);
  nor (_23216_, _04803_, _03491_);
  and (_23217_, _23216_, _06409_);
  and (_23218_, _23217_, _23215_);
  or (_23219_, _23218_, _23211_);
  nor (_23221_, _15279_, _15278_);
  nor (_23222_, _15503_, \oc8051_golden_model_1.ACC [3]);
  and (_23223_, _15503_, \oc8051_golden_model_1.ACC [3]);
  nor (_23224_, _23223_, _23222_);
  nor (_23225_, _23201_, \oc8051_golden_model_1.ACC [6]);
  and (_23226_, _23201_, \oc8051_golden_model_1.ACC [6]);
  nor (_23227_, _23226_, _23225_);
  and (_23228_, _23227_, _23224_);
  nor (_23229_, _23227_, _23224_);
  nor (_23230_, _23229_, _23228_);
  nor (_23232_, _23230_, _23221_);
  and (_23233_, _23230_, _23221_);
  or (_23234_, _23233_, _23232_);
  and (_23235_, _23234_, _08587_);
  not (_23236_, _06377_);
  nor (_23237_, _12332_, _12003_);
  and (_23238_, _12332_, _12003_);
  nor (_23239_, _23238_, _23237_);
  and (_23240_, _23239_, _12538_);
  nor (_23241_, _23239_, _12538_);
  or (_23243_, _23241_, _23240_);
  nand (_23244_, _23243_, _12738_);
  or (_23245_, _23243_, _12738_);
  and (_23246_, _23245_, _23244_);
  nor (_23247_, _13146_, _12816_);
  and (_23248_, _13146_, _12816_);
  nor (_23249_, _23248_, _23247_);
  nor (_23250_, _23249_, _13352_);
  and (_23251_, _23249_, _13352_);
  nor (_23252_, _23251_, _23250_);
  not (_23254_, _23252_);
  nor (_23255_, _23254_, _23246_);
  and (_23256_, _23254_, _23246_);
  nor (_23257_, _23256_, _23255_);
  nor (_23258_, _23257_, _23236_);
  and (_23259_, _23257_, _23236_);
  or (_23260_, _23259_, _23258_);
  and (_23261_, _23260_, _03783_);
  nor (_23262_, _04749_, _04722_);
  and (_23263_, _23262_, _11707_);
  or (_23265_, _23263_, _23211_);
  not (_23266_, _03613_);
  and (_23267_, _11671_, _23266_);
  and (_23268_, _23267_, _03598_);
  or (_23269_, _23268_, _23211_);
  nor (_23270_, _06787_, _06638_);
  not (_23271_, _23270_);
  nand (_23272_, _23271_, _12203_);
  or (_23273_, _23271_, _12203_);
  and (_23274_, _23273_, _23272_);
  nor (_23276_, _06789_, _06731_);
  nand (_23277_, _23276_, _06456_);
  or (_23278_, _23276_, _06456_);
  and (_23279_, _23278_, _23277_);
  and (_23280_, _23279_, _23274_);
  nor (_23281_, _23279_, _23274_);
  or (_23282_, _23281_, _23280_);
  nor (_23283_, _23282_, _06069_);
  and (_23284_, _23282_, _06069_);
  or (_23285_, _23284_, _23283_);
  or (_23287_, _23285_, _08067_);
  and (_23288_, _06772_, _05469_);
  nor (_23289_, _06772_, _05469_);
  nor (_23290_, _23289_, _23288_);
  and (_23291_, _12205_, _05777_);
  nor (_23292_, _12205_, _05777_);
  nor (_23293_, _23292_, _23291_);
  nor (_23294_, _06766_, _05836_);
  nor (_23295_, _23294_, _23293_);
  and (_23296_, _23294_, _23293_);
  nor (_23298_, _23296_, _23295_);
  or (_23299_, _23298_, _23290_);
  nand (_23300_, _23298_, _23290_);
  and (_23301_, _23300_, _23299_);
  and (_23302_, _23301_, _08079_);
  nor (_23303_, _04729_, _03981_);
  and (_23304_, _23303_, \oc8051_golden_model_1.PSW [0]);
  not (_23305_, _23303_);
  and (_23306_, _23305_, _23211_);
  or (_23307_, _23306_, _23304_);
  and (_23309_, _23307_, _08078_);
  or (_23310_, _23309_, _08066_);
  or (_23311_, _23310_, _23302_);
  and (_23312_, _06072_, _03235_);
  and (_23313_, _23312_, _23311_);
  and (_23314_, _23313_, _23287_);
  and (_23315_, _23211_, _06073_);
  or (_23316_, _23315_, _04422_);
  or (_23317_, _23316_, _23314_);
  nor (_23318_, _23227_, \oc8051_golden_model_1.ACC [7]);
  and (_23320_, _23227_, \oc8051_golden_model_1.ACC [7]);
  nor (_23321_, _23320_, _23318_);
  nor (_23322_, _23321_, _23274_);
  and (_23323_, _23321_, _23274_);
  or (_23324_, _23323_, _23322_);
  or (_23325_, _23324_, _05966_);
  and (_23326_, _23325_, _04081_);
  and (_23327_, _23326_, _23317_);
  not (_23328_, _16816_);
  not (_23329_, _14988_);
  nor (_23331_, _15232_, _23329_);
  and (_23332_, _15232_, _23329_);
  nor (_23333_, _23332_, _23331_);
  and (_23334_, _23333_, _15497_);
  nor (_23335_, _23333_, _15497_);
  nor (_23336_, _23335_, _23334_);
  and (_23337_, _23336_, _16497_);
  nor (_23338_, _23336_, _16497_);
  or (_23339_, _23338_, _23337_);
  nor (_23340_, _16167_, _15855_);
  and (_23342_, _16167_, _15855_);
  nor (_23343_, _23342_, _23340_);
  and (_23344_, _23343_, _23339_);
  nor (_23345_, _23343_, _23339_);
  nor (_23346_, _23345_, _23344_);
  nor (_23347_, _23346_, _23328_);
  and (_23348_, _23346_, _23328_);
  or (_23349_, _23348_, _23347_);
  and (_23350_, _23349_, _08091_);
  nor (_23351_, _23349_, _08091_);
  or (_23352_, _23351_, _23350_);
  and (_23353_, _23352_, _03610_);
  or (_23354_, _23353_, _08089_);
  or (_23355_, _23354_, _23327_);
  and (_23356_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_23357_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_23358_, _23357_, _23356_);
  and (_23359_, _23358_, _15238_);
  nor (_23360_, _23358_, _15238_);
  nor (_23361_, _23360_, _23359_);
  nor (_23363_, _15861_, _07484_);
  and (_23364_, _15861_, _07484_);
  nor (_23365_, _23364_, _23363_);
  and (_23366_, _23365_, _23361_);
  nor (_23367_, _23365_, _23361_);
  nor (_23368_, _23367_, _23366_);
  nor (_23369_, _23368_, _16504_);
  and (_23370_, _23368_, _16504_);
  or (_23371_, _23370_, _23369_);
  nor (_23372_, _16835_, _08114_);
  and (_23374_, _16835_, _08114_);
  nor (_23375_, _23374_, _23372_);
  nor (_23376_, _23375_, _23371_);
  and (_23377_, _23375_, _23371_);
  or (_23378_, _23377_, _09882_);
  or (_23379_, _23378_, _23376_);
  and (_23380_, _23379_, _23355_);
  or (_23381_, _23380_, _09895_);
  or (_23382_, _23211_, _09896_);
  and (_23383_, _23382_, _04055_);
  and (_23384_, _23383_, _23381_);
  and (_23385_, _15245_, _14994_);
  nor (_23386_, _15245_, _14994_);
  or (_23387_, _23386_, _23385_);
  nor (_23388_, _16841_, _16179_);
  and (_23389_, _16841_, _16179_);
  nor (_23390_, _23389_, _23388_);
  nor (_23391_, _23390_, _23387_);
  and (_23392_, _23390_, _23387_);
  or (_23393_, _23392_, _23391_);
  not (_23394_, _16508_);
  nor (_23395_, _15867_, _15511_);
  and (_23396_, _15867_, _15511_);
  nor (_23397_, _23396_, _23395_);
  nor (_23398_, _23397_, _23394_);
  and (_23399_, _23397_, _23394_);
  nor (_23400_, _23399_, _23398_);
  and (_23401_, _23400_, _23393_);
  nor (_23402_, _23400_, _23393_);
  nor (_23403_, _23402_, _23401_);
  and (_23404_, _23403_, _08120_);
  nor (_23405_, _23403_, _08120_);
  or (_23406_, _23405_, _23404_);
  and (_23407_, _23406_, _03715_);
  or (_23408_, _23407_, _23384_);
  and (_23409_, _23408_, _03230_);
  and (_23410_, _23211_, _04768_);
  or (_23411_, _23410_, _23409_);
  or (_23412_, _23411_, _03723_);
  and (_23413_, _15213_, _14971_);
  nor (_23414_, _15213_, _14971_);
  nor (_23415_, _23414_, _23413_);
  and (_23416_, _23415_, _15481_);
  nor (_23417_, _23415_, _15481_);
  or (_23418_, _23417_, _23416_);
  and (_23419_, _23418_, _15818_);
  nor (_23420_, _23418_, _15818_);
  or (_23421_, _23420_, _23419_);
  and (_23422_, _23421_, _16131_);
  nor (_23423_, _23421_, _16131_);
  or (_23424_, _23423_, _23422_);
  and (_23425_, _23424_, _16461_);
  nor (_23426_, _23424_, _16461_);
  or (_23427_, _23426_, _23425_);
  and (_23428_, _23427_, _16793_);
  nor (_23429_, _23427_, _16793_);
  or (_23430_, _23429_, _23428_);
  and (_23431_, _23430_, _07910_);
  nor (_23432_, _23430_, _07910_);
  or (_23433_, _23432_, _23431_);
  or (_23435_, _23433_, _03996_);
  and (_23436_, _23435_, _08062_);
  and (_23437_, _23436_, _23412_);
  not (_23438_, _08062_);
  and (_23439_, _23301_, _23438_);
  or (_23440_, _23439_, _23437_);
  and (_23441_, _23440_, _08061_);
  and (_23442_, _23301_, _04759_);
  or (_23443_, _23442_, _04443_);
  or (_23444_, _23443_, _23441_);
  or (_23446_, _23285_, _08128_);
  and (_23447_, _23446_, _03737_);
  and (_23448_, _23447_, _23444_);
  not (_23449_, _08285_);
  nor (_23450_, _08271_, _08260_);
  and (_23451_, _08271_, _08260_);
  nor (_23452_, _23451_, _23450_);
  nor (_23453_, _23452_, _23449_);
  and (_23454_, _23452_, _23449_);
  nor (_23455_, _23454_, _23453_);
  and (_23456_, _08235_, _08218_);
  nor (_23457_, _23456_, _08517_);
  and (_23458_, _08248_, _08203_);
  nor (_23459_, _08248_, _08203_);
  or (_23460_, _23459_, _23458_);
  and (_23461_, _23460_, _23457_);
  nor (_23462_, _23460_, _23457_);
  nor (_23463_, _23462_, _23461_);
  nor (_23464_, _23463_, _23455_);
  and (_23465_, _23463_, _23455_);
  nor (_23467_, _23465_, _23464_);
  or (_23468_, _23467_, _06133_);
  nand (_23469_, _23467_, _06133_);
  and (_23470_, _23469_, _03729_);
  and (_23471_, _23470_, _23468_);
  or (_23472_, _23471_, _11668_);
  or (_23473_, _23472_, _23448_);
  or (_23474_, _23211_, _11666_);
  and (_23475_, _23474_, _03736_);
  and (_23476_, _23475_, _23473_);
  nand (_23478_, _23193_, _03714_);
  nand (_23479_, _23478_, _23268_);
  or (_23480_, _23479_, _23476_);
  nand (_23481_, _23480_, _23269_);
  not (_23482_, _03606_);
  and (_23483_, _03618_, _23482_);
  and (_23484_, _23483_, _09856_);
  and (_23485_, _11358_, _23484_);
  nand (_23486_, _23485_, _23481_);
  or (_23487_, _23485_, _23211_);
  and (_23489_, _23487_, _06840_);
  and (_23490_, _23489_, _23486_);
  nor (_23491_, _15837_, _23329_);
  and (_23492_, _15837_, _23329_);
  nor (_23493_, _23492_, _23491_);
  and (_23494_, _23493_, _16204_);
  nor (_23495_, _23493_, _16204_);
  nor (_23496_, _23495_, _23494_);
  nor (_23497_, _16868_, _08145_);
  and (_23498_, _16868_, _08145_);
  nor (_23500_, _23498_, _23497_);
  not (_23501_, _23500_);
  nor (_23502_, _23501_, _23496_);
  and (_23503_, _23501_, _23496_);
  nor (_23504_, _23503_, _23502_);
  not (_23505_, _15534_);
  and (_23506_, _23505_, _15268_);
  nor (_23507_, _23505_, _15268_);
  nor (_23508_, _23507_, _23506_);
  and (_23509_, _23508_, _16482_);
  nor (_23510_, _23508_, _16482_);
  or (_23511_, _23510_, _23509_);
  nand (_23512_, _23511_, _23504_);
  or (_23513_, _23511_, _23504_);
  and (_23514_, _23513_, _03719_);
  nand (_23515_, _23514_, _23512_);
  nand (_23516_, _23515_, _23263_);
  or (_23517_, _23516_, _23490_);
  nand (_23518_, _23517_, _23265_);
  nor (_23519_, _04463_, _04753_);
  and (_23521_, _23519_, _11353_);
  nand (_23522_, _23521_, _23518_);
  or (_23523_, _23521_, _23211_);
  and (_23524_, _23523_, _06875_);
  and (_23525_, _23524_, _23522_);
  nor (_23526_, _03753_, _11727_);
  and (_23527_, _23526_, _08848_);
  nor (_23528_, _15274_, _15020_);
  and (_23529_, _15274_, _15020_);
  or (_23530_, _23529_, _23528_);
  nor (_23532_, _23530_, _15539_);
  and (_23533_, _23530_, _15539_);
  nor (_23534_, _23533_, _23532_);
  nor (_23535_, _23534_, _15895_);
  and (_23536_, _23534_, _15895_);
  nor (_23537_, _23536_, _23535_);
  not (_23538_, _23537_);
  nor (_23539_, _23538_, _16210_);
  and (_23540_, _23538_, _16210_);
  nor (_23541_, _23540_, _23539_);
  nor (_23543_, _23541_, _16537_);
  and (_23544_, _23541_, _16537_);
  or (_23545_, _23544_, _23543_);
  and (_23546_, _23545_, _16873_);
  nor (_23547_, _23545_, _16873_);
  nor (_23548_, _23547_, _23546_);
  or (_23549_, _23548_, _08150_);
  nand (_23550_, _23548_, _08150_);
  and (_23551_, _23550_, _06869_);
  nand (_23552_, _23551_, _23549_);
  nand (_23554_, _23552_, _23527_);
  or (_23555_, _23554_, _23525_);
  or (_23556_, _23527_, _23211_);
  and (_23557_, _23556_, _09668_);
  and (_23558_, _23557_, _23555_);
  nand (_23559_, _23211_, _03752_);
  nand (_23560_, _23559_, _08059_);
  or (_23561_, _23560_, _23558_);
  not (_23562_, _08180_);
  nor (_23563_, _15285_, _08170_);
  and (_23565_, _15285_, _08170_);
  nor (_23566_, _23565_, _23563_);
  or (_23567_, _23566_, _15911_);
  nand (_23568_, _23566_, _15911_);
  and (_23569_, _23568_, _23567_);
  or (_23570_, _23569_, _15557_);
  nand (_23571_, _23569_, _15557_);
  and (_23572_, _23571_, _23570_);
  nor (_23573_, _23572_, _16229_);
  and (_23574_, _23572_, _16229_);
  nor (_23575_, _23574_, _23573_);
  nor (_23576_, _23575_, _16554_);
  and (_23577_, _23575_, _16554_);
  or (_23578_, _23577_, _23576_);
  nor (_23579_, _23578_, _16890_);
  and (_23580_, _23578_, _16890_);
  nor (_23581_, _23580_, _23579_);
  nor (_23582_, _23581_, _23562_);
  and (_23583_, _23581_, _23562_);
  or (_23584_, _23583_, _23582_);
  or (_23586_, _23584_, _08059_);
  and (_23587_, _23586_, _23561_);
  or (_23588_, _23587_, _08051_);
  nor (_23589_, _15293_, _15029_);
  and (_23590_, _15293_, _15029_);
  or (_23591_, _23590_, _23589_);
  and (_23592_, _23591_, _15573_);
  nor (_23593_, _23591_, _15573_);
  or (_23594_, _23593_, _23592_);
  nor (_23595_, _23594_, _15930_);
  and (_23597_, _23594_, _15930_);
  nor (_23598_, _23597_, _23595_);
  or (_23599_, _23598_, _16152_);
  nand (_23600_, _23598_, _16152_);
  and (_23601_, _23600_, _23599_);
  nor (_23602_, _23601_, _16576_);
  and (_23603_, _23601_, _16576_);
  or (_23604_, _23603_, _23602_);
  nor (_23605_, _23604_, _16812_);
  and (_23606_, _23604_, _16812_);
  nor (_23608_, _23606_, _23605_);
  nor (_23609_, _23608_, _08050_);
  and (_23610_, _23608_, _08050_);
  or (_23611_, _23610_, _10201_);
  or (_23612_, _23611_, _23609_);
  and (_23613_, _23612_, _03766_);
  and (_23614_, _23613_, _23588_);
  not (_23615_, _08330_);
  not (_23616_, _16134_);
  and (_23617_, _15301_, _15034_);
  nor (_23619_, _15301_, _15034_);
  nor (_23620_, _23619_, _23617_);
  nor (_23621_, _23620_, _15583_);
  and (_23622_, _23620_, _15583_);
  nor (_23623_, _23622_, _23621_);
  nor (_23624_, _23623_, _15940_);
  and (_23625_, _23623_, _15940_);
  or (_23626_, _23625_, _23624_);
  and (_23627_, _23626_, _23616_);
  nor (_23628_, _23626_, _23616_);
  nor (_23630_, _23628_, _23627_);
  and (_23631_, _23630_, _16582_);
  nor (_23632_, _23630_, _16582_);
  or (_23633_, _23632_, _23631_);
  nor (_23634_, _23633_, _16796_);
  and (_23635_, _23633_, _16796_);
  or (_23636_, _23635_, _23634_);
  and (_23637_, _23636_, _23615_);
  nor (_23638_, _23636_, _23615_);
  or (_23639_, _23638_, _23637_);
  and (_23640_, _23639_, _03761_);
  or (_23641_, _23640_, _07913_);
  or (_23642_, _23641_, _23614_);
  not (_23643_, _07974_);
  nand (_23644_, _15309_, _23643_);
  nand (_23645_, _23644_, _07975_);
  nor (_23646_, _23645_, _15599_);
  and (_23647_, _23645_, _15599_);
  nor (_23648_, _23647_, _23646_);
  nand (_23649_, _23648_, _15831_);
  or (_23651_, _23648_, _15831_);
  and (_23652_, _23651_, _23649_);
  or (_23653_, _23652_, _16248_);
  nand (_23654_, _23652_, _16248_);
  and (_23655_, _23654_, _23653_);
  nor (_23656_, _23655_, _16476_);
  and (_23657_, _23655_, _16476_);
  or (_23658_, _23657_, _23656_);
  nor (_23659_, _23658_, _16907_);
  and (_23660_, _23658_, _16907_);
  nor (_23662_, _23660_, _23659_);
  not (_23663_, _23662_);
  nor (_23664_, _23663_, _07984_);
  and (_23665_, _23663_, _07984_);
  or (_23666_, _23665_, _23664_);
  or (_23667_, _23666_, _07914_);
  and (_23668_, _23667_, _23642_);
  or (_23669_, _23668_, _07912_);
  or (_23670_, _05223_, _05210_);
  nor (_23671_, _05206_, _03550_);
  and (_23673_, _23671_, _23670_);
  nor (_23674_, _23671_, _23670_);
  or (_23675_, _23674_, _23673_);
  nor (_23676_, _05261_, _05233_);
  not (_23677_, _23676_);
  nor (_23678_, _05227_, _05219_);
  and (_23679_, _23678_, _23677_);
  nor (_23680_, _23678_, _23677_);
  nor (_23681_, _23680_, _23679_);
  nor (_23682_, _23681_, _23675_);
  and (_23684_, _23681_, _23675_);
  or (_23685_, _23684_, _23682_);
  or (_23686_, _23685_, _03248_);
  and (_23687_, _23686_, _03710_);
  and (_23688_, _23687_, _23669_);
  nor (_23689_, _03625_, _03224_);
  not (_23690_, _23689_);
  not (_23691_, _08341_);
  and (_23692_, _15317_, _15044_);
  nor (_23693_, _15317_, _15044_);
  or (_23695_, _23693_, _23692_);
  nor (_23696_, _15951_, _15607_);
  and (_23697_, _15951_, _15607_);
  nor (_23698_, _23697_, _23696_);
  nor (_23699_, _23698_, _23695_);
  and (_23700_, _23698_, _23695_);
  nor (_23701_, _23700_, _23699_);
  not (_23702_, _16916_);
  nor (_23703_, _16593_, _16257_);
  and (_23704_, _16593_, _16257_);
  nor (_23705_, _23704_, _23703_);
  nor (_23706_, _23705_, _23702_);
  and (_23707_, _23705_, _23702_);
  nor (_23708_, _23707_, _23706_);
  nor (_23709_, _23708_, _23701_);
  and (_23710_, _23708_, _23701_);
  or (_23711_, _23710_, _23709_);
  nand (_23712_, _23711_, _23691_);
  and (_23713_, _23711_, _03505_);
  or (_23714_, _23713_, _08342_);
  and (_23716_, _23714_, _23712_);
  or (_23717_, _23716_, _23690_);
  or (_23718_, _23717_, _23688_);
  or (_23719_, _23689_, _23211_);
  and (_23720_, _23719_, _23718_);
  or (_23721_, _23720_, _10658_);
  and (_23722_, _23433_, _06834_);
  or (_23723_, _23722_, _06838_);
  and (_23724_, _23723_, _23721_);
  and (_23725_, _23433_, _06833_);
  or (_23727_, _23725_, _04481_);
  or (_23728_, _23727_, _23724_);
  and (_23729_, _15324_, _15051_);
  nor (_23730_, _15324_, _15051_);
  nor (_23731_, _23730_, _23729_);
  not (_23732_, _15959_);
  and (_23733_, _23732_, _15614_);
  nor (_23734_, _23732_, _15614_);
  nor (_23735_, _23734_, _23733_);
  nor (_23736_, _23735_, _23731_);
  and (_23738_, _23735_, _23731_);
  or (_23739_, _23738_, _23736_);
  not (_23740_, _16600_);
  and (_23741_, _23740_, _16265_);
  nor (_23742_, _23740_, _16265_);
  nor (_23743_, _23742_, _23741_);
  nand (_23744_, _23743_, _16924_);
  or (_23745_, _23743_, _16924_);
  and (_23746_, _23745_, _23744_);
  or (_23747_, _23746_, _23739_);
  nand (_23749_, _23746_, _23739_);
  and (_23750_, _23749_, _23747_);
  nor (_23751_, _23750_, _08348_);
  and (_23752_, _23750_, _08348_);
  or (_23753_, _23752_, _07400_);
  or (_23754_, _23753_, _23751_);
  and (_23755_, _23754_, _03589_);
  and (_23756_, _23755_, _23728_);
  and (_23757_, _15329_, _15056_);
  nor (_23758_, _15329_, _15056_);
  nor (_23760_, _23758_, _23757_);
  and (_23761_, _23760_, _15619_);
  nor (_23762_, _23760_, _15619_);
  or (_23763_, _23762_, _23761_);
  and (_23764_, _23763_, _15965_);
  nor (_23765_, _23763_, _15965_);
  or (_23766_, _23765_, _23764_);
  not (_23767_, _16606_);
  and (_23768_, _23767_, _16270_);
  nor (_23769_, _23767_, _16270_);
  nor (_23770_, _23769_, _23768_);
  not (_23771_, _16929_);
  and (_23772_, _23771_, _08353_);
  nor (_23773_, _23771_, _08353_);
  nor (_23774_, _23773_, _23772_);
  or (_23775_, _23774_, _23770_);
  nand (_23776_, _23774_, _23770_);
  and (_23777_, _23776_, _23775_);
  or (_23778_, _23777_, _23766_);
  nand (_23779_, _23777_, _23766_);
  and (_23781_, _23779_, _03222_);
  and (_23782_, _23781_, _23778_);
  or (_23783_, _23782_, _07405_);
  or (_23784_, _23783_, _23756_);
  and (_23785_, _07463_, _16935_);
  nor (_23786_, _07463_, _16935_);
  nor (_23787_, _23786_, _23785_);
  nor (_23788_, _07604_, _07547_);
  and (_23789_, _07604_, _07547_);
  nor (_23790_, _23789_, _23788_);
  nor (_23792_, _23790_, _07493_);
  and (_23793_, _23790_, _07493_);
  nor (_23794_, _23793_, _23792_);
  nor (_23795_, _23794_, _23787_);
  and (_23796_, _23794_, _23787_);
  nor (_23797_, _23796_, _23795_);
  not (_23798_, _23797_);
  nor (_23799_, _07674_, _07424_);
  and (_23800_, _07674_, _07424_);
  nor (_23801_, _23800_, _23799_);
  nor (_23803_, _23801_, _23798_);
  and (_23804_, _23801_, _23798_);
  nor (_23805_, _23804_, _23803_);
  and (_23806_, _23805_, _07760_);
  nor (_23807_, _23805_, _07760_);
  or (_23808_, _23807_, _07411_);
  or (_23809_, _23808_, _23806_);
  and (_23810_, _23809_, _03217_);
  and (_23811_, _23810_, _23784_);
  nand (_23812_, _23685_, _03216_);
  nor (_23814_, _11764_, _04754_);
  and (_23815_, _23814_, _11760_);
  and (_23816_, _23815_, _04734_);
  and (_23817_, _05889_, _04733_);
  and (_23818_, _23817_, _23816_);
  nand (_23819_, _23818_, _23812_);
  or (_23820_, _23819_, _23811_);
  or (_23821_, _23818_, _23211_);
  and (_23822_, _23821_, _05886_);
  and (_23823_, _23822_, _23820_);
  nor (_23825_, _15339_, _14959_);
  and (_23826_, _15339_, _14959_);
  or (_23827_, _23826_, _23825_);
  nor (_23828_, _15976_, _15630_);
  and (_23829_, _15976_, _15630_);
  nor (_23830_, _23829_, _23828_);
  nor (_23831_, _23830_, _23827_);
  and (_23832_, _23830_, _23827_);
  or (_23833_, _23832_, _23831_);
  nor (_23834_, _16445_, _16281_);
  and (_23835_, _16445_, _16281_);
  nor (_23836_, _23835_, _23834_);
  and (_23837_, _23836_, _16780_);
  nor (_23838_, _23836_, _16780_);
  nor (_23839_, _23838_, _23837_);
  nor (_23840_, _23839_, _23833_);
  and (_23841_, _23839_, _23833_);
  nor (_23842_, _23841_, _23840_);
  and (_23843_, _23842_, _08366_);
  nor (_23844_, _23842_, _08366_);
  or (_23846_, _23844_, _23843_);
  and (_23847_, _23846_, _03601_);
  or (_23848_, _23847_, _23823_);
  and (_23849_, _23848_, _08364_);
  nand (_23850_, _23685_, _08363_);
  and (_23851_, _11815_, _11348_);
  and (_23852_, _23851_, _11820_);
  nand (_23853_, _23852_, _23850_);
  or (_23854_, _23853_, _23849_);
  or (_23855_, _23852_, _23211_);
  and (_23857_, _23855_, _11343_);
  and (_23858_, _23857_, _23854_);
  nor (_23859_, _15799_, _08676_);
  and (_23860_, _15799_, _08676_);
  nor (_23861_, _23860_, _23859_);
  and (_23862_, _15072_, _08680_);
  nor (_23863_, _23862_, _15550_);
  nor (_23864_, _23863_, _23861_);
  and (_23865_, _23863_, _23861_);
  nor (_23866_, _23865_, _23864_);
  nor (_23868_, _16453_, _08669_);
  and (_23869_, _16453_, _08669_);
  nor (_23870_, _23869_, _23868_);
  nor (_23871_, _23870_, _23866_);
  and (_23872_, _23870_, _23866_);
  nor (_23873_, _23872_, _23871_);
  not (_23874_, _23873_);
  and (_23875_, _08664_, _08376_);
  nor (_23876_, _08664_, _08376_);
  nor (_23877_, _23876_, _23875_);
  nor (_23879_, _23877_, _23874_);
  and (_23880_, _23877_, _23874_);
  or (_23881_, _23880_, _23879_);
  and (_23882_, _23881_, _11344_);
  or (_23883_, _23882_, _08392_);
  or (_23884_, _23883_, _23858_);
  nor (_23885_, _15921_, _08640_);
  and (_23886_, _15921_, _08640_);
  nor (_23887_, _23886_, _23885_);
  and (_23888_, _15083_, _08644_);
  nor (_23890_, _23888_, _15568_);
  nor (_23891_, _23890_, _23887_);
  and (_23892_, _23890_, _23887_);
  nor (_23893_, _23892_, _23891_);
  nor (_23894_, _08630_, _08634_);
  and (_23895_, _08630_, _08634_);
  nor (_23896_, _23895_, _23894_);
  nor (_23897_, _23896_, _23893_);
  and (_23898_, _23896_, _23893_);
  nor (_23899_, _23898_, _23897_);
  nor (_23900_, _23899_, _08627_);
  and (_23901_, _23899_, _08627_);
  or (_23902_, _23901_, _23900_);
  and (_23903_, _23902_, _08400_);
  nor (_23904_, _23902_, _08400_);
  or (_23905_, _23904_, _23903_);
  or (_23906_, _23905_, _08393_);
  and (_23907_, _23906_, _03779_);
  and (_23908_, _23907_, _23884_);
  nor (_23909_, _12739_, _12539_);
  and (_23911_, _12739_, _12539_);
  nor (_23912_, _23911_, _23909_);
  nor (_23913_, _12333_, _12128_);
  and (_23914_, _12333_, _12128_);
  nor (_23915_, _23914_, _23913_);
  not (_23916_, _23915_);
  and (_23917_, _23916_, _23912_);
  nor (_23918_, _23916_, _23912_);
  nor (_23919_, _23918_, _23917_);
  or (_23920_, _23919_, _12817_);
  nand (_23922_, _23919_, _12817_);
  and (_23923_, _23922_, _23920_);
  or (_23924_, _23923_, _13147_);
  nand (_23925_, _23923_, _13147_);
  and (_23926_, _23925_, _23924_);
  or (_23927_, _23926_, _13353_);
  nand (_23928_, _23926_, _13353_);
  and (_23929_, _23928_, _23927_);
  nor (_23930_, _23929_, _06378_);
  and (_23931_, _23929_, _06378_);
  or (_23933_, _23931_, _23930_);
  and (_23934_, _23933_, _03778_);
  or (_23935_, _23934_, _07904_);
  or (_23936_, _23935_, _23908_);
  and (_23937_, _16734_, _08737_);
  and (_23938_, _10026_, _08738_);
  nor (_23939_, _23938_, _23937_);
  not (_23940_, _10058_);
  nor (_23941_, _08753_, _23940_);
  and (_23942_, _08753_, _23940_);
  nor (_23944_, _23942_, _23941_);
  and (_23945_, _10030_, _08748_);
  nor (_23946_, _23945_, _10031_);
  and (_23947_, _23946_, _23944_);
  nor (_23948_, _23946_, _23944_);
  nor (_23949_, _23948_, _23947_);
  nor (_23950_, _23949_, _08743_);
  and (_23951_, _23949_, _08743_);
  or (_23952_, _23951_, _23950_);
  nor (_23953_, _23952_, _23939_);
  and (_23955_, _23952_, _23939_);
  nor (_23956_, _23955_, _23953_);
  nand (_23957_, _23956_, _08407_);
  or (_23958_, _23956_, _08407_);
  and (_23959_, _23958_, _23957_);
  or (_23960_, _23959_, _07905_);
  and (_23961_, _23960_, _07766_);
  and (_23962_, _23961_, _23936_);
  and (_23963_, _15209_, _14965_);
  nor (_23964_, _15209_, _14965_);
  nor (_23966_, _23964_, _23963_);
  and (_23967_, _23966_, _15474_);
  nor (_23968_, _23966_, _15474_);
  or (_23969_, _23968_, _23967_);
  nand (_23970_, _23969_, _15813_);
  or (_23971_, _23969_, _15813_);
  and (_23972_, _23971_, _23970_);
  nor (_23973_, _16784_, _16450_);
  and (_23974_, _16784_, _16450_);
  nor (_23975_, _23974_, _23973_);
  not (_23977_, _16124_);
  and (_23978_, _23977_, _07902_);
  nor (_23979_, _23977_, _07902_);
  nor (_23980_, _23979_, _23978_);
  nor (_23981_, _23980_, _23975_);
  and (_23982_, _23980_, _23975_);
  nor (_23983_, _23982_, _23981_);
  nand (_23984_, _23983_, _23972_);
  or (_23985_, _23983_, _23972_);
  and (_23986_, _23985_, _03600_);
  and (_23988_, _23986_, _23984_);
  or (_23989_, _23988_, _23962_);
  and (_23990_, _23989_, _07778_);
  nor (_23991_, _11841_, _03182_);
  nand (_23992_, _23211_, _03780_);
  or (_23993_, _23992_, _05254_);
  nand (_23994_, _23993_, _23991_);
  or (_23995_, _23994_, _23990_);
  or (_23996_, _23991_, _23211_);
  and (_23997_, _23996_, _08414_);
  and (_23999_, _23997_, _08416_);
  and (_24000_, _23999_, _23995_);
  or (_24001_, _08681_, _08678_);
  nand (_24002_, _08681_, _08678_);
  and (_24003_, _24002_, _24001_);
  nor (_24004_, _08672_, _08674_);
  and (_24005_, _08672_, _08674_);
  nor (_24006_, _24005_, _24004_);
  and (_24007_, _24006_, _24003_);
  nor (_24008_, _24006_, _24003_);
  nor (_24010_, _24008_, _24007_);
  and (_24011_, _08662_, _08375_);
  or (_24012_, _24011_, _10329_);
  nor (_24013_, _08665_, _08667_);
  and (_24014_, _08665_, _08667_);
  nor (_24015_, _24014_, _24013_);
  not (_24016_, _24015_);
  and (_24017_, _24016_, _24012_);
  nor (_24018_, _24016_, _24012_);
  nor (_24019_, _24018_, _24017_);
  nor (_24021_, _24019_, _24010_);
  and (_24022_, _24019_, _24010_);
  or (_24023_, _24022_, _24021_);
  and (_24024_, _24023_, _08421_);
  or (_24025_, _24024_, _08420_);
  or (_24026_, _24025_, _24000_);
  not (_24027_, _08638_);
  or (_24028_, _08645_, _08642_);
  nand (_24029_, _08645_, _08642_);
  and (_24030_, _24029_, _24028_);
  nand (_24032_, _24030_, _24027_);
  or (_24033_, _24030_, _24027_);
  and (_24034_, _24033_, _24032_);
  nor (_24035_, _24034_, _08635_);
  and (_24036_, _24034_, _08635_);
  or (_24037_, _24036_, _24035_);
  not (_24038_, _08628_);
  nor (_24039_, _08632_, _08625_);
  and (_24040_, _08632_, _08625_);
  nor (_24041_, _24040_, _24039_);
  nor (_24043_, _24041_, _24038_);
  and (_24044_, _24041_, _24038_);
  nor (_24045_, _24044_, _24043_);
  nor (_24046_, _24045_, _24037_);
  and (_24047_, _24045_, _24037_);
  nor (_24048_, _24047_, _24046_);
  and (_24049_, _24048_, _08399_);
  nor (_24050_, _24048_, _08399_);
  or (_24051_, _24050_, _24049_);
  or (_24052_, _24051_, _08425_);
  and (_24054_, _24052_, _03789_);
  and (_24055_, _24054_, _24026_);
  nor (_24056_, _12331_, _12005_);
  and (_24057_, _12331_, _12005_);
  nor (_24058_, _24057_, _24056_);
  not (_24059_, _24058_);
  not (_24060_, _12737_);
  and (_24061_, _24060_, _12537_);
  nor (_24062_, _24060_, _12537_);
  nor (_24063_, _24062_, _24061_);
  nor (_24065_, _24063_, _24059_);
  and (_24066_, _24063_, _24059_);
  nor (_24067_, _24066_, _24065_);
  not (_24068_, _13351_);
  nor (_24069_, _13145_, _12815_);
  and (_24070_, _13145_, _12815_);
  nor (_24071_, _24070_, _24069_);
  nor (_24072_, _24071_, _24068_);
  and (_24073_, _24071_, _24068_);
  nor (_24074_, _24073_, _24072_);
  not (_24076_, _24074_);
  nor (_24077_, _24076_, _24067_);
  and (_24078_, _24076_, _24067_);
  nor (_24079_, _24078_, _24077_);
  or (_24080_, _24079_, _06376_);
  nand (_24081_, _24079_, _06376_);
  and (_24082_, _24081_, _03788_);
  and (_24083_, _24082_, _24080_);
  or (_24084_, _24083_, _08429_);
  or (_24085_, _24084_, _24055_);
  not (_24087_, _08741_);
  or (_24088_, _08750_, _08751_);
  nand (_24089_, _08750_, _08751_);
  and (_24090_, _24089_, _24088_);
  not (_24091_, _08744_);
  and (_24092_, _24091_, _08746_);
  nor (_24093_, _24091_, _08746_);
  nor (_24094_, _24093_, _24092_);
  not (_24095_, _24094_);
  and (_24096_, _24095_, _24090_);
  nor (_24098_, _24095_, _24090_);
  nor (_24099_, _24098_, _24096_);
  nand (_24100_, _24099_, _24087_);
  or (_24101_, _24099_, _24087_);
  and (_24102_, _24101_, _24100_);
  or (_24103_, _24102_, _08739_);
  nand (_24104_, _24102_, _08739_);
  and (_24105_, _24104_, _24103_);
  or (_24106_, _24105_, _08735_);
  nand (_24107_, _24105_, _08735_);
  and (_24109_, _24107_, _24106_);
  nor (_24110_, _24109_, _08405_);
  and (_24111_, _24109_, _08405_);
  or (_24112_, _24111_, _24110_);
  or (_24113_, _24112_, _08435_);
  and (_24114_, _24113_, _07777_);
  and (_24115_, _24114_, _24085_);
  and (_24116_, _11338_, _10753_);
  nor (_24117_, _15687_, _14960_);
  and (_24118_, _15687_, _14960_);
  nor (_24120_, _24118_, _24117_);
  nor (_24121_, _16781_, _16333_);
  and (_24122_, _16781_, _16333_);
  nor (_24123_, _24122_, _24121_);
  and (_24124_, _24123_, _24120_);
  nor (_24125_, _24123_, _24120_);
  nor (_24126_, _24125_, _24124_);
  nor (_24127_, _16447_, _16017_);
  and (_24128_, _16447_, _16017_);
  nor (_24129_, _24128_, _24127_);
  nor (_24131_, _15206_, _08439_);
  and (_24132_, _15206_, _08439_);
  nor (_24133_, _24132_, _24131_);
  and (_24134_, _24133_, _24129_);
  nor (_24135_, _24133_, _24129_);
  nor (_24136_, _24135_, _24134_);
  not (_24137_, _24136_);
  nand (_24138_, _24137_, _24126_);
  or (_24139_, _24137_, _24126_);
  and (_24140_, _24139_, _03622_);
  nand (_24142_, _24140_, _24138_);
  nand (_24143_, _24142_, _24116_);
  or (_24144_, _24143_, _24115_);
  or (_24145_, _23211_, _24116_);
  and (_24146_, _24145_, _08447_);
  and (_24147_, _24146_, _24144_);
  nor (_24148_, _15071_, _08679_);
  and (_24149_, _15071_, _08679_);
  nor (_24150_, _24149_, _24148_);
  and (_24151_, _24150_, _08675_);
  nor (_24153_, _24150_, _08675_);
  or (_24154_, _24153_, _24151_);
  nand (_24155_, _24154_, _08673_);
  or (_24156_, _24154_, _08673_);
  and (_24157_, _24156_, _24155_);
  not (_24158_, _08666_);
  nor (_24159_, _08668_, _08663_);
  and (_24160_, _08668_, _08663_);
  nor (_24161_, _24160_, _24159_);
  nor (_24162_, _24161_, _24158_);
  and (_24164_, _24161_, _24158_);
  nor (_24165_, _24164_, _24162_);
  and (_24166_, _24165_, _24157_);
  nor (_24167_, _24165_, _24157_);
  or (_24168_, _24167_, _24166_);
  and (_24169_, _24168_, _08374_);
  nor (_24170_, _24168_, _08374_);
  or (_24171_, _24170_, _24169_);
  and (_24172_, _24171_, _08446_);
  or (_24173_, _24172_, _08450_);
  or (_24175_, _24173_, _24147_);
  not (_24176_, _08398_);
  nor (_24177_, _15082_, _08643_);
  and (_24178_, _15082_, _08643_);
  nor (_24179_, _24178_, _24177_);
  and (_24180_, _24179_, _08639_);
  nor (_24181_, _24179_, _08639_);
  or (_24182_, _24181_, _24180_);
  nand (_24183_, _24182_, _08637_);
  or (_24184_, _24182_, _08637_);
  and (_24187_, _24184_, _24183_);
  nor (_24188_, _08633_, _08626_);
  and (_24189_, _08633_, _08626_);
  nor (_24190_, _24189_, _24188_);
  and (_24191_, _24190_, _08629_);
  nor (_24192_, _24190_, _08629_);
  nor (_24193_, _24192_, _24191_);
  and (_24194_, _24193_, _24187_);
  nor (_24195_, _24193_, _24187_);
  or (_24196_, _24195_, _24194_);
  nor (_24199_, _24196_, _24176_);
  and (_24200_, _24196_, _24176_);
  nor (_24201_, _24200_, _24199_);
  nand (_24202_, _24201_, _08450_);
  and (_24203_, _24202_, _03784_);
  and (_24204_, _24203_, _24175_);
  or (_24205_, _24204_, _23261_);
  and (_24206_, _24205_, _08461_);
  nor (_24207_, _08752_, _10057_);
  and (_24208_, _08752_, _10057_);
  nor (_24211_, _24208_, _24207_);
  not (_24212_, _24211_);
  not (_24213_, _08745_);
  and (_24214_, _24213_, _08747_);
  nor (_24215_, _24213_, _08747_);
  nor (_24216_, _24215_, _24214_);
  nor (_24217_, _24216_, _24212_);
  and (_24218_, _24216_, _24212_);
  nor (_24219_, _24218_, _24217_);
  and (_24220_, _24219_, _08742_);
  nor (_24223_, _24219_, _08742_);
  or (_24224_, _24223_, _24220_);
  and (_24225_, _24224_, _08740_);
  nor (_24226_, _24224_, _08740_);
  or (_24227_, _24226_, _24225_);
  and (_24228_, _24227_, _08736_);
  nor (_24229_, _24227_, _08736_);
  or (_24230_, _24229_, _24228_);
  and (_24231_, _24230_, _08406_);
  nor (_24232_, _24230_, _08406_);
  or (_24235_, _24232_, _24231_);
  and (_24236_, _24235_, _08458_);
  or (_24237_, _24236_, _24206_);
  and (_24238_, _24237_, _07795_);
  and (_24239_, _11881_, _11877_);
  nor (_24240_, _15401_, _15144_);
  and (_24241_, _15401_, _15144_);
  or (_24242_, _24241_, _24240_);
  nor (_24243_, _16037_, _15710_);
  and (_24244_, _16037_, _15710_);
  nor (_24247_, _24244_, _24243_);
  nor (_24248_, _24247_, _24242_);
  and (_24249_, _24247_, _24242_);
  nor (_24250_, _24249_, _24248_);
  not (_24251_, _24250_);
  nor (_24252_, _17004_, _16442_);
  and (_24253_, _17004_, _16442_);
  nor (_24254_, _24253_, _24252_);
  not (_24255_, _16352_);
  and (_24256_, _24255_, _08470_);
  nor (_24259_, _24255_, _08470_);
  nor (_24260_, _24259_, _24256_);
  nor (_24261_, _24260_, _24254_);
  and (_24262_, _24260_, _24254_);
  nor (_24263_, _24262_, _24261_);
  nand (_24264_, _24263_, _24251_);
  or (_24265_, _24263_, _24251_);
  and (_24266_, _24265_, _03624_);
  nand (_24267_, _24266_, _24264_);
  nand (_24268_, _24267_, _24239_);
  or (_24270_, _24268_, _24238_);
  or (_24271_, _23211_, _24239_);
  and (_24272_, _24271_, _07898_);
  and (_24273_, _24272_, _24270_);
  not (_24274_, _15805_);
  nor (_24275_, _15406_, _08170_);
  and (_24276_, _15406_, _08170_);
  or (_24277_, _24276_, _24275_);
  nor (_24278_, _24277_, _15716_);
  and (_24279_, _24277_, _15716_);
  nor (_24281_, _24279_, _24278_);
  and (_24282_, _24281_, _24274_);
  nor (_24283_, _24281_, _24274_);
  nor (_24284_, _24283_, _24282_);
  nor (_24285_, _24284_, _16357_);
  and (_24286_, _24284_, _16357_);
  or (_24287_, _24286_, _24285_);
  and (_24288_, _24287_, _16684_);
  nor (_24289_, _24287_, _16684_);
  nor (_24290_, _24289_, _24288_);
  nor (_24292_, _24290_, _17010_);
  and (_24293_, _24290_, _17010_);
  or (_24294_, _24293_, _24292_);
  nor (_24295_, _24294_, _07890_);
  and (_24296_, _24294_, _07890_);
  or (_24297_, _24296_, _24295_);
  and (_24298_, _24297_, _08468_);
  or (_24299_, _24298_, _08475_);
  or (_24300_, _24299_, _24273_);
  not (_24301_, _16690_);
  not (_24303_, _16045_);
  nor (_24304_, _15411_, _15029_);
  and (_24305_, _15411_, _15029_);
  or (_24306_, _24305_, _24304_);
  nor (_24307_, _24306_, _15721_);
  and (_24308_, _24306_, _15721_);
  nor (_24309_, _24308_, _24307_);
  and (_24310_, _24309_, _24303_);
  nor (_24311_, _24309_, _24303_);
  nor (_24312_, _24311_, _24310_);
  nor (_24314_, _24312_, _16363_);
  and (_24315_, _24312_, _16363_);
  or (_24316_, _24315_, _24314_);
  nor (_24317_, _24316_, _24301_);
  and (_24318_, _24316_, _24301_);
  nor (_24319_, _24318_, _24317_);
  and (_24320_, _24319_, _17015_);
  nor (_24321_, _24319_, _17015_);
  or (_24322_, _24321_, _24320_);
  not (_24323_, _24322_);
  nor (_24325_, _24323_, _08502_);
  and (_24326_, _24323_, _08502_);
  or (_24327_, _24326_, _24325_);
  or (_24328_, _24327_, _08477_);
  and (_24329_, _24328_, _03777_);
  and (_24330_, _24329_, _24300_);
  nor (_24331_, _15416_, _15034_);
  and (_24332_, _15416_, _15034_);
  or (_24333_, _24332_, _24331_);
  nor (_24334_, _24333_, _15727_);
  and (_24336_, _24333_, _15727_);
  nor (_24337_, _24336_, _24334_);
  nor (_24338_, _24337_, _16050_);
  and (_24339_, _24337_, _16050_);
  or (_24340_, _24339_, _24338_);
  nor (_24341_, _24340_, _16368_);
  and (_24342_, _24340_, _16368_);
  or (_24343_, _24342_, _24341_);
  nor (_24344_, _24343_, _16695_);
  and (_24345_, _24343_, _16695_);
  or (_24347_, _24345_, _24344_);
  and (_24348_, _24347_, _17021_);
  nor (_24349_, _24347_, _17021_);
  or (_24350_, _24349_, _24348_);
  or (_24351_, _24350_, _08583_);
  nand (_24352_, _24350_, _08583_);
  and (_24353_, _24352_, _03776_);
  and (_24354_, _24353_, _24351_);
  or (_24355_, _24354_, _08506_);
  or (_24356_, _24355_, _24330_);
  not (_24358_, _08613_);
  and (_24359_, _15421_, _07974_);
  and (_24360_, _23643_, _07972_);
  nor (_24361_, _24360_, _24359_);
  nor (_24362_, _24361_, _15732_);
  and (_24363_, _24361_, _15732_);
  nor (_24364_, _24363_, _24362_);
  or (_24365_, _24364_, _16056_);
  nand (_24366_, _24364_, _16056_);
  and (_24367_, _24366_, _24365_);
  nor (_24369_, _24367_, _16374_);
  and (_24370_, _24367_, _16374_);
  nor (_24371_, _24370_, _24369_);
  nor (_24372_, _24371_, _16701_);
  and (_24373_, _24371_, _16701_);
  or (_24374_, _24373_, _24372_);
  and (_24375_, _24374_, _17026_);
  nor (_24376_, _24374_, _17026_);
  nor (_24377_, _24376_, _24375_);
  nor (_24378_, _24377_, _24358_);
  and (_24380_, _24377_, _24358_);
  or (_24381_, _24380_, _24378_);
  or (_24382_, _24381_, _08589_);
  and (_24383_, _24382_, _08588_);
  and (_24384_, _24383_, _24356_);
  or (_24385_, _24384_, _23235_);
  and (_24386_, _10774_, _11903_);
  and (_24387_, _24386_, _24385_);
  not (_24388_, _24386_);
  nand (_24389_, _24388_, _23211_);
  nand (_24391_, _24389_, _16706_);
  or (_24392_, _24391_, _24387_);
  not (_24393_, _15071_);
  and (_24394_, _24393_, _08680_);
  nor (_24395_, _24393_, _08680_);
  nor (_24396_, _24395_, _24394_);
  and (_24397_, _24396_, _15741_);
  nor (_24398_, _24396_, _15741_);
  nor (_24399_, _24398_, _24397_);
  and (_24400_, _24399_, _15802_);
  nor (_24402_, _24399_, _15802_);
  or (_24403_, _24402_, _24400_);
  and (_24404_, _24403_, _16383_);
  nor (_24405_, _24403_, _16383_);
  nor (_24406_, _24405_, _24404_);
  nor (_24407_, _24406_, _16715_);
  and (_24408_, _24406_, _16715_);
  nor (_24409_, _24408_, _24407_);
  and (_24410_, _24409_, _17035_);
  nor (_24411_, _24409_, _17035_);
  or (_24413_, _24411_, _24410_);
  nor (_24414_, _24413_, _08696_);
  and (_24415_, _24413_, _08696_);
  or (_24416_, _24415_, _24414_);
  or (_24417_, _24416_, _16706_);
  and (_24418_, _24417_, _16712_);
  and (_24419_, _24418_, _24392_);
  and (_24420_, _24416_, _16710_);
  or (_24421_, _24420_, _08620_);
  or (_24422_, _24421_, _24419_);
  not (_24424_, _08660_);
  and (_24425_, _15082_, _08644_);
  nor (_24426_, _15082_, _08644_);
  or (_24427_, _24426_, _24425_);
  and (_24428_, _24427_, _15747_);
  nor (_24429_, _24427_, _15747_);
  nor (_24430_, _24429_, _24428_);
  nor (_24431_, _24430_, _16068_);
  and (_24432_, _24430_, _16068_);
  or (_24433_, _24432_, _24431_);
  nor (_24435_, _24433_, _16388_);
  and (_24436_, _24433_, _16388_);
  or (_24437_, _24436_, _24435_);
  and (_24438_, _24437_, _16724_);
  nor (_24439_, _24437_, _16724_);
  nor (_24440_, _24439_, _24438_);
  nor (_24441_, _24440_, _17041_);
  and (_24442_, _24440_, _17041_);
  or (_24443_, _24442_, _24441_);
  nor (_24444_, _24443_, _24424_);
  and (_24446_, _24443_, _24424_);
  or (_24447_, _24446_, _24444_);
  or (_24448_, _24447_, _08624_);
  and (_24449_, _24448_, _03518_);
  and (_24450_, _24449_, _24422_);
  nor (_24451_, _15436_, _08318_);
  and (_24452_, _15436_, _08318_);
  or (_24453_, _24452_, _24451_);
  nor (_24454_, _24453_, _15752_);
  and (_24455_, _24453_, _15752_);
  nor (_24457_, _24455_, _24454_);
  and (_24458_, _24457_, _16075_);
  nor (_24459_, _24457_, _16075_);
  nor (_24460_, _24459_, _24458_);
  and (_24461_, _24460_, _16394_);
  nor (_24462_, _24460_, _16394_);
  nor (_24463_, _24462_, _24461_);
  nor (_24464_, _24463_, _16729_);
  and (_24465_, _24463_, _16729_);
  or (_24466_, _24465_, _24464_);
  nor (_24468_, _24466_, _17046_);
  and (_24469_, _24466_, _17046_);
  or (_24470_, _24469_, _24468_);
  or (_24471_, _24470_, _08728_);
  nand (_24472_, _24470_, _08728_);
  and (_24473_, _24472_, _03517_);
  and (_24474_, _24473_, _24471_);
  or (_24475_, _24474_, _24450_);
  and (_24476_, _24475_, _08734_);
  and (_24477_, _15441_, _23940_);
  nor (_24479_, _24477_, _23941_);
  and (_24480_, _24479_, _15758_);
  nor (_24481_, _24479_, _15758_);
  nor (_24482_, _24481_, _24480_);
  nor (_24483_, _24482_, _16081_);
  and (_24484_, _24482_, _16081_);
  nor (_24485_, _24484_, _24483_);
  nor (_24486_, _24485_, _16399_);
  and (_24487_, _24485_, _16399_);
  or (_24488_, _24487_, _24486_);
  nor (_24490_, _24488_, _16737_);
  and (_24491_, _24488_, _16737_);
  or (_24492_, _24491_, _24490_);
  nor (_24493_, _24492_, _17052_);
  and (_24494_, _24492_, _17052_);
  or (_24495_, _24494_, _24493_);
  nor (_24496_, _24495_, _08768_);
  and (_24497_, _24495_, _08768_);
  or (_24498_, _24497_, _24496_);
  nand (_24499_, _24498_, _08701_);
  nand (_24501_, _24499_, _23218_);
  or (_24502_, _24501_, _24476_);
  and (_24503_, _24502_, _23219_);
  or (_24504_, _24503_, _03815_);
  or (_24505_, _23352_, _04246_);
  and (_24506_, _24505_, _08776_);
  and (_24507_, _24506_, _24504_);
  not (_24508_, _08781_);
  and (_24509_, _15503_, _24508_);
  and (_24510_, _24509_, \oc8051_golden_model_1.ACC [3]);
  nor (_24512_, _24509_, \oc8051_golden_model_1.ACC [3]);
  nor (_24513_, _24512_, _24510_);
  and (_24514_, _24513_, _16412_);
  nor (_24515_, _24513_, _16412_);
  nor (_24516_, _24515_, _24514_);
  and (_24517_, _16748_, _07433_);
  nor (_24518_, _16748_, _07433_);
  nor (_24519_, _24518_, _24517_);
  nor (_24520_, _24519_, _24516_);
  and (_24521_, _24519_, _24516_);
  or (_24523_, _24521_, _24520_);
  or (_24524_, _24523_, _08788_);
  nand (_24525_, _24523_, _08788_);
  and (_24526_, _24525_, _24524_);
  and (_24527_, _24526_, _08775_);
  or (_24528_, _24527_, _24507_);
  and (_24529_, _24528_, _10359_);
  and (_24530_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_24531_, _24530_, _08110_);
  nand (_24532_, _24531_, _23230_);
  or (_24534_, _24531_, _23230_);
  and (_24535_, _24534_, _24532_);
  nand (_24536_, _24535_, _08780_);
  nand (_24537_, _24536_, _04540_);
  or (_24538_, _24537_, _24529_);
  or (_24539_, _23211_, _04540_);
  and (_24540_, _24539_, _03823_);
  and (_24541_, _24540_, _24538_);
  or (_24542_, _24541_, _23194_);
  and (_24543_, _24542_, _11955_);
  and (_24545_, _23211_, _11956_);
  or (_24546_, _24545_, _04552_);
  or (_24547_, _24546_, _24543_);
  or (_24548_, _23211_, _06785_);
  and (_24549_, _24548_, _03514_);
  and (_24550_, _24549_, _24547_);
  or (_24551_, _24550_, _23170_);
  and (_24552_, _24551_, _08799_);
  nor (_24553_, _11975_, _03196_);
  nor (_24554_, _08805_, _03631_);
  and (_24556_, _24554_, _24553_);
  not (_24557_, _08806_);
  and (_24558_, _15503_, _24557_);
  and (_24559_, _24558_, _07578_);
  nor (_24560_, _24558_, _07578_);
  nor (_24561_, _24560_, _24559_);
  nor (_24562_, _17080_, _16430_);
  and (_24563_, _17080_, _16430_);
  or (_24564_, _24563_, _24562_);
  or (_24565_, _24564_, _24561_);
  nand (_24567_, _24564_, _24561_);
  and (_24568_, _24567_, _24565_);
  nor (_24569_, _16767_, _08813_);
  and (_24570_, _16767_, _08813_);
  nor (_24571_, _24570_, _24569_);
  not (_24572_, _24571_);
  nand (_24573_, _24572_, _24568_);
  or (_24574_, _24572_, _24568_);
  and (_24575_, _24574_, _08798_);
  nand (_24576_, _24575_, _24573_);
  nand (_24578_, _24576_, _24556_);
  or (_24579_, _24578_, _24552_);
  or (_24580_, _24556_, _23211_);
  and (_24581_, _24580_, _43000_);
  and (_24582_, _24581_, _24579_);
  or (_24583_, _24582_, _23144_);
  and (_43570_, _24583_, _41806_);
  or (_24584_, _05245_, \oc8051_golden_model_1.PSW [1]);
  and (_24585_, _12213_, _05245_);
  not (_24586_, _24585_);
  and (_24588_, _24586_, _24584_);
  or (_24589_, _24588_, _04081_);
  nand (_24590_, _05245_, _03274_);
  and (_24591_, _24590_, _24584_);
  and (_24592_, _24591_, _04409_);
  not (_24593_, \oc8051_golden_model_1.PSW [1]);
  nor (_24594_, _04409_, _24593_);
  or (_24595_, _24594_, _03610_);
  or (_24596_, _24595_, _24592_);
  and (_24597_, _24596_, _04055_);
  and (_24599_, _24597_, _24589_);
  and (_24600_, _12224_, _05901_);
  nor (_24601_, _05901_, _24593_);
  or (_24602_, _24601_, _03723_);
  or (_24603_, _24602_, _24600_);
  and (_24604_, _24603_, _14265_);
  or (_24605_, _24604_, _24599_);
  nor (_24606_, _05245_, _24593_);
  and (_24607_, _05245_, _06764_);
  or (_24608_, _24607_, _24606_);
  or (_24610_, _24608_, _03996_);
  and (_24611_, _24610_, _24605_);
  or (_24612_, _24611_, _03729_);
  or (_24613_, _24591_, _03737_);
  and (_24614_, _24613_, _03736_);
  and (_24615_, _24614_, _24612_);
  and (_24616_, _12211_, _05901_);
  or (_24617_, _24616_, _24601_);
  and (_24618_, _24617_, _03714_);
  or (_24619_, _24618_, _03719_);
  or (_24622_, _24619_, _24615_);
  and (_24623_, _24600_, _12239_);
  or (_24624_, _24601_, _06840_);
  or (_24625_, _24624_, _24623_);
  and (_24626_, _24625_, _24622_);
  and (_24627_, _24626_, _03710_);
  not (_24628_, _05901_);
  nor (_24629_, _12256_, _24628_);
  or (_24630_, _24601_, _24629_);
  and (_24631_, _24630_, _03505_);
  or (_24633_, _24631_, _07390_);
  or (_24634_, _24633_, _24627_);
  or (_24635_, _24608_, _06838_);
  and (_24636_, _24635_, _24634_);
  or (_24637_, _24636_, _04481_);
  and (_24638_, _06501_, _05245_);
  or (_24639_, _24606_, _07400_);
  or (_24640_, _24639_, _24638_);
  and (_24641_, _24640_, _03589_);
  and (_24642_, _24641_, _24637_);
  nor (_24644_, _12313_, _09661_);
  or (_24645_, _24644_, _24606_);
  and (_24646_, _24645_, _03222_);
  or (_24647_, _24646_, _24642_);
  and (_24648_, _24647_, _03602_);
  or (_24649_, _12327_, _09661_);
  and (_24650_, _24649_, _03600_);
  nand (_24651_, _05245_, _04303_);
  and (_24652_, _24651_, _03601_);
  or (_24653_, _24652_, _24650_);
  and (_24655_, _24653_, _24584_);
  or (_24656_, _24655_, _24648_);
  and (_24657_, _24656_, _07778_);
  or (_24658_, _12333_, _09661_);
  and (_24659_, _24584_, _03780_);
  and (_24660_, _24659_, _24658_);
  or (_24661_, _24660_, _24657_);
  and (_24662_, _24661_, _07777_);
  or (_24663_, _12207_, _09661_);
  and (_24664_, _24584_, _03622_);
  and (_24666_, _24664_, _24663_);
  or (_24667_, _24666_, _24662_);
  and (_24668_, _24667_, _06828_);
  or (_24669_, _24606_, _05618_);
  and (_24670_, _24591_, _03790_);
  and (_24671_, _24670_, _24669_);
  or (_24672_, _24671_, _24668_);
  and (_24673_, _24672_, _03786_);
  or (_24674_, _24651_, _05618_);
  and (_24675_, _24584_, _03624_);
  and (_24677_, _24675_, _24674_);
  or (_24678_, _24590_, _05618_);
  and (_24679_, _24584_, _03785_);
  and (_24680_, _24679_, _24678_);
  or (_24681_, _24680_, _03815_);
  or (_24682_, _24681_, _24677_);
  or (_24683_, _24682_, _24673_);
  or (_24684_, _24588_, _04246_);
  and (_24685_, _24684_, _03823_);
  and (_24686_, _24685_, _24683_);
  and (_24688_, _24617_, _03453_);
  or (_24689_, _24688_, _03447_);
  or (_24690_, _24689_, _24686_);
  or (_24691_, _24606_, _03514_);
  or (_24692_, _24691_, _24585_);
  and (_24693_, _24692_, _24690_);
  or (_24694_, _24693_, _43004_);
  or (_24695_, _43000_, \oc8051_golden_model_1.PSW [1]);
  and (_24696_, _24695_, _41806_);
  and (_43571_, _24696_, _24694_);
  and (_24698_, _07821_, \oc8051_golden_model_1.ACC [7]);
  nor (_24699_, _07821_, \oc8051_golden_model_1.ACC [7]);
  nor (_24700_, _24699_, _10295_);
  nor (_24701_, _24700_, _24698_);
  nand (_24702_, _24701_, _07890_);
  and (_24703_, _24698_, _07887_);
  nor (_24704_, _24703_, _07898_);
  and (_24705_, _24704_, _24702_);
  not (_24706_, \oc8051_golden_model_1.PSW [2]);
  nor (_24707_, _05245_, _24706_);
  not (_24709_, _24707_);
  or (_24710_, _12519_, _09661_);
  and (_24711_, _24710_, _24709_);
  or (_24712_, _24711_, _03589_);
  or (_24713_, _09661_, _04875_);
  and (_24714_, _24713_, _24709_);
  and (_24715_, _24714_, _07390_);
  not (_24716_, _08050_);
  nor (_24717_, _07987_, \oc8051_golden_model_1.ACC [7]);
  and (_24718_, _07987_, \oc8051_golden_model_1.ACC [7]);
  nor (_24720_, _24718_, _24717_);
  and (_24721_, _24720_, _10197_);
  nor (_24722_, _24720_, _10197_);
  or (_24723_, _24722_, _24721_);
  or (_24724_, _24723_, _24716_);
  nand (_24725_, _24723_, _24716_);
  and (_24726_, _24725_, _24724_);
  and (_24727_, _24726_, _08051_);
  not (_24728_, _07822_);
  and (_24729_, _10183_, _24728_);
  nor (_24731_, _10183_, _24728_);
  nor (_24732_, _24731_, _24729_);
  nor (_24733_, _24732_, _08177_);
  and (_24734_, _24732_, _08177_);
  or (_24735_, _24734_, _24733_);
  or (_24736_, _24735_, _08059_);
  nor (_24737_, _05901_, _24706_);
  and (_24738_, _12409_, _05901_);
  nor (_24739_, _24738_, _24737_);
  or (_24740_, _24739_, _03736_);
  and (_24742_, _24714_, _03723_);
  nor (_24743_, _12416_, _09661_);
  nor (_24744_, _24743_, _24707_);
  and (_24745_, _24744_, _03610_);
  and (_24746_, _05245_, \oc8051_golden_model_1.ACC [2]);
  nor (_24747_, _24746_, _24707_);
  or (_24748_, _24747_, _09029_);
  or (_24749_, _04409_, _24706_);
  and (_24750_, _24749_, _04081_);
  and (_24751_, _24750_, _24748_);
  or (_24753_, _24751_, _03715_);
  or (_24754_, _24753_, _24745_);
  not (_24755_, _24737_);
  nand (_24756_, _12411_, _05901_);
  and (_24757_, _24756_, _24755_);
  or (_24758_, _24757_, _04055_);
  and (_24759_, _24758_, _03996_);
  and (_24760_, _24759_, _24754_);
  or (_24761_, _24760_, _24742_);
  and (_24762_, _24761_, _03737_);
  and (_24764_, _24747_, _03729_);
  or (_24765_, _24764_, _03714_);
  or (_24766_, _24765_, _24762_);
  and (_24767_, _24766_, _24740_);
  or (_24768_, _24767_, _03719_);
  and (_24769_, _24755_, _10084_);
  or (_24770_, _24769_, _06840_);
  or (_24771_, _24770_, _24757_);
  and (_24772_, _24771_, _06875_);
  and (_24773_, _24772_, _24768_);
  or (_24775_, _14294_, _14181_);
  or (_24776_, _24775_, _14408_);
  or (_24777_, _24776_, _14527_);
  or (_24778_, _24777_, _14643_);
  or (_24779_, _24778_, _14758_);
  or (_24780_, _24779_, _07386_);
  nor (_24781_, _24780_, _14875_);
  or (_24782_, _24781_, _08060_);
  or (_24783_, _24782_, _24773_);
  and (_24784_, _24783_, _10201_);
  and (_24786_, _24784_, _24736_);
  or (_24787_, _24786_, _03761_);
  or (_24788_, _24787_, _24727_);
  nor (_24789_, _08520_, \oc8051_golden_model_1.ACC [7]);
  and (_24790_, _08520_, \oc8051_golden_model_1.ACC [7]);
  nor (_24791_, _24790_, _24789_);
  not (_24792_, _24791_);
  or (_24793_, _24792_, _10227_);
  nand (_24794_, _24792_, _10227_);
  and (_24795_, _24794_, _24793_);
  nand (_24797_, _24795_, _23615_);
  or (_24798_, _24795_, _23615_);
  and (_24799_, _24798_, _24797_);
  or (_24800_, _24799_, _03766_);
  and (_24801_, _24800_, _07914_);
  and (_24802_, _24801_, _24788_);
  nor (_24803_, _07919_, \oc8051_golden_model_1.ACC [7]);
  and (_24804_, _07919_, \oc8051_golden_model_1.ACC [7]);
  nor (_24805_, _24804_, _24803_);
  nor (_24806_, _24805_, _10239_);
  and (_24808_, _24805_, _10239_);
  or (_24809_, _24808_, _24806_);
  or (_24810_, _24809_, _07984_);
  nand (_24811_, _24809_, _07984_);
  and (_24812_, _24811_, _24810_);
  and (_24813_, _24812_, _07913_);
  or (_24814_, _24813_, _03505_);
  or (_24815_, _24814_, _24802_);
  or (_24816_, _12461_, _24628_);
  and (_24817_, _24816_, _24755_);
  or (_24819_, _24817_, _03710_);
  and (_24820_, _24819_, _06838_);
  and (_24821_, _24820_, _24815_);
  or (_24822_, _24821_, _24715_);
  and (_24823_, _24822_, _07400_);
  nand (_24824_, _06637_, _05245_);
  nor (_24825_, _24707_, _07400_);
  and (_24826_, _24825_, _24824_);
  or (_24827_, _24826_, _03222_);
  or (_24828_, _24827_, _24823_);
  and (_24830_, _24828_, _24712_);
  or (_24831_, _24830_, _07405_);
  nor (_24832_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and (_24833_, _24832_, _07431_);
  nand (_24834_, _24833_, _07405_);
  and (_24835_, _24834_, _03602_);
  and (_24836_, _24835_, _24831_);
  nand (_24837_, _12533_, _05245_);
  nor (_24838_, _24707_, _07766_);
  and (_24839_, _24838_, _24837_);
  and (_24841_, _05245_, _06332_);
  nor (_24842_, _24841_, _24707_);
  and (_24843_, _24842_, _03601_);
  or (_24844_, _24843_, _03780_);
  or (_24845_, _24844_, _24839_);
  or (_24846_, _24845_, _24836_);
  nand (_24847_, _12539_, _05245_);
  and (_24848_, _24847_, _24709_);
  or (_24849_, _24848_, _07778_);
  and (_24850_, _24849_, _24846_);
  or (_24852_, _24850_, _03622_);
  and (_24853_, _24709_, _05717_);
  or (_24854_, _24842_, _07777_);
  or (_24855_, _24854_, _24853_);
  and (_24856_, _24855_, _24852_);
  or (_24857_, _24856_, _03790_);
  or (_24858_, _24747_, _06828_);
  or (_24859_, _24858_, _24853_);
  and (_24860_, _24859_, _07795_);
  and (_24861_, _24860_, _24857_);
  or (_24863_, _12532_, _09661_);
  nor (_24864_, _24707_, _07795_);
  and (_24865_, _24864_, _24863_);
  or (_24866_, _24865_, _03785_);
  or (_24867_, _24866_, _24861_);
  or (_24868_, _12538_, _09661_);
  and (_24869_, _24868_, _24709_);
  or (_24870_, _24869_, _07793_);
  and (_24871_, _24870_, _07898_);
  and (_24872_, _24871_, _24867_);
  or (_24874_, _24872_, _24705_);
  and (_24875_, _24874_, _08477_);
  nand (_24876_, _24718_, _08499_);
  nor (_24877_, _24717_, _10301_);
  nor (_24878_, _24877_, _24718_);
  nand (_24879_, _24878_, _08502_);
  and (_24880_, _24879_, _24876_);
  and (_24881_, _24880_, _08475_);
  or (_24882_, _24881_, _03776_);
  or (_24883_, _24882_, _24875_);
  nand (_24885_, _24790_, _08580_);
  nor (_24886_, _24792_, _10307_);
  nor (_24887_, _24886_, _24790_);
  nand (_24888_, _24887_, _08583_);
  and (_24889_, _24888_, _24885_);
  or (_24890_, _24889_, _03777_);
  and (_24891_, _24890_, _08589_);
  and (_24892_, _24891_, _24883_);
  nand (_24893_, _24804_, _08610_);
  nor (_24894_, _24803_, _10313_);
  or (_24896_, _24804_, _24358_);
  or (_24897_, _24896_, _24894_);
  and (_24898_, _24897_, _24893_);
  and (_24899_, _24898_, _08506_);
  or (_24900_, _24899_, _08618_);
  or (_24901_, _24900_, _24892_);
  nor (_24902_, _08693_, _08374_);
  nand (_24903_, _10331_, _08618_);
  or (_24904_, _24903_, _24902_);
  and (_24905_, _24904_, _08624_);
  nand (_24907_, _24905_, _24901_);
  nor (_24908_, _08657_, _24176_);
  and (_24909_, _08657_, _08399_);
  or (_24910_, _24909_, _08624_);
  or (_24911_, _24910_, _24908_);
  and (_24912_, _24911_, _08702_);
  and (_24913_, _24912_, _24907_);
  or (_24914_, _08725_, _08188_);
  and (_24915_, _24914_, _10354_);
  or (_24916_, _08765_, _08406_);
  and (_24918_, _10349_, _24916_);
  or (_24919_, _24918_, _03815_);
  or (_24920_, _24919_, _24915_);
  or (_24921_, _24920_, _24913_);
  nand (_24922_, _24744_, _03815_);
  and (_24923_, _24922_, _03823_);
  and (_24924_, _24923_, _24921_);
  nor (_24925_, _24739_, _03823_);
  or (_24926_, _24925_, _03447_);
  or (_24927_, _24926_, _24924_);
  and (_24929_, _12592_, _05245_);
  or (_24930_, _24707_, _03514_);
  or (_24931_, _24930_, _24929_);
  and (_24932_, _24931_, _24927_);
  or (_24933_, _24932_, _43004_);
  or (_24934_, _43000_, \oc8051_golden_model_1.PSW [2]);
  and (_24935_, _24934_, _41806_);
  and (_43572_, _24935_, _24933_);
  nor (_24936_, _05245_, _05018_);
  and (_24937_, _05245_, _06276_);
  nor (_24939_, _24937_, _24936_);
  and (_24940_, _24939_, _03601_);
  nor (_24941_, _09661_, _05005_);
  nor (_24942_, _24941_, _24936_);
  and (_24943_, _24942_, _07390_);
  and (_24944_, _05245_, \oc8051_golden_model_1.ACC [3]);
  nor (_24945_, _24944_, _24936_);
  nor (_24946_, _24945_, _09029_);
  nor (_24947_, _04409_, _05018_);
  or (_24948_, _24947_, _24946_);
  and (_24950_, _24948_, _04081_);
  nor (_24951_, _12627_, _09661_);
  nor (_24952_, _24951_, _24936_);
  nor (_24953_, _24952_, _04081_);
  or (_24954_, _24953_, _24950_);
  and (_24955_, _24954_, _04055_);
  nor (_24956_, _05901_, _05018_);
  and (_24957_, _12631_, _05901_);
  nor (_24958_, _24957_, _24956_);
  nor (_24959_, _24958_, _04055_);
  or (_24961_, _24959_, _03723_);
  or (_24962_, _24961_, _24955_);
  nand (_24963_, _24942_, _03723_);
  and (_24964_, _24963_, _24962_);
  and (_24965_, _24964_, _03737_);
  nor (_24966_, _24945_, _03737_);
  or (_24967_, _24966_, _24965_);
  and (_24968_, _24967_, _03736_);
  and (_24969_, _12641_, _05901_);
  nor (_24970_, _24969_, _24956_);
  nor (_24972_, _24970_, _03736_);
  or (_24973_, _24972_, _03719_);
  or (_24974_, _24973_, _24968_);
  nor (_24975_, _24956_, _12648_);
  nor (_24976_, _24975_, _24958_);
  or (_24977_, _24976_, _06840_);
  and (_24978_, _24977_, _03710_);
  and (_24979_, _24978_, _24974_);
  nor (_24980_, _12612_, _24628_);
  nor (_24981_, _24980_, _24956_);
  nor (_24983_, _24981_, _03710_);
  nor (_24984_, _24983_, _07390_);
  not (_24985_, _24984_);
  nor (_24986_, _24985_, _24979_);
  nor (_24987_, _24986_, _24943_);
  nor (_24988_, _24987_, _04481_);
  and (_24989_, _06592_, _05245_);
  nor (_24990_, _24936_, _07400_);
  not (_24991_, _24990_);
  nor (_24992_, _24991_, _24989_);
  or (_24994_, _24992_, _03222_);
  nor (_24995_, _24994_, _24988_);
  nor (_24996_, _12718_, _09661_);
  nor (_24997_, _24936_, _24996_);
  nor (_24998_, _24997_, _03589_);
  or (_24999_, _24998_, _03601_);
  nor (_25000_, _24999_, _24995_);
  nor (_25001_, _25000_, _24940_);
  or (_25002_, _25001_, _03600_);
  and (_25003_, _12733_, _05245_);
  or (_25005_, _25003_, _24936_);
  or (_25006_, _25005_, _07766_);
  and (_25007_, _25006_, _07778_);
  and (_25008_, _25007_, _25002_);
  and (_25009_, _12739_, _05245_);
  nor (_25010_, _25009_, _24936_);
  nor (_25011_, _25010_, _07778_);
  nor (_25012_, _25011_, _25008_);
  nor (_25013_, _25012_, _03622_);
  nor (_25014_, _24936_, _05567_);
  not (_25016_, _25014_);
  nor (_25017_, _24939_, _07777_);
  and (_25018_, _25017_, _25016_);
  nor (_25019_, _25018_, _25013_);
  nor (_25020_, _25019_, _03790_);
  nor (_25021_, _24945_, _06828_);
  and (_25022_, _25021_, _25016_);
  nor (_25023_, _25022_, _03624_);
  not (_25024_, _25023_);
  nor (_25025_, _25024_, _25020_);
  nor (_25027_, _12732_, _09661_);
  or (_25028_, _24936_, _07795_);
  nor (_25029_, _25028_, _25027_);
  or (_25030_, _25029_, _03785_);
  nor (_25031_, _25030_, _25025_);
  nor (_25032_, _12738_, _09661_);
  nor (_25033_, _25032_, _24936_);
  nor (_25034_, _25033_, _07793_);
  or (_25035_, _25034_, _25031_);
  and (_25036_, _25035_, _04246_);
  nor (_25038_, _24952_, _04246_);
  or (_25039_, _25038_, _25036_);
  and (_25040_, _25039_, _03823_);
  nor (_25041_, _24970_, _03823_);
  or (_25042_, _25041_, _25040_);
  and (_25043_, _25042_, _03514_);
  and (_25044_, _12794_, _05245_);
  nor (_25045_, _25044_, _24936_);
  nor (_25046_, _25045_, _03514_);
  or (_25047_, _25046_, _25043_);
  or (_25049_, _25047_, _43004_);
  or (_25050_, _43000_, \oc8051_golden_model_1.PSW [3]);
  and (_25051_, _25050_, _41806_);
  and (_43573_, _25051_, _25049_);
  not (_25052_, \oc8051_golden_model_1.PSW [4]);
  nor (_25053_, _05245_, _25052_);
  nor (_25054_, _05777_, _09661_);
  nor (_25055_, _25054_, _25053_);
  and (_25056_, _25055_, _07390_);
  nor (_25057_, _05901_, _25052_);
  and (_25059_, _12827_, _05901_);
  nor (_25060_, _25059_, _25057_);
  nor (_25061_, _25060_, _03736_);
  and (_25062_, _05245_, \oc8051_golden_model_1.ACC [4]);
  nor (_25063_, _25062_, _25053_);
  nor (_25064_, _25063_, _09029_);
  nor (_25065_, _04409_, _25052_);
  or (_25066_, _25065_, _25064_);
  and (_25067_, _25066_, _04081_);
  nor (_25068_, _12841_, _09661_);
  nor (_25070_, _25068_, _25053_);
  nor (_25071_, _25070_, _04081_);
  or (_25072_, _25071_, _25067_);
  and (_25073_, _25072_, _04055_);
  and (_25074_, _12845_, _05901_);
  nor (_25075_, _25074_, _25057_);
  nor (_25076_, _25075_, _04055_);
  or (_25077_, _25076_, _03723_);
  or (_25078_, _25077_, _25073_);
  nand (_25079_, _25055_, _03723_);
  and (_25081_, _25079_, _25078_);
  and (_25082_, _25081_, _03737_);
  nor (_25083_, _25063_, _03737_);
  or (_25084_, _25083_, _25082_);
  and (_25085_, _25084_, _03736_);
  nor (_25086_, _25085_, _25061_);
  nor (_25087_, _25086_, _03719_);
  nor (_25088_, _25057_, _12860_);
  or (_25089_, _25075_, _06840_);
  nor (_25090_, _25089_, _25088_);
  nor (_25092_, _25090_, _25087_);
  nor (_25093_, _25092_, _03505_);
  nor (_25094_, _12825_, _24628_);
  nor (_25095_, _25094_, _25057_);
  nor (_25096_, _25095_, _03710_);
  nor (_25097_, _25096_, _07390_);
  not (_25098_, _25097_);
  nor (_25099_, _25098_, _25093_);
  nor (_25100_, _25099_, _25056_);
  nor (_25101_, _25100_, _04481_);
  and (_25102_, _06730_, _05245_);
  nor (_25103_, _25053_, _07400_);
  not (_25104_, _25103_);
  nor (_25105_, _25104_, _25102_);
  nor (_25106_, _25105_, _03222_);
  not (_25107_, _25106_);
  nor (_25108_, _25107_, _25101_);
  nor (_25109_, _12933_, _09661_);
  nor (_25110_, _25109_, _25053_);
  nor (_25111_, _25110_, _03589_);
  or (_25114_, _25111_, _08828_);
  or (_25115_, _25114_, _25108_);
  and (_25116_, _12821_, _05245_);
  or (_25117_, _25053_, _07766_);
  or (_25118_, _25117_, _25116_);
  and (_25119_, _06298_, _05245_);
  nor (_25120_, _25119_, _25053_);
  and (_25121_, _25120_, _03601_);
  nor (_25122_, _25121_, _03780_);
  and (_25123_, _25122_, _25118_);
  and (_25125_, _25123_, _25115_);
  and (_25126_, _12817_, _05245_);
  nor (_25127_, _25126_, _25053_);
  nor (_25128_, _25127_, _07778_);
  nor (_25129_, _25128_, _25125_);
  nor (_25130_, _25129_, _03622_);
  nor (_25131_, _25053_, _05825_);
  not (_25132_, _25131_);
  nor (_25133_, _25120_, _07777_);
  and (_25134_, _25133_, _25132_);
  nor (_25136_, _25134_, _25130_);
  nor (_25137_, _25136_, _03790_);
  nor (_25138_, _25063_, _06828_);
  and (_25139_, _25138_, _25132_);
  nor (_25140_, _25139_, _03624_);
  not (_25141_, _25140_);
  nor (_25142_, _25141_, _25137_);
  nor (_25143_, _12819_, _09661_);
  or (_25144_, _25053_, _07795_);
  nor (_25145_, _25144_, _25143_);
  or (_25146_, _25145_, _03785_);
  nor (_25147_, _25146_, _25142_);
  nor (_25148_, _12816_, _09661_);
  nor (_25149_, _25148_, _25053_);
  nor (_25150_, _25149_, _07793_);
  or (_25151_, _25150_, _25147_);
  and (_25152_, _25151_, _04246_);
  nor (_25153_, _25070_, _04246_);
  or (_25154_, _25153_, _25152_);
  and (_25155_, _25154_, _03823_);
  nor (_25158_, _25060_, _03823_);
  or (_25159_, _25158_, _25155_);
  and (_25160_, _25159_, _03514_);
  and (_25161_, _13003_, _05245_);
  nor (_25162_, _25161_, _25053_);
  nor (_25163_, _25162_, _03514_);
  or (_25164_, _25163_, _25160_);
  or (_25165_, _25164_, _43004_);
  or (_25166_, _43000_, \oc8051_golden_model_1.PSW [4]);
  and (_25167_, _25166_, _41806_);
  and (_43574_, _25167_, _25165_);
  not (_25169_, \oc8051_golden_model_1.PSW [5]);
  nor (_25170_, _05245_, _25169_);
  and (_25171_, _06684_, _05245_);
  or (_25172_, _25171_, _25170_);
  and (_25173_, _25172_, _04481_);
  and (_25174_, _05245_, \oc8051_golden_model_1.ACC [5]);
  nor (_25175_, _25174_, _25170_);
  nor (_25176_, _25175_, _09029_);
  nor (_25177_, _04409_, _25169_);
  or (_25178_, _25177_, _25176_);
  and (_25179_, _25178_, _04081_);
  nor (_25180_, _13014_, _09661_);
  nor (_25181_, _25180_, _25170_);
  nor (_25182_, _25181_, _04081_);
  or (_25183_, _25182_, _25179_);
  and (_25184_, _25183_, _04055_);
  nor (_25185_, _05901_, _25169_);
  and (_25186_, _13037_, _05901_);
  nor (_25187_, _25186_, _25185_);
  nor (_25190_, _25187_, _04055_);
  or (_25191_, _25190_, _03723_);
  or (_25192_, _25191_, _25184_);
  nor (_25193_, _05469_, _09661_);
  nor (_25194_, _25193_, _25170_);
  nand (_25195_, _25194_, _03723_);
  and (_25196_, _25195_, _25192_);
  and (_25197_, _25196_, _03737_);
  nor (_25198_, _25175_, _03737_);
  or (_25199_, _25198_, _25197_);
  and (_25201_, _25199_, _03736_);
  and (_25202_, _13047_, _05901_);
  nor (_25203_, _25202_, _25185_);
  nor (_25204_, _25203_, _03736_);
  or (_25205_, _25204_, _25201_);
  and (_25206_, _25205_, _06840_);
  nor (_25207_, _25185_, _13054_);
  nor (_25208_, _25207_, _25187_);
  and (_25209_, _25208_, _03719_);
  or (_25210_, _25209_, _25206_);
  and (_25212_, _25210_, _03710_);
  nor (_25213_, _13020_, _24628_);
  nor (_25214_, _25213_, _25185_);
  nor (_25215_, _25214_, _03710_);
  nor (_25216_, _25215_, _07390_);
  not (_25217_, _25216_);
  nor (_25218_, _25217_, _25212_);
  and (_25219_, _25194_, _07390_);
  or (_25220_, _25219_, _04481_);
  nor (_25221_, _25220_, _25218_);
  or (_25223_, _25221_, _25173_);
  and (_25224_, _25223_, _03589_);
  nor (_25225_, _13127_, _09661_);
  nor (_25226_, _25225_, _25170_);
  nor (_25227_, _25226_, _03589_);
  or (_25228_, _25227_, _08828_);
  or (_25229_, _25228_, _25224_);
  and (_25230_, _13141_, _05245_);
  or (_25231_, _25170_, _07766_);
  or (_25232_, _25231_, _25230_);
  and (_25233_, _06306_, _05245_);
  nor (_25234_, _25233_, _25170_);
  and (_25235_, _25234_, _03601_);
  nor (_25236_, _25235_, _03780_);
  and (_25237_, _25236_, _25232_);
  and (_25238_, _25237_, _25229_);
  and (_25239_, _13147_, _05245_);
  nor (_25240_, _25239_, _25170_);
  nor (_25241_, _25240_, _07778_);
  nor (_25242_, _25241_, _25238_);
  nor (_25245_, _25242_, _03622_);
  nor (_25246_, _25170_, _05518_);
  not (_25247_, _25246_);
  nor (_25248_, _25234_, _07777_);
  and (_25249_, _25248_, _25247_);
  nor (_25250_, _25249_, _25245_);
  nor (_25251_, _25250_, _03790_);
  nor (_25252_, _25175_, _06828_);
  and (_25253_, _25252_, _25247_);
  nor (_25254_, _25253_, _03624_);
  not (_25256_, _25254_);
  nor (_25257_, _25256_, _25251_);
  nor (_25258_, _13140_, _09661_);
  or (_25259_, _25170_, _07795_);
  nor (_25260_, _25259_, _25258_);
  or (_25261_, _25260_, _03785_);
  nor (_25262_, _25261_, _25257_);
  nor (_25263_, _13146_, _09661_);
  nor (_25264_, _25263_, _25170_);
  nor (_25265_, _25264_, _07793_);
  or (_25267_, _25265_, _25262_);
  and (_25268_, _25267_, _04246_);
  nor (_25269_, _25181_, _04246_);
  or (_25270_, _25269_, _25268_);
  and (_25271_, _25270_, _03823_);
  nor (_25272_, _25203_, _03823_);
  or (_25273_, _25272_, _25271_);
  and (_25274_, _25273_, _03514_);
  and (_25275_, _13199_, _05245_);
  nor (_25276_, _25275_, _25170_);
  nor (_25278_, _25276_, _03514_);
  or (_25279_, _25278_, _25274_);
  or (_25280_, _25279_, _43004_);
  or (_25281_, _43000_, \oc8051_golden_model_1.PSW [5]);
  and (_25282_, _25281_, _41806_);
  and (_43575_, _25282_, _25280_);
  not (_25283_, _08574_);
  nor (_25284_, _25283_, _08516_);
  nor (_25285_, _25284_, _03777_);
  nor (_25286_, _05245_, _15859_);
  nor (_25288_, _05363_, _09661_);
  nor (_25289_, _25288_, _25286_);
  and (_25290_, _25289_, _07390_);
  nor (_25291_, _08516_, _03766_);
  not (_25292_, _25291_);
  nor (_25293_, _25292_, _10223_);
  nor (_25294_, _08042_, _08006_);
  or (_25295_, _25294_, _10201_);
  or (_25296_, _08059_, _07834_);
  nor (_25297_, _25296_, _08173_);
  nor (_25299_, _05901_, _15859_);
  and (_25300_, _13253_, _05901_);
  nor (_25301_, _25300_, _25299_);
  nor (_25302_, _25301_, _03736_);
  and (_25303_, _05245_, \oc8051_golden_model_1.ACC [6]);
  nor (_25304_, _25303_, _25286_);
  nor (_25305_, _25304_, _09029_);
  nor (_25306_, _04409_, _15859_);
  or (_25307_, _25306_, _25305_);
  and (_25308_, _25307_, _04081_);
  nor (_25310_, _13242_, _09661_);
  nor (_25311_, _25310_, _25286_);
  nor (_25312_, _25311_, _04081_);
  or (_25313_, _25312_, _25308_);
  and (_25314_, _25313_, _04055_);
  and (_25315_, _13229_, _05901_);
  nor (_25316_, _25315_, _25299_);
  nor (_25317_, _25316_, _04055_);
  or (_25318_, _25317_, _03723_);
  or (_25319_, _25318_, _25314_);
  nand (_25321_, _25289_, _03723_);
  and (_25322_, _25321_, _25319_);
  and (_25323_, _25322_, _03737_);
  nor (_25324_, _25304_, _03737_);
  or (_25325_, _25324_, _25323_);
  and (_25326_, _25325_, _03736_);
  nor (_25327_, _25326_, _25302_);
  nor (_25328_, _25327_, _03719_);
  nor (_25329_, _25299_, _13260_);
  or (_25330_, _25329_, _06840_);
  nor (_25332_, _25330_, _25316_);
  or (_25333_, _25332_, _08060_);
  nor (_25334_, _25333_, _25328_);
  or (_25335_, _25334_, _25297_);
  or (_25336_, _25335_, _08051_);
  and (_25337_, _25336_, _03766_);
  and (_25338_, _25337_, _25295_);
  nor (_25339_, _25338_, _25293_);
  nor (_25340_, _25339_, _07913_);
  or (_25341_, _07916_, _07914_);
  nor (_25343_, _25341_, _07977_);
  or (_25344_, _25343_, _03505_);
  nor (_25345_, _25344_, _25340_);
  nor (_25346_, _13226_, _24628_);
  nor (_25347_, _25346_, _25299_);
  nor (_25348_, _25347_, _03710_);
  nor (_25349_, _25348_, _07390_);
  not (_25350_, _25349_);
  nor (_25351_, _25350_, _25345_);
  nor (_25352_, _25351_, _25290_);
  nor (_25354_, _25352_, _04481_);
  and (_25355_, _06455_, _05245_);
  nor (_25356_, _25286_, _07400_);
  not (_25357_, _25356_);
  nor (_25358_, _25357_, _25355_);
  nor (_25359_, _25358_, _03222_);
  not (_25360_, _25359_);
  nor (_25361_, _25360_, _25354_);
  nor (_25362_, _13332_, _09661_);
  nor (_25363_, _25362_, _25286_);
  nor (_25364_, _25363_, _03589_);
  or (_25365_, _25364_, _08828_);
  or (_25366_, _25365_, _25361_);
  and (_25367_, _13347_, _05245_);
  or (_25368_, _25286_, _07766_);
  or (_25369_, _25368_, _25367_);
  and (_25370_, _13339_, _05245_);
  nor (_25371_, _25370_, _25286_);
  and (_25372_, _25371_, _03601_);
  nor (_25373_, _25372_, _03780_);
  and (_25376_, _25373_, _25369_);
  and (_25377_, _25376_, _25366_);
  and (_25378_, _13353_, _05245_);
  nor (_25379_, _25378_, _25286_);
  nor (_25380_, _25379_, _07778_);
  nor (_25381_, _25380_, _25377_);
  nor (_25382_, _25381_, _03622_);
  nor (_25383_, _25286_, _05412_);
  not (_25384_, _25383_);
  nor (_25385_, _25371_, _07777_);
  and (_25387_, _25385_, _25384_);
  nor (_25388_, _25387_, _25382_);
  nor (_25389_, _25388_, _03790_);
  nor (_25390_, _25304_, _06828_);
  and (_25391_, _25390_, _25384_);
  or (_25392_, _25391_, _25389_);
  and (_25393_, _25392_, _07795_);
  nor (_25394_, _13346_, _09661_);
  nor (_25395_, _25394_, _25286_);
  nor (_25396_, _25395_, _07795_);
  or (_25398_, _25396_, _25393_);
  and (_25399_, _25398_, _07793_);
  not (_25400_, _07897_);
  nor (_25401_, _13352_, _09661_);
  nor (_25402_, _25401_, _25286_);
  nor (_25403_, _25402_, _07793_);
  nor (_25404_, _25403_, _25400_);
  not (_25405_, _25404_);
  nor (_25406_, _25405_, _25399_);
  not (_25407_, _07834_);
  and (_25409_, _07881_, _25407_);
  nor (_25410_, _25409_, _07891_);
  nor (_25411_, _25410_, _07898_);
  nor (_25412_, _25411_, _25406_);
  nor (_25413_, _25409_, _07892_);
  nor (_25414_, _25413_, _08475_);
  not (_25415_, _25414_);
  nor (_25416_, _25415_, _25412_);
  nor (_25417_, _08477_, _08006_);
  and (_25418_, _25417_, _08493_);
  nor (_25420_, _25418_, _03776_);
  not (_25421_, _25420_);
  nor (_25422_, _25421_, _25416_);
  nor (_25423_, _25422_, _25285_);
  nor (_25424_, _25423_, _08506_);
  not (_25425_, _07916_);
  and (_25426_, _08604_, _25425_);
  nor (_25427_, _25426_, _08589_);
  nor (_25428_, _25427_, _11907_);
  not (_25429_, _25428_);
  nor (_25431_, _25429_, _25424_);
  and (_25432_, _08687_, _08618_);
  nor (_25433_, _08651_, _08624_);
  or (_25434_, _25433_, _03517_);
  nor (_25435_, _25434_, _25432_);
  not (_25436_, _25435_);
  nor (_25437_, _25436_, _25431_);
  and (_25438_, _08719_, _03517_);
  or (_25439_, _25438_, _08701_);
  nor (_25440_, _25439_, _25437_);
  nor (_25442_, _08759_, _08734_);
  nor (_25443_, _25442_, _25440_);
  and (_25444_, _25443_, _04246_);
  nor (_25445_, _25311_, _04246_);
  or (_25446_, _25445_, _25444_);
  and (_25447_, _25446_, _03823_);
  nor (_25448_, _25301_, _03823_);
  or (_25449_, _25448_, _25447_);
  and (_25450_, _25449_, _03514_);
  and (_25451_, _13402_, _05245_);
  nor (_25453_, _25286_, _25451_);
  nor (_25454_, _25453_, _03514_);
  or (_25455_, _25454_, _25450_);
  or (_25456_, _25455_, _43004_);
  or (_25457_, _43000_, \oc8051_golden_model_1.PSW [6]);
  and (_25458_, _25457_, _41806_);
  and (_43576_, _25458_, _25456_);
  not (_25459_, \oc8051_golden_model_1.PCON [0]);
  nor (_25460_, _05212_, _25459_);
  nor (_25461_, _05666_, _10377_);
  nor (_25463_, _25461_, _25460_);
  and (_25464_, _25463_, _17166_);
  and (_25465_, _05212_, \oc8051_golden_model_1.ACC [0]);
  nor (_25466_, _25465_, _25460_);
  nor (_25467_, _25466_, _03737_);
  nor (_25468_, _25467_, _07390_);
  nor (_25469_, _25463_, _04081_);
  nor (_25470_, _04409_, _25459_);
  nor (_25471_, _25466_, _09029_);
  nor (_25472_, _25471_, _25470_);
  nor (_25474_, _25472_, _03610_);
  or (_25475_, _25474_, _03723_);
  nor (_25476_, _25475_, _25469_);
  or (_25477_, _25476_, _03729_);
  and (_25478_, _25477_, _25468_);
  and (_25479_, _05212_, _04620_);
  and (_25480_, _06838_, _03996_);
  or (_25481_, _25480_, _25460_);
  nor (_25482_, _25481_, _25479_);
  nor (_25483_, _25482_, _25478_);
  nor (_25485_, _25483_, _04481_);
  and (_25486_, _06546_, _05212_);
  nor (_25487_, _25460_, _07400_);
  not (_25488_, _25487_);
  nor (_25489_, _25488_, _25486_);
  nor (_25490_, _25489_, _25485_);
  nor (_25491_, _25490_, _03222_);
  nor (_25492_, _12109_, _10377_);
  or (_25493_, _25460_, _03589_);
  nor (_25494_, _25493_, _25492_);
  or (_25496_, _25494_, _03601_);
  nor (_25497_, _25496_, _25491_);
  and (_25498_, _05212_, _06274_);
  nor (_25499_, _25498_, _25460_);
  nand (_25500_, _25499_, _07766_);
  and (_25501_, _25500_, _08828_);
  nor (_25502_, _25501_, _25497_);
  and (_25503_, _12124_, _05212_);
  nor (_25504_, _25503_, _25460_);
  and (_25505_, _25504_, _03600_);
  nor (_25507_, _25505_, _25502_);
  nor (_25508_, _25507_, _03780_);
  and (_25509_, _12128_, _05212_);
  or (_25510_, _25460_, _07778_);
  nor (_25511_, _25510_, _25509_);
  or (_25512_, _25511_, _03622_);
  nor (_25513_, _25512_, _25508_);
  or (_25514_, _25499_, _07777_);
  nor (_25515_, _25514_, _25461_);
  nor (_25516_, _25515_, _25513_);
  nor (_25518_, _25516_, _03790_);
  and (_25519_, _12005_, _05212_);
  or (_25520_, _25519_, _25460_);
  and (_25521_, _25520_, _03790_);
  or (_25522_, _25521_, _25518_);
  and (_25523_, _25522_, _07795_);
  nor (_25524_, _12122_, _10377_);
  nor (_25525_, _25524_, _25460_);
  nor (_25526_, _25525_, _07795_);
  or (_25527_, _25526_, _25523_);
  and (_25529_, _25527_, _07793_);
  nor (_25530_, _12003_, _10377_);
  nor (_25531_, _25530_, _25460_);
  nor (_25532_, _25531_, _07793_);
  nor (_25533_, _25532_, _17166_);
  not (_25534_, _25533_);
  nor (_25535_, _25534_, _25529_);
  nor (_25536_, _25535_, _25464_);
  or (_25537_, _25536_, _43004_);
  or (_25538_, _43000_, \oc8051_golden_model_1.PCON [0]);
  and (_25539_, _25538_, _41806_);
  and (_43579_, _25539_, _25537_);
  and (_25540_, _06501_, _05212_);
  not (_25541_, \oc8051_golden_model_1.PCON [1]);
  nor (_25542_, _05212_, _25541_);
  nor (_25543_, _25542_, _07400_);
  not (_25544_, _25543_);
  nor (_25545_, _25544_, _25540_);
  not (_25546_, _25545_);
  nor (_25547_, _05212_, \oc8051_golden_model_1.PCON [1]);
  and (_25550_, _05212_, _03274_);
  nor (_25551_, _25550_, _25547_);
  and (_25552_, _25551_, _03729_);
  and (_25553_, _25551_, _04409_);
  nor (_25554_, _04409_, _25541_);
  or (_25555_, _25554_, _25553_);
  and (_25556_, _25555_, _04081_);
  and (_25557_, _12213_, _05212_);
  nor (_25558_, _25557_, _25547_);
  and (_25559_, _25558_, _03610_);
  or (_25561_, _25559_, _25556_);
  and (_25562_, _25561_, _03996_);
  and (_25563_, _05212_, _06764_);
  nor (_25564_, _25563_, _25542_);
  nor (_25565_, _25564_, _03996_);
  nor (_25566_, _25565_, _25562_);
  nor (_25567_, _25566_, _03729_);
  or (_25568_, _25567_, _07390_);
  nor (_25569_, _25568_, _25552_);
  and (_25570_, _25564_, _07390_);
  nor (_25572_, _25570_, _25569_);
  nor (_25573_, _25572_, _04481_);
  nor (_25574_, _25573_, _03222_);
  and (_25575_, _25574_, _25546_);
  not (_25576_, _25547_);
  and (_25577_, _12313_, _05212_);
  nor (_25578_, _25577_, _03589_);
  and (_25579_, _25578_, _25576_);
  nor (_25580_, _25579_, _25575_);
  nor (_25581_, _25580_, _08828_);
  nor (_25583_, _12327_, _10377_);
  nor (_25584_, _25583_, _07766_);
  and (_25585_, _05212_, _04303_);
  nor (_25586_, _25585_, _05886_);
  nor (_25587_, _25586_, _25584_);
  nor (_25588_, _25587_, _25547_);
  nor (_25589_, _25588_, _25581_);
  nor (_25590_, _25589_, _03780_);
  nor (_25591_, _12333_, _10377_);
  nor (_25592_, _25591_, _07778_);
  and (_25594_, _25592_, _25576_);
  nor (_25595_, _25594_, _25590_);
  nor (_25596_, _25595_, _03622_);
  nor (_25597_, _12207_, _10377_);
  nor (_25598_, _25597_, _07777_);
  and (_25599_, _25598_, _25576_);
  nor (_25600_, _25599_, _25596_);
  nor (_25601_, _25600_, _03790_);
  nor (_25602_, _25542_, _05618_);
  nor (_25603_, _25602_, _06828_);
  and (_25605_, _25603_, _25551_);
  nor (_25606_, _25605_, _25601_);
  or (_25607_, _25606_, _18499_);
  and (_25608_, _25585_, _05617_);
  or (_25609_, _25547_, _07795_);
  or (_25610_, _25609_, _25608_);
  and (_25611_, _25550_, _05617_);
  or (_25612_, _25547_, _07793_);
  or (_25613_, _25612_, _25611_);
  and (_25614_, _25613_, _04246_);
  and (_25616_, _25614_, _25610_);
  and (_25617_, _25616_, _25607_);
  nor (_25618_, _25558_, _04246_);
  nor (_25619_, _25618_, _25617_);
  and (_25620_, _25619_, _03514_);
  nor (_25621_, _25557_, _25542_);
  nor (_25622_, _25621_, _03514_);
  or (_25623_, _25622_, _25620_);
  or (_25624_, _25623_, _43004_);
  or (_25625_, _43000_, \oc8051_golden_model_1.PCON [1]);
  and (_25627_, _25625_, _41806_);
  and (_43580_, _25627_, _25624_);
  not (_25628_, \oc8051_golden_model_1.PCON [2]);
  nor (_25629_, _05212_, _25628_);
  nor (_25630_, _12538_, _10377_);
  nor (_25631_, _25630_, _25629_);
  nor (_25632_, _25631_, _07793_);
  and (_25633_, _12539_, _05212_);
  nor (_25634_, _25633_, _25629_);
  nor (_25635_, _25634_, _07778_);
  nor (_25637_, _10377_, _04875_);
  nor (_25638_, _25637_, _25629_);
  and (_25639_, _25638_, _07390_);
  and (_25640_, _05212_, \oc8051_golden_model_1.ACC [2]);
  nor (_25641_, _25640_, _25629_);
  nor (_25642_, _25641_, _03737_);
  nor (_25643_, _25641_, _09029_);
  nor (_25644_, _04409_, _25628_);
  or (_25645_, _25644_, _25643_);
  and (_25646_, _25645_, _04081_);
  nor (_25648_, _12416_, _10377_);
  nor (_25649_, _25648_, _25629_);
  nor (_25650_, _25649_, _04081_);
  or (_25651_, _25650_, _25646_);
  and (_25652_, _25651_, _03996_);
  nor (_25653_, _25638_, _03996_);
  nor (_25654_, _25653_, _25652_);
  nor (_25655_, _25654_, _03729_);
  or (_25656_, _25655_, _07390_);
  nor (_25657_, _25656_, _25642_);
  nor (_25659_, _25657_, _25639_);
  nor (_25660_, _25659_, _04481_);
  and (_25661_, _06637_, _05212_);
  nor (_25662_, _25629_, _07400_);
  not (_25663_, _25662_);
  nor (_25664_, _25663_, _25661_);
  nor (_25665_, _25664_, _03222_);
  not (_25666_, _25665_);
  nor (_25667_, _25666_, _25660_);
  nor (_25668_, _12519_, _10377_);
  nor (_25670_, _25668_, _25629_);
  nor (_25671_, _25670_, _03589_);
  or (_25672_, _25671_, _08828_);
  or (_25673_, _25672_, _25667_);
  and (_25674_, _12533_, _05212_);
  or (_25675_, _25629_, _07766_);
  or (_25676_, _25675_, _25674_);
  and (_25677_, _05212_, _06332_);
  nor (_25678_, _25677_, _25629_);
  and (_25679_, _25678_, _03601_);
  nor (_25681_, _25679_, _03780_);
  and (_25682_, _25681_, _25676_);
  and (_25683_, _25682_, _25673_);
  nor (_25684_, _25683_, _25635_);
  nor (_25685_, _25684_, _03622_);
  nor (_25686_, _25629_, _05718_);
  not (_25687_, _25686_);
  nor (_25688_, _25678_, _07777_);
  and (_25689_, _25688_, _25687_);
  nor (_25690_, _25689_, _25685_);
  nor (_25692_, _25690_, _03790_);
  nor (_25693_, _25641_, _06828_);
  and (_25694_, _25693_, _25687_);
  nor (_25695_, _25694_, _03624_);
  not (_25696_, _25695_);
  nor (_25697_, _25696_, _25692_);
  nor (_25698_, _12532_, _10377_);
  or (_25699_, _25629_, _07795_);
  nor (_25700_, _25699_, _25698_);
  or (_25701_, _25700_, _03785_);
  nor (_25703_, _25701_, _25697_);
  nor (_25704_, _25703_, _25632_);
  nor (_25705_, _25704_, _03815_);
  nor (_25706_, _25649_, _04246_);
  or (_25707_, _25706_, _03447_);
  nor (_25708_, _25707_, _25705_);
  and (_25709_, _12592_, _05212_);
  or (_25710_, _25629_, _03514_);
  nor (_25711_, _25710_, _25709_);
  nor (_25712_, _25711_, _25708_);
  or (_25714_, _25712_, _43004_);
  or (_25715_, _43000_, \oc8051_golden_model_1.PCON [2]);
  and (_25716_, _25715_, _41806_);
  and (_43581_, _25716_, _25714_);
  not (_25717_, \oc8051_golden_model_1.PCON [3]);
  nor (_25718_, _05212_, _25717_);
  nor (_25719_, _12738_, _10377_);
  nor (_25720_, _25719_, _25718_);
  nor (_25721_, _25720_, _07793_);
  and (_25722_, _12739_, _05212_);
  nor (_25724_, _25722_, _25718_);
  nor (_25725_, _25724_, _07778_);
  and (_25726_, _06592_, _05212_);
  or (_25727_, _25726_, _25718_);
  and (_25728_, _25727_, _04481_);
  and (_25729_, _05212_, \oc8051_golden_model_1.ACC [3]);
  nor (_25730_, _25729_, _25718_);
  nor (_25731_, _25730_, _03737_);
  nor (_25732_, _25730_, _09029_);
  nor (_25733_, _04409_, _25717_);
  or (_25734_, _25733_, _25732_);
  and (_25735_, _25734_, _04081_);
  nor (_25736_, _12627_, _10377_);
  nor (_25737_, _25736_, _25718_);
  nor (_25738_, _25737_, _04081_);
  or (_25739_, _25738_, _25735_);
  and (_25740_, _25739_, _03996_);
  nor (_25741_, _10377_, _05005_);
  nor (_25742_, _25741_, _25718_);
  nor (_25743_, _25742_, _03996_);
  nor (_25746_, _25743_, _25740_);
  nor (_25747_, _25746_, _03729_);
  or (_25748_, _25747_, _07390_);
  nor (_25749_, _25748_, _25731_);
  and (_25750_, _25742_, _07390_);
  or (_25751_, _25750_, _04481_);
  nor (_25752_, _25751_, _25749_);
  or (_25753_, _25752_, _25728_);
  and (_25754_, _25753_, _03589_);
  nor (_25755_, _12718_, _10377_);
  nor (_25757_, _25755_, _25718_);
  nor (_25758_, _25757_, _03589_);
  or (_25759_, _25758_, _08828_);
  or (_25760_, _25759_, _25754_);
  and (_25761_, _12733_, _05212_);
  or (_25762_, _25718_, _07766_);
  or (_25763_, _25762_, _25761_);
  and (_25764_, _05212_, _06276_);
  nor (_25765_, _25764_, _25718_);
  and (_25766_, _25765_, _03601_);
  nor (_25768_, _25766_, _03780_);
  and (_25769_, _25768_, _25763_);
  and (_25770_, _25769_, _25760_);
  nor (_25771_, _25770_, _25725_);
  nor (_25772_, _25771_, _03622_);
  nor (_25773_, _25718_, _05567_);
  not (_25774_, _25773_);
  nor (_25775_, _25765_, _07777_);
  and (_25776_, _25775_, _25774_);
  nor (_25777_, _25776_, _25772_);
  nor (_25779_, _25777_, _03790_);
  nor (_25780_, _25730_, _06828_);
  and (_25781_, _25780_, _25774_);
  or (_25782_, _25781_, _25779_);
  and (_25783_, _25782_, _07795_);
  nor (_25784_, _12732_, _10377_);
  nor (_25785_, _25784_, _25718_);
  nor (_25786_, _25785_, _07795_);
  or (_25787_, _25786_, _25783_);
  and (_25788_, _25787_, _07793_);
  nor (_25790_, _25788_, _25721_);
  nor (_25791_, _25790_, _03815_);
  nor (_25792_, _25737_, _04246_);
  or (_25793_, _25792_, _03447_);
  nor (_25794_, _25793_, _25791_);
  and (_25795_, _12794_, _05212_);
  nor (_25796_, _25795_, _25718_);
  and (_25797_, _25796_, _03447_);
  nor (_25798_, _25797_, _25794_);
  or (_25799_, _25798_, _43004_);
  or (_25801_, _43000_, \oc8051_golden_model_1.PCON [3]);
  and (_25802_, _25801_, _41806_);
  and (_43582_, _25802_, _25799_);
  not (_25803_, \oc8051_golden_model_1.PCON [4]);
  nor (_25804_, _05212_, _25803_);
  nor (_25805_, _12816_, _10377_);
  nor (_25806_, _25805_, _25804_);
  nor (_25807_, _25806_, _07793_);
  and (_25808_, _12817_, _05212_);
  nor (_25809_, _25808_, _25804_);
  nor (_25811_, _25809_, _07778_);
  and (_25812_, _06298_, _05212_);
  nor (_25813_, _25812_, _25804_);
  and (_25814_, _25813_, _03601_);
  and (_25815_, _05212_, \oc8051_golden_model_1.ACC [4]);
  nor (_25816_, _25815_, _25804_);
  nor (_25817_, _25816_, _03737_);
  nor (_25818_, _25816_, _09029_);
  nor (_25819_, _04409_, _25803_);
  or (_25820_, _25819_, _25818_);
  and (_25822_, _25820_, _04081_);
  nor (_25823_, _12841_, _10377_);
  nor (_25824_, _25823_, _25804_);
  nor (_25825_, _25824_, _04081_);
  or (_25826_, _25825_, _25822_);
  and (_25827_, _25826_, _03996_);
  nor (_25828_, _05777_, _10377_);
  nor (_25829_, _25828_, _25804_);
  nor (_25830_, _25829_, _03996_);
  nor (_25831_, _25830_, _25827_);
  nor (_25833_, _25831_, _03729_);
  or (_25834_, _25833_, _07390_);
  nor (_25835_, _25834_, _25817_);
  and (_25836_, _25829_, _07390_);
  nor (_25837_, _25836_, _25835_);
  nor (_25838_, _25837_, _04481_);
  and (_25839_, _06730_, _05212_);
  nor (_25840_, _25804_, _07400_);
  not (_25841_, _25840_);
  nor (_25842_, _25841_, _25839_);
  or (_25844_, _25842_, _03222_);
  nor (_25845_, _25844_, _25838_);
  nor (_25846_, _12933_, _10377_);
  nor (_25847_, _25846_, _25804_);
  nor (_25848_, _25847_, _03589_);
  or (_25849_, _25848_, _03601_);
  nor (_25850_, _25849_, _25845_);
  nor (_25851_, _25850_, _25814_);
  or (_25852_, _25851_, _03600_);
  and (_25853_, _12821_, _05212_);
  or (_25855_, _25853_, _25804_);
  or (_25856_, _25855_, _07766_);
  and (_25857_, _25856_, _07778_);
  and (_25858_, _25857_, _25852_);
  nor (_25859_, _25858_, _25811_);
  nor (_25860_, _25859_, _03622_);
  nor (_25861_, _25804_, _05825_);
  not (_25862_, _25861_);
  nor (_25863_, _25813_, _07777_);
  and (_25864_, _25863_, _25862_);
  nor (_25866_, _25864_, _25860_);
  nor (_25867_, _25866_, _03790_);
  nor (_25868_, _25816_, _06828_);
  and (_25869_, _25868_, _25862_);
  or (_25870_, _25869_, _25867_);
  and (_25871_, _25870_, _07795_);
  nor (_25872_, _12819_, _10377_);
  nor (_25873_, _25872_, _25804_);
  nor (_25874_, _25873_, _07795_);
  or (_25875_, _25874_, _25871_);
  and (_25877_, _25875_, _07793_);
  nor (_25878_, _25877_, _25807_);
  nor (_25879_, _25878_, _03815_);
  nor (_25880_, _25824_, _04246_);
  or (_25881_, _25880_, _03447_);
  nor (_25882_, _25881_, _25879_);
  and (_25883_, _13003_, _05212_);
  or (_25884_, _25804_, _03514_);
  nor (_25885_, _25884_, _25883_);
  nor (_25886_, _25885_, _25882_);
  or (_25888_, _25886_, _43004_);
  or (_25889_, _43000_, \oc8051_golden_model_1.PCON [4]);
  and (_25890_, _25889_, _41806_);
  and (_43583_, _25890_, _25888_);
  not (_25891_, \oc8051_golden_model_1.PCON [5]);
  nor (_25892_, _05212_, _25891_);
  nor (_25893_, _13146_, _10377_);
  nor (_25894_, _25893_, _25892_);
  nor (_25895_, _25894_, _07793_);
  and (_25896_, _13147_, _05212_);
  nor (_25898_, _25896_, _25892_);
  nor (_25899_, _25898_, _07778_);
  and (_25900_, _06684_, _05212_);
  or (_25901_, _25900_, _25892_);
  and (_25902_, _25901_, _04481_);
  and (_25903_, _05212_, \oc8051_golden_model_1.ACC [5]);
  nor (_25904_, _25903_, _25892_);
  nor (_25905_, _25904_, _03737_);
  nor (_25906_, _25904_, _09029_);
  nor (_25907_, _04409_, _25891_);
  or (_25909_, _25907_, _25906_);
  and (_25910_, _25909_, _04081_);
  nor (_25911_, _13014_, _10377_);
  nor (_25912_, _25911_, _25892_);
  nor (_25913_, _25912_, _04081_);
  or (_25914_, _25913_, _25910_);
  and (_25915_, _25914_, _03996_);
  nor (_25916_, _05469_, _10377_);
  nor (_25917_, _25916_, _25892_);
  nor (_25918_, _25917_, _03996_);
  nor (_25920_, _25918_, _25915_);
  nor (_25921_, _25920_, _03729_);
  or (_25922_, _25921_, _07390_);
  nor (_25923_, _25922_, _25905_);
  and (_25924_, _25917_, _07390_);
  or (_25925_, _25924_, _04481_);
  nor (_25926_, _25925_, _25923_);
  or (_25927_, _25926_, _25902_);
  and (_25928_, _25927_, _03589_);
  nor (_25929_, _13127_, _10377_);
  nor (_25931_, _25929_, _25892_);
  nor (_25932_, _25931_, _03589_);
  or (_25933_, _25932_, _08828_);
  or (_25934_, _25933_, _25928_);
  and (_25935_, _13141_, _05212_);
  or (_25936_, _25892_, _07766_);
  or (_25937_, _25936_, _25935_);
  and (_25938_, _06306_, _05212_);
  nor (_25939_, _25938_, _25892_);
  and (_25940_, _25939_, _03601_);
  nor (_25942_, _25940_, _03780_);
  and (_25943_, _25942_, _25937_);
  and (_25944_, _25943_, _25934_);
  nor (_25945_, _25944_, _25899_);
  nor (_25946_, _25945_, _03622_);
  nor (_25947_, _25892_, _05518_);
  not (_25948_, _25947_);
  nor (_25949_, _25939_, _07777_);
  and (_25950_, _25949_, _25948_);
  nor (_25951_, _25950_, _25946_);
  nor (_25953_, _25951_, _03790_);
  nor (_25954_, _25904_, _06828_);
  and (_25955_, _25954_, _25948_);
  nor (_25956_, _25955_, _03624_);
  not (_25957_, _25956_);
  nor (_25958_, _25957_, _25953_);
  nor (_25959_, _13140_, _10377_);
  or (_25960_, _25892_, _07795_);
  nor (_25961_, _25960_, _25959_);
  or (_25962_, _25961_, _03785_);
  nor (_25964_, _25962_, _25958_);
  nor (_25965_, _25964_, _25895_);
  nor (_25966_, _25965_, _03815_);
  nor (_25967_, _25912_, _04246_);
  or (_25968_, _25967_, _03447_);
  nor (_25969_, _25968_, _25966_);
  and (_25970_, _13199_, _05212_);
  or (_25971_, _25892_, _03514_);
  nor (_25972_, _25971_, _25970_);
  nor (_25973_, _25972_, _25969_);
  or (_25975_, _25973_, _43004_);
  or (_25976_, _43000_, \oc8051_golden_model_1.PCON [5]);
  and (_25977_, _25976_, _41806_);
  and (_43584_, _25977_, _25975_);
  not (_25978_, \oc8051_golden_model_1.PCON [6]);
  nor (_25979_, _05212_, _25978_);
  nor (_25980_, _13352_, _10377_);
  nor (_25981_, _25980_, _25979_);
  nor (_25982_, _25981_, _07793_);
  and (_25983_, _13353_, _05212_);
  nor (_25985_, _25983_, _25979_);
  nor (_25986_, _25985_, _07778_);
  and (_25987_, _06455_, _05212_);
  or (_25988_, _25987_, _25979_);
  and (_25989_, _25988_, _04481_);
  and (_25990_, _05212_, \oc8051_golden_model_1.ACC [6]);
  nor (_25991_, _25990_, _25979_);
  nor (_25992_, _25991_, _03737_);
  nor (_25993_, _25991_, _09029_);
  nor (_25994_, _04409_, _25978_);
  or (_25996_, _25994_, _25993_);
  and (_25997_, _25996_, _04081_);
  nor (_25998_, _13242_, _10377_);
  nor (_25999_, _25998_, _25979_);
  nor (_26000_, _25999_, _04081_);
  or (_26001_, _26000_, _25997_);
  and (_26002_, _26001_, _03996_);
  nor (_26003_, _05363_, _10377_);
  nor (_26004_, _26003_, _25979_);
  nor (_26005_, _26004_, _03996_);
  nor (_26007_, _26005_, _26002_);
  nor (_26008_, _26007_, _03729_);
  or (_26009_, _26008_, _07390_);
  nor (_26010_, _26009_, _25992_);
  and (_26011_, _26004_, _07390_);
  or (_26012_, _26011_, _04481_);
  nor (_26013_, _26012_, _26010_);
  or (_26014_, _26013_, _25989_);
  and (_26015_, _26014_, _03589_);
  nor (_26016_, _13332_, _10377_);
  nor (_26018_, _26016_, _25979_);
  nor (_26019_, _26018_, _03589_);
  or (_26020_, _26019_, _08828_);
  or (_26021_, _26020_, _26015_);
  and (_26022_, _13347_, _05212_);
  or (_26023_, _25979_, _07766_);
  or (_26024_, _26023_, _26022_);
  and (_26025_, _13339_, _05212_);
  nor (_26026_, _26025_, _25979_);
  and (_26027_, _26026_, _03601_);
  nor (_26029_, _26027_, _03780_);
  and (_26030_, _26029_, _26024_);
  and (_26031_, _26030_, _26021_);
  nor (_26032_, _26031_, _25986_);
  nor (_26033_, _26032_, _03622_);
  nor (_26034_, _25979_, _05412_);
  not (_26035_, _26034_);
  nor (_26036_, _26026_, _07777_);
  and (_26037_, _26036_, _26035_);
  nor (_26038_, _26037_, _26033_);
  nor (_26040_, _26038_, _03790_);
  nor (_26041_, _25991_, _06828_);
  and (_26042_, _26041_, _26035_);
  or (_26043_, _26042_, _26040_);
  and (_26044_, _26043_, _07795_);
  nor (_26045_, _13346_, _10377_);
  nor (_26046_, _26045_, _25979_);
  nor (_26047_, _26046_, _07795_);
  or (_26048_, _26047_, _26044_);
  and (_26049_, _26048_, _07793_);
  nor (_26051_, _26049_, _25982_);
  nor (_26052_, _26051_, _03815_);
  nor (_26053_, _25999_, _04246_);
  or (_26054_, _26053_, _03447_);
  nor (_26055_, _26054_, _26052_);
  and (_26056_, _13402_, _05212_);
  or (_26057_, _25979_, _03514_);
  nor (_26058_, _26057_, _26056_);
  nor (_26059_, _26058_, _26055_);
  or (_26060_, _26059_, _43004_);
  or (_26062_, _43000_, \oc8051_golden_model_1.PCON [6]);
  and (_26063_, _26062_, _41806_);
  and (_43585_, _26063_, _26060_);
  not (_26064_, \oc8051_golden_model_1.SBUF [0]);
  nor (_26065_, _05221_, _26064_);
  nor (_26066_, _05666_, _10458_);
  nor (_26067_, _26066_, _26065_);
  and (_26068_, _26067_, _17166_);
  and (_26069_, _05221_, \oc8051_golden_model_1.ACC [0]);
  nor (_26070_, _26069_, _26065_);
  nor (_26072_, _26070_, _03737_);
  nor (_26073_, _26072_, _07390_);
  nor (_26074_, _26067_, _04081_);
  nor (_26075_, _04409_, _26064_);
  nor (_26076_, _26070_, _09029_);
  nor (_26077_, _26076_, _26075_);
  nor (_26078_, _26077_, _03610_);
  or (_26079_, _26078_, _03723_);
  nor (_26080_, _26079_, _26074_);
  or (_26081_, _26080_, _03729_);
  and (_26082_, _26081_, _26073_);
  and (_26083_, _05221_, _04620_);
  or (_26084_, _26065_, _25480_);
  nor (_26085_, _26084_, _26083_);
  nor (_26086_, _26085_, _26082_);
  nor (_26087_, _26086_, _04481_);
  and (_26088_, _06546_, _05221_);
  nor (_26089_, _26065_, _07400_);
  not (_26090_, _26089_);
  nor (_26091_, _26090_, _26088_);
  nor (_26094_, _26091_, _26087_);
  nor (_26095_, _26094_, _03222_);
  nor (_26096_, _12109_, _10458_);
  or (_26097_, _26065_, _03589_);
  nor (_26098_, _26097_, _26096_);
  or (_26099_, _26098_, _03601_);
  nor (_26100_, _26099_, _26095_);
  and (_26101_, _05221_, _06274_);
  nor (_26102_, _26101_, _26065_);
  nand (_26103_, _26102_, _07766_);
  and (_26105_, _26103_, _08828_);
  nor (_26106_, _26105_, _26100_);
  and (_26107_, _12124_, _05221_);
  nor (_26108_, _26107_, _26065_);
  and (_26109_, _26108_, _03600_);
  nor (_26110_, _26109_, _26106_);
  nor (_26111_, _26110_, _03780_);
  and (_26112_, _12128_, _05221_);
  or (_26113_, _26065_, _07778_);
  nor (_26114_, _26113_, _26112_);
  or (_26116_, _26114_, _03622_);
  nor (_26117_, _26116_, _26111_);
  or (_26118_, _26102_, _07777_);
  nor (_26119_, _26118_, _26066_);
  nor (_26120_, _26119_, _26117_);
  nor (_26121_, _26120_, _03790_);
  nor (_26122_, _26065_, _05666_);
  or (_26123_, _26122_, _06828_);
  nor (_26124_, _26123_, _26070_);
  or (_26125_, _26124_, _26121_);
  and (_26127_, _26125_, _07795_);
  nor (_26128_, _12122_, _10458_);
  nor (_26129_, _26128_, _26065_);
  nor (_26130_, _26129_, _07795_);
  or (_26131_, _26130_, _26127_);
  and (_26132_, _26131_, _07793_);
  nor (_26133_, _12003_, _10458_);
  nor (_26134_, _26133_, _26065_);
  nor (_26135_, _26134_, _07793_);
  nor (_26136_, _26135_, _17166_);
  not (_26138_, _26136_);
  nor (_26139_, _26138_, _26132_);
  nor (_26140_, _26139_, _26068_);
  or (_26141_, _26140_, _43004_);
  or (_26142_, _43000_, \oc8051_golden_model_1.SBUF [0]);
  and (_26143_, _26142_, _41806_);
  and (_43588_, _26143_, _26141_);
  and (_26144_, _06501_, _05221_);
  not (_26145_, \oc8051_golden_model_1.SBUF [1]);
  nor (_26146_, _05221_, _26145_);
  nor (_26148_, _26146_, _07400_);
  not (_26149_, _26148_);
  nor (_26150_, _26149_, _26144_);
  not (_26151_, _26150_);
  and (_26152_, _05221_, _06764_);
  nor (_26153_, _26152_, _26146_);
  and (_26154_, _26153_, _07390_);
  nor (_26155_, _05221_, \oc8051_golden_model_1.SBUF [1]);
  and (_26156_, _05221_, _03274_);
  nor (_26157_, _26156_, _26155_);
  and (_26159_, _26157_, _03729_);
  and (_26160_, _26157_, _04409_);
  nor (_26161_, _04409_, _26145_);
  or (_26162_, _26161_, _26160_);
  and (_26163_, _26162_, _04081_);
  and (_26164_, _12213_, _05221_);
  nor (_26165_, _26164_, _26155_);
  and (_26166_, _26165_, _03610_);
  or (_26167_, _26166_, _26163_);
  and (_26168_, _26167_, _03996_);
  nor (_26170_, _26153_, _03996_);
  nor (_26171_, _26170_, _26168_);
  nor (_26172_, _26171_, _03729_);
  or (_26173_, _26172_, _07390_);
  nor (_26174_, _26173_, _26159_);
  nor (_26175_, _26174_, _26154_);
  nor (_26176_, _26175_, _04481_);
  nor (_26177_, _26176_, _03222_);
  and (_26178_, _26177_, _26151_);
  not (_26179_, _26155_);
  and (_26181_, _12313_, _05221_);
  nor (_26182_, _26181_, _03589_);
  and (_26183_, _26182_, _26179_);
  nor (_26184_, _26183_, _26178_);
  nor (_26185_, _26184_, _08828_);
  nor (_26186_, _12327_, _10458_);
  nor (_26187_, _26186_, _07766_);
  and (_26188_, _05221_, _04303_);
  nor (_26189_, _26188_, _05886_);
  nor (_26190_, _26189_, _26187_);
  nor (_26191_, _26190_, _26155_);
  nor (_26192_, _26191_, _26185_);
  nor (_26193_, _26192_, _03780_);
  nor (_26194_, _12333_, _10458_);
  nor (_26195_, _26194_, _07778_);
  and (_26196_, _26195_, _26179_);
  nor (_26197_, _26196_, _26193_);
  nor (_26198_, _26197_, _03622_);
  nor (_26199_, _12207_, _10458_);
  nor (_26200_, _26199_, _07777_);
  and (_26203_, _26200_, _26179_);
  nor (_26204_, _26203_, _26198_);
  nor (_26205_, _26204_, _03790_);
  nor (_26206_, _26146_, _05618_);
  nor (_26207_, _26206_, _06828_);
  and (_26208_, _26207_, _26157_);
  nor (_26209_, _26208_, _26205_);
  or (_26210_, _26209_, _18499_);
  and (_26211_, _26188_, _05617_);
  nor (_26212_, _26211_, _07795_);
  and (_26214_, _26212_, _26179_);
  nand (_26215_, _26156_, _05617_);
  nor (_26216_, _26155_, _07793_);
  and (_26217_, _26216_, _26215_);
  or (_26218_, _26217_, _03815_);
  nor (_26219_, _26218_, _26214_);
  and (_26220_, _26219_, _26210_);
  nor (_26221_, _26165_, _04246_);
  nor (_26222_, _26221_, _26220_);
  and (_26223_, _26222_, _03514_);
  nor (_26225_, _26164_, _26146_);
  nor (_26226_, _26225_, _03514_);
  or (_26227_, _26226_, _26223_);
  or (_26228_, _26227_, _43004_);
  or (_26229_, _43000_, \oc8051_golden_model_1.SBUF [1]);
  and (_26230_, _26229_, _41806_);
  and (_43589_, _26230_, _26228_);
  not (_26231_, \oc8051_golden_model_1.SBUF [2]);
  nor (_26232_, _05221_, _26231_);
  nor (_26233_, _12538_, _10458_);
  nor (_26235_, _26233_, _26232_);
  nor (_26236_, _26235_, _07793_);
  and (_26237_, _12539_, _05221_);
  nor (_26238_, _26237_, _26232_);
  nor (_26239_, _26238_, _07778_);
  nor (_26240_, _10458_, _04875_);
  nor (_26241_, _26240_, _26232_);
  and (_26242_, _26241_, _07390_);
  and (_26243_, _05221_, \oc8051_golden_model_1.ACC [2]);
  nor (_26244_, _26243_, _26232_);
  nor (_26246_, _26244_, _03737_);
  nor (_26247_, _26244_, _09029_);
  nor (_26248_, _04409_, _26231_);
  or (_26249_, _26248_, _26247_);
  and (_26250_, _26249_, _04081_);
  nor (_26251_, _12416_, _10458_);
  nor (_26252_, _26251_, _26232_);
  nor (_26253_, _26252_, _04081_);
  or (_26254_, _26253_, _26250_);
  and (_26255_, _26254_, _03996_);
  nor (_26257_, _26241_, _03996_);
  nor (_26258_, _26257_, _26255_);
  nor (_26259_, _26258_, _03729_);
  or (_26260_, _26259_, _07390_);
  nor (_26261_, _26260_, _26246_);
  nor (_26262_, _26261_, _26242_);
  nor (_26263_, _26262_, _04481_);
  and (_26264_, _06637_, _05221_);
  nor (_26265_, _26232_, _07400_);
  not (_26266_, _26265_);
  nor (_26268_, _26266_, _26264_);
  nor (_26269_, _26268_, _03222_);
  not (_26270_, _26269_);
  nor (_26271_, _26270_, _26263_);
  nor (_26272_, _12519_, _10458_);
  nor (_26273_, _26272_, _26232_);
  nor (_26274_, _26273_, _03589_);
  or (_26275_, _26274_, _08828_);
  or (_26276_, _26275_, _26271_);
  and (_26277_, _12533_, _05221_);
  or (_26279_, _26232_, _07766_);
  or (_26280_, _26279_, _26277_);
  and (_26281_, _05221_, _06332_);
  nor (_26282_, _26281_, _26232_);
  and (_26283_, _26282_, _03601_);
  nor (_26284_, _26283_, _03780_);
  and (_26285_, _26284_, _26280_);
  and (_26286_, _26285_, _26276_);
  nor (_26287_, _26286_, _26239_);
  nor (_26288_, _26287_, _03622_);
  nor (_26290_, _26232_, _05718_);
  not (_26291_, _26290_);
  nor (_26292_, _26282_, _07777_);
  and (_26293_, _26292_, _26291_);
  nor (_26294_, _26293_, _26288_);
  nor (_26295_, _26294_, _03790_);
  nor (_26296_, _26244_, _06828_);
  and (_26297_, _26296_, _26291_);
  nor (_26298_, _26297_, _03624_);
  not (_26299_, _26298_);
  nor (_26301_, _26299_, _26295_);
  nor (_26302_, _12532_, _10458_);
  or (_26303_, _26232_, _07795_);
  nor (_26304_, _26303_, _26302_);
  or (_26305_, _26304_, _03785_);
  nor (_26306_, _26305_, _26301_);
  nor (_26307_, _26306_, _26236_);
  nor (_26308_, _26307_, _03815_);
  nor (_26309_, _26252_, _04246_);
  or (_26310_, _26309_, _03447_);
  nor (_26312_, _26310_, _26308_);
  and (_26313_, _12592_, _05221_);
  or (_26314_, _26232_, _03514_);
  nor (_26315_, _26314_, _26313_);
  nor (_26316_, _26315_, _26312_);
  or (_26317_, _26316_, _43004_);
  or (_26318_, _43000_, \oc8051_golden_model_1.SBUF [2]);
  and (_26319_, _26318_, _41806_);
  and (_43590_, _26319_, _26317_);
  not (_26320_, \oc8051_golden_model_1.SBUF [3]);
  nor (_26322_, _05221_, _26320_);
  nor (_26323_, _12738_, _10458_);
  nor (_26324_, _26323_, _26322_);
  nor (_26325_, _26324_, _07793_);
  and (_26326_, _12739_, _05221_);
  nor (_26327_, _26326_, _26322_);
  nor (_26328_, _26327_, _07778_);
  and (_26329_, _06592_, _05221_);
  or (_26330_, _26329_, _26322_);
  and (_26331_, _26330_, _04481_);
  and (_26333_, _05221_, \oc8051_golden_model_1.ACC [3]);
  nor (_26334_, _26333_, _26322_);
  nor (_26335_, _26334_, _03737_);
  nor (_26336_, _26334_, _09029_);
  nor (_26337_, _04409_, _26320_);
  or (_26338_, _26337_, _26336_);
  and (_26339_, _26338_, _04081_);
  nor (_26340_, _12627_, _10458_);
  nor (_26341_, _26340_, _26322_);
  nor (_26342_, _26341_, _04081_);
  or (_26344_, _26342_, _26339_);
  and (_26345_, _26344_, _03996_);
  nor (_26346_, _10458_, _05005_);
  nor (_26347_, _26346_, _26322_);
  nor (_26348_, _26347_, _03996_);
  nor (_26349_, _26348_, _26345_);
  nor (_26350_, _26349_, _03729_);
  or (_26351_, _26350_, _07390_);
  nor (_26352_, _26351_, _26335_);
  and (_26353_, _26347_, _07390_);
  or (_26355_, _26353_, _04481_);
  nor (_26356_, _26355_, _26352_);
  or (_26357_, _26356_, _26331_);
  and (_26358_, _26357_, _03589_);
  nor (_26359_, _12718_, _10458_);
  nor (_26360_, _26359_, _26322_);
  nor (_26361_, _26360_, _03589_);
  or (_26362_, _26361_, _08828_);
  or (_26363_, _26362_, _26358_);
  and (_26364_, _12733_, _05221_);
  or (_26366_, _26322_, _07766_);
  or (_26367_, _26366_, _26364_);
  and (_26368_, _05221_, _06276_);
  nor (_26369_, _26368_, _26322_);
  and (_26370_, _26369_, _03601_);
  nor (_26371_, _26370_, _03780_);
  and (_26372_, _26371_, _26367_);
  and (_26373_, _26372_, _26363_);
  nor (_26374_, _26373_, _26328_);
  nor (_26375_, _26374_, _03622_);
  nor (_26377_, _26322_, _05567_);
  not (_26378_, _26377_);
  nor (_26379_, _26369_, _07777_);
  and (_26380_, _26379_, _26378_);
  nor (_26381_, _26380_, _26375_);
  nor (_26382_, _26381_, _03790_);
  nor (_26383_, _26334_, _06828_);
  and (_26384_, _26383_, _26378_);
  nor (_26385_, _26384_, _03624_);
  not (_26386_, _26385_);
  nor (_26388_, _26386_, _26382_);
  nor (_26389_, _12732_, _10458_);
  or (_26390_, _26322_, _07795_);
  nor (_26391_, _26390_, _26389_);
  or (_26392_, _26391_, _03785_);
  nor (_26393_, _26392_, _26388_);
  nor (_26394_, _26393_, _26325_);
  nor (_26395_, _26394_, _03815_);
  nor (_26396_, _26341_, _04246_);
  or (_26397_, _26396_, _03447_);
  nor (_26399_, _26397_, _26395_);
  and (_26400_, _12794_, _05221_);
  or (_26401_, _26322_, _03514_);
  nor (_26402_, _26401_, _26400_);
  nor (_26403_, _26402_, _26399_);
  or (_26404_, _26403_, _43004_);
  or (_26405_, _43000_, \oc8051_golden_model_1.SBUF [3]);
  and (_26406_, _26405_, _41806_);
  and (_43591_, _26406_, _26404_);
  not (_26407_, \oc8051_golden_model_1.SBUF [4]);
  nor (_26409_, _05221_, _26407_);
  nor (_26410_, _12816_, _10458_);
  nor (_26411_, _26410_, _26409_);
  nor (_26412_, _26411_, _07793_);
  and (_26413_, _12817_, _05221_);
  nor (_26414_, _26413_, _26409_);
  nor (_26415_, _26414_, _07778_);
  and (_26416_, _06298_, _05221_);
  nor (_26417_, _26416_, _26409_);
  and (_26418_, _26417_, _03601_);
  nor (_26420_, _05777_, _10458_);
  nor (_26421_, _26420_, _26409_);
  and (_26422_, _26421_, _07390_);
  and (_26423_, _05221_, \oc8051_golden_model_1.ACC [4]);
  nor (_26424_, _26423_, _26409_);
  nor (_26425_, _26424_, _03737_);
  nor (_26426_, _26424_, _09029_);
  nor (_26427_, _04409_, _26407_);
  or (_26428_, _26427_, _26426_);
  and (_26429_, _26428_, _04081_);
  nor (_26431_, _12841_, _10458_);
  nor (_26432_, _26431_, _26409_);
  nor (_26433_, _26432_, _04081_);
  or (_26434_, _26433_, _26429_);
  and (_26435_, _26434_, _03996_);
  nor (_26436_, _26421_, _03996_);
  nor (_26437_, _26436_, _26435_);
  nor (_26438_, _26437_, _03729_);
  or (_26439_, _26438_, _07390_);
  nor (_26440_, _26439_, _26425_);
  nor (_26442_, _26440_, _26422_);
  nor (_26443_, _26442_, _04481_);
  and (_26444_, _06730_, _05221_);
  nor (_26445_, _26409_, _07400_);
  not (_26446_, _26445_);
  nor (_26447_, _26446_, _26444_);
  or (_26448_, _26447_, _03222_);
  nor (_26449_, _26448_, _26443_);
  nor (_26450_, _12933_, _10458_);
  nor (_26451_, _26450_, _26409_);
  nor (_26453_, _26451_, _03589_);
  or (_26454_, _26453_, _03601_);
  nor (_26455_, _26454_, _26449_);
  nor (_26456_, _26455_, _26418_);
  or (_26457_, _26456_, _03600_);
  and (_26458_, _12821_, _05221_);
  or (_26459_, _26458_, _26409_);
  or (_26460_, _26459_, _07766_);
  and (_26461_, _26460_, _07778_);
  and (_26462_, _26461_, _26457_);
  nor (_26464_, _26462_, _26415_);
  nor (_26465_, _26464_, _03622_);
  nor (_26466_, _26409_, _05825_);
  not (_26467_, _26466_);
  nor (_26468_, _26417_, _07777_);
  and (_26469_, _26468_, _26467_);
  nor (_26470_, _26469_, _26465_);
  nor (_26471_, _26470_, _03790_);
  nor (_26472_, _26424_, _06828_);
  and (_26473_, _26472_, _26467_);
  nor (_26475_, _26473_, _03624_);
  not (_26476_, _26475_);
  nor (_26477_, _26476_, _26471_);
  nor (_26478_, _12819_, _10458_);
  or (_26479_, _26409_, _07795_);
  nor (_26480_, _26479_, _26478_);
  or (_26481_, _26480_, _03785_);
  nor (_26482_, _26481_, _26477_);
  nor (_26483_, _26482_, _26412_);
  nor (_26484_, _26483_, _03815_);
  nor (_26486_, _26432_, _04246_);
  or (_26487_, _26486_, _03447_);
  nor (_26488_, _26487_, _26484_);
  and (_26489_, _13003_, _05221_);
  or (_26490_, _26409_, _03514_);
  nor (_26491_, _26490_, _26489_);
  nor (_26492_, _26491_, _26488_);
  or (_26493_, _26492_, _43004_);
  or (_26494_, _43000_, \oc8051_golden_model_1.SBUF [4]);
  and (_26495_, _26494_, _41806_);
  and (_43592_, _26495_, _26493_);
  not (_26497_, \oc8051_golden_model_1.SBUF [5]);
  nor (_26498_, _05221_, _26497_);
  nor (_26499_, _13146_, _10458_);
  nor (_26500_, _26499_, _26498_);
  nor (_26501_, _26500_, _07793_);
  and (_26502_, _13147_, _05221_);
  nor (_26503_, _26502_, _26498_);
  nor (_26504_, _26503_, _07778_);
  and (_26505_, _06684_, _05221_);
  or (_26507_, _26505_, _26498_);
  and (_26508_, _26507_, _04481_);
  and (_26509_, _05221_, \oc8051_golden_model_1.ACC [5]);
  nor (_26510_, _26509_, _26498_);
  nor (_26511_, _26510_, _03737_);
  nor (_26512_, _26510_, _09029_);
  nor (_26513_, _04409_, _26497_);
  or (_26514_, _26513_, _26512_);
  and (_26515_, _26514_, _04081_);
  nor (_26516_, _13014_, _10458_);
  nor (_26518_, _26516_, _26498_);
  nor (_26519_, _26518_, _04081_);
  or (_26520_, _26519_, _26515_);
  and (_26521_, _26520_, _03996_);
  nor (_26522_, _05469_, _10458_);
  nor (_26523_, _26522_, _26498_);
  nor (_26524_, _26523_, _03996_);
  nor (_26525_, _26524_, _26521_);
  nor (_26526_, _26525_, _03729_);
  or (_26527_, _26526_, _07390_);
  nor (_26529_, _26527_, _26511_);
  and (_26530_, _26523_, _07390_);
  or (_26531_, _26530_, _04481_);
  nor (_26532_, _26531_, _26529_);
  or (_26533_, _26532_, _26508_);
  and (_26534_, _26533_, _03589_);
  nor (_26535_, _13127_, _10458_);
  nor (_26536_, _26535_, _26498_);
  nor (_26537_, _26536_, _03589_);
  or (_26538_, _26537_, _08828_);
  or (_26540_, _26538_, _26534_);
  and (_26541_, _13141_, _05221_);
  or (_26542_, _26498_, _07766_);
  or (_26543_, _26542_, _26541_);
  and (_26544_, _06306_, _05221_);
  nor (_26545_, _26544_, _26498_);
  and (_26546_, _26545_, _03601_);
  nor (_26547_, _26546_, _03780_);
  and (_26548_, _26547_, _26543_);
  and (_26549_, _26548_, _26540_);
  nor (_26551_, _26549_, _26504_);
  nor (_26552_, _26551_, _03622_);
  nor (_26553_, _26498_, _05518_);
  not (_26554_, _26553_);
  nor (_26555_, _26545_, _07777_);
  and (_26556_, _26555_, _26554_);
  nor (_26557_, _26556_, _26552_);
  nor (_26558_, _26557_, _03790_);
  nor (_26559_, _26510_, _06828_);
  and (_26560_, _26559_, _26554_);
  nor (_26562_, _26560_, _03624_);
  not (_26563_, _26562_);
  nor (_26564_, _26563_, _26558_);
  nor (_26565_, _13140_, _10458_);
  or (_26566_, _26498_, _07795_);
  nor (_26567_, _26566_, _26565_);
  or (_26568_, _26567_, _03785_);
  nor (_26569_, _26568_, _26564_);
  nor (_26570_, _26569_, _26501_);
  nor (_26571_, _26570_, _03815_);
  nor (_26573_, _26518_, _04246_);
  or (_26574_, _26573_, _03447_);
  nor (_26575_, _26574_, _26571_);
  and (_26576_, _13199_, _05221_);
  or (_26577_, _26498_, _03514_);
  nor (_26578_, _26577_, _26576_);
  nor (_26579_, _26578_, _26575_);
  or (_26580_, _26579_, _43004_);
  or (_26581_, _43000_, \oc8051_golden_model_1.SBUF [5]);
  and (_26582_, _26581_, _41806_);
  and (_43594_, _26582_, _26580_);
  not (_26584_, \oc8051_golden_model_1.SBUF [6]);
  nor (_26585_, _05221_, _26584_);
  nor (_26586_, _13352_, _10458_);
  nor (_26587_, _26586_, _26585_);
  nor (_26588_, _26587_, _07793_);
  and (_26589_, _13353_, _05221_);
  nor (_26590_, _26589_, _26585_);
  nor (_26591_, _26590_, _07778_);
  and (_26592_, _06455_, _05221_);
  or (_26594_, _26592_, _26585_);
  and (_26595_, _26594_, _04481_);
  and (_26596_, _05221_, \oc8051_golden_model_1.ACC [6]);
  nor (_26597_, _26596_, _26585_);
  nor (_26598_, _26597_, _03737_);
  nor (_26599_, _26597_, _09029_);
  nor (_26600_, _04409_, _26584_);
  or (_26601_, _26600_, _26599_);
  and (_26602_, _26601_, _04081_);
  nor (_26603_, _13242_, _10458_);
  nor (_26605_, _26603_, _26585_);
  nor (_26606_, _26605_, _04081_);
  or (_26607_, _26606_, _26602_);
  and (_26608_, _26607_, _03996_);
  nor (_26609_, _05363_, _10458_);
  nor (_26610_, _26609_, _26585_);
  nor (_26611_, _26610_, _03996_);
  nor (_26612_, _26611_, _26608_);
  nor (_26613_, _26612_, _03729_);
  or (_26614_, _26613_, _07390_);
  nor (_26616_, _26614_, _26598_);
  and (_26617_, _26610_, _07390_);
  or (_26618_, _26617_, _04481_);
  nor (_26619_, _26618_, _26616_);
  or (_26620_, _26619_, _26595_);
  and (_26621_, _26620_, _03589_);
  nor (_26622_, _13332_, _10458_);
  nor (_26623_, _26622_, _26585_);
  nor (_26624_, _26623_, _03589_);
  or (_26625_, _26624_, _08828_);
  or (_26627_, _26625_, _26621_);
  and (_26628_, _13347_, _05221_);
  or (_26629_, _26585_, _07766_);
  or (_26630_, _26629_, _26628_);
  and (_26631_, _13339_, _05221_);
  nor (_26632_, _26631_, _26585_);
  and (_26633_, _26632_, _03601_);
  nor (_26634_, _26633_, _03780_);
  and (_26635_, _26634_, _26630_);
  and (_26636_, _26635_, _26627_);
  nor (_26637_, _26636_, _26591_);
  nor (_26638_, _26637_, _03622_);
  nor (_26639_, _26585_, _05412_);
  not (_26640_, _26639_);
  nor (_26641_, _26632_, _07777_);
  and (_26642_, _26641_, _26640_);
  nor (_26643_, _26642_, _26638_);
  nor (_26644_, _26643_, _03790_);
  nor (_26645_, _26597_, _06828_);
  and (_26646_, _26645_, _26640_);
  nor (_26649_, _26646_, _03624_);
  not (_26650_, _26649_);
  nor (_26651_, _26650_, _26644_);
  nor (_26652_, _13346_, _10458_);
  or (_26653_, _26585_, _07795_);
  nor (_26654_, _26653_, _26652_);
  or (_26655_, _26654_, _03785_);
  nor (_26656_, _26655_, _26651_);
  nor (_26657_, _26656_, _26588_);
  nor (_26658_, _26657_, _03815_);
  nor (_26660_, _26605_, _04246_);
  or (_26661_, _26660_, _03447_);
  nor (_26662_, _26661_, _26658_);
  and (_26663_, _13402_, _05221_);
  or (_26664_, _26585_, _03514_);
  nor (_26665_, _26664_, _26663_);
  nor (_26666_, _26665_, _26662_);
  or (_26667_, _26666_, _43004_);
  or (_26668_, _43000_, \oc8051_golden_model_1.SBUF [6]);
  and (_26669_, _26668_, _41806_);
  and (_43595_, _26669_, _26667_);
  not (_26671_, \oc8051_golden_model_1.SCON [0]);
  nor (_26672_, _05275_, _26671_);
  and (_26673_, _12128_, _05275_);
  nor (_26674_, _26673_, _26672_);
  nor (_26675_, _26674_, _07778_);
  and (_26676_, _05275_, _06274_);
  nor (_26677_, _26676_, _26672_);
  and (_26678_, _26677_, _03601_);
  and (_26679_, _05275_, _04620_);
  nor (_26681_, _26679_, _26672_);
  and (_26682_, _26681_, _07390_);
  and (_26683_, _05275_, \oc8051_golden_model_1.ACC [0]);
  nor (_26684_, _26683_, _26672_);
  nor (_26685_, _26684_, _09029_);
  nor (_26686_, _04409_, _26671_);
  or (_26687_, _26686_, _26685_);
  and (_26688_, _26687_, _04081_);
  nor (_26689_, _05666_, _10539_);
  nor (_26690_, _26689_, _26672_);
  nor (_26692_, _26690_, _04081_);
  or (_26693_, _26692_, _26688_);
  and (_26694_, _26693_, _04055_);
  nor (_26695_, _05922_, _26671_);
  and (_26696_, _12021_, _05922_);
  nor (_26697_, _26696_, _26695_);
  nor (_26698_, _26697_, _04055_);
  nor (_26699_, _26698_, _26694_);
  nor (_26700_, _26699_, _03723_);
  nor (_26701_, _26681_, _03996_);
  or (_26703_, _26701_, _26700_);
  and (_26704_, _26703_, _03737_);
  nor (_26705_, _26684_, _03737_);
  or (_26706_, _26705_, _26704_);
  and (_26707_, _26706_, _03736_);
  and (_26708_, _26672_, _03714_);
  or (_26709_, _26708_, _26707_);
  and (_26710_, _26709_, _06840_);
  nor (_26711_, _26690_, _06840_);
  or (_26712_, _26711_, _26710_);
  and (_26714_, _26712_, _03710_);
  nor (_26715_, _12052_, _10576_);
  nor (_26716_, _26715_, _26695_);
  nor (_26717_, _26716_, _03710_);
  or (_26718_, _26717_, _07390_);
  nor (_26719_, _26718_, _26714_);
  nor (_26720_, _26719_, _26682_);
  nor (_26721_, _26720_, _04481_);
  and (_26722_, _06546_, _05275_);
  nor (_26723_, _26672_, _07400_);
  not (_26725_, _26723_);
  nor (_26726_, _26725_, _26722_);
  or (_26727_, _26726_, _03222_);
  nor (_26728_, _26727_, _26721_);
  nor (_26729_, _12109_, _10539_);
  nor (_26730_, _26729_, _26672_);
  nor (_26731_, _26730_, _03589_);
  or (_26732_, _26731_, _03601_);
  nor (_26733_, _26732_, _26728_);
  nor (_26734_, _26733_, _26678_);
  or (_26736_, _26734_, _03600_);
  and (_26737_, _12124_, _05275_);
  or (_26738_, _26737_, _26672_);
  or (_26739_, _26738_, _07766_);
  and (_26740_, _26739_, _07778_);
  and (_26741_, _26740_, _26736_);
  nor (_26742_, _26741_, _26675_);
  nor (_26743_, _26742_, _03622_);
  or (_26744_, _26677_, _07777_);
  nor (_26745_, _26744_, _26689_);
  nor (_26747_, _26745_, _26743_);
  nor (_26748_, _26747_, _03790_);
  and (_26749_, _12005_, _05275_);
  or (_26750_, _26749_, _26672_);
  and (_26751_, _26750_, _03790_);
  or (_26752_, _26751_, _26748_);
  and (_26753_, _26752_, _07795_);
  nor (_26754_, _12122_, _10539_);
  nor (_26755_, _26754_, _26672_);
  nor (_26756_, _26755_, _07795_);
  or (_26758_, _26756_, _26753_);
  and (_26759_, _26758_, _07793_);
  nor (_26760_, _12003_, _10539_);
  nor (_26761_, _26760_, _26672_);
  nor (_26762_, _26761_, _07793_);
  or (_26763_, _26762_, _26759_);
  and (_26764_, _26763_, _04246_);
  nor (_26765_, _26690_, _04246_);
  or (_26766_, _26765_, _26764_);
  and (_26767_, _26766_, _03823_);
  and (_26769_, _26672_, _03453_);
  nor (_26770_, _26769_, _03447_);
  not (_26771_, _26770_);
  nor (_26772_, _26771_, _26767_);
  and (_26773_, _26690_, _03447_);
  or (_26774_, _26773_, _26772_);
  nand (_26775_, _26774_, _43000_);
  or (_26776_, _43000_, \oc8051_golden_model_1.SCON [0]);
  and (_26777_, _26776_, _41806_);
  and (_43596_, _26777_, _26775_);
  not (_26779_, \oc8051_golden_model_1.SCON [1]);
  nor (_26780_, _05275_, _26779_);
  and (_26781_, _06501_, _05275_);
  or (_26782_, _26781_, _26780_);
  and (_26783_, _26782_, _04481_);
  nor (_26784_, _05275_, \oc8051_golden_model_1.SCON [1]);
  and (_26785_, _05275_, _03274_);
  nor (_26786_, _26785_, _26784_);
  and (_26787_, _26786_, _04409_);
  nor (_26788_, _04409_, _26779_);
  or (_26790_, _26788_, _26787_);
  and (_26791_, _26790_, _04081_);
  and (_26792_, _12213_, _05275_);
  nor (_26793_, _26792_, _26784_);
  and (_26794_, _26793_, _03610_);
  or (_26795_, _26794_, _26791_);
  and (_26796_, _26795_, _04055_);
  and (_26797_, _12224_, _05922_);
  nor (_26798_, _05922_, _26779_);
  or (_26799_, _26798_, _03723_);
  or (_26801_, _26799_, _26797_);
  and (_26802_, _26801_, _14265_);
  nor (_26803_, _26802_, _26796_);
  and (_26804_, _05275_, _06764_);
  nor (_26805_, _26804_, _26780_);
  and (_26806_, _26805_, _03723_);
  nor (_26807_, _26806_, _26803_);
  and (_26808_, _26807_, _03737_);
  and (_26809_, _26786_, _03729_);
  or (_26810_, _26809_, _26808_);
  and (_26812_, _26810_, _03736_);
  and (_26813_, _12211_, _05922_);
  nor (_26814_, _26813_, _26798_);
  nor (_26815_, _26814_, _03736_);
  or (_26816_, _26815_, _26812_);
  and (_26817_, _26816_, _06840_);
  and (_26818_, _26797_, _12239_);
  or (_26819_, _26818_, _26798_);
  and (_26820_, _26819_, _03719_);
  or (_26821_, _26820_, _26817_);
  and (_26823_, _26821_, _03710_);
  nor (_26824_, _12256_, _10576_);
  nor (_26825_, _26798_, _26824_);
  nor (_26826_, _26825_, _03710_);
  or (_26827_, _26826_, _07390_);
  nor (_26828_, _26827_, _26823_);
  and (_26829_, _26805_, _07390_);
  or (_26830_, _26829_, _04481_);
  nor (_26831_, _26830_, _26828_);
  or (_26832_, _26831_, _26783_);
  and (_26834_, _26832_, _03589_);
  nor (_26835_, _12313_, _10539_);
  nor (_26836_, _26835_, _26780_);
  nor (_26837_, _26836_, _03589_);
  nor (_26838_, _26837_, _26834_);
  nor (_26839_, _26838_, _08828_);
  not (_26840_, _26784_);
  nor (_26841_, _12327_, _10539_);
  nor (_26842_, _26841_, _07766_);
  and (_26843_, _05275_, _04303_);
  nor (_26845_, _26843_, _05886_);
  or (_26846_, _26845_, _26842_);
  and (_26847_, _26846_, _26840_);
  nor (_26848_, _26847_, _26839_);
  nor (_26849_, _26848_, _03780_);
  nor (_26850_, _12333_, _10539_);
  nor (_26851_, _26850_, _07778_);
  and (_26852_, _26851_, _26840_);
  nor (_26853_, _26852_, _26849_);
  nor (_26854_, _26853_, _03622_);
  nor (_26856_, _12207_, _10539_);
  nor (_26857_, _26856_, _07777_);
  and (_26858_, _26857_, _26840_);
  nor (_26859_, _26858_, _26854_);
  nor (_26860_, _26859_, _03790_);
  nor (_26861_, _26780_, _05618_);
  nor (_26862_, _26861_, _06828_);
  and (_26863_, _26862_, _26786_);
  nor (_26864_, _26863_, _26860_);
  or (_26865_, _26864_, _18499_);
  and (_26867_, _26785_, _05617_);
  nor (_26868_, _26867_, _07793_);
  and (_26869_, _26868_, _26840_);
  nor (_26870_, _26869_, _03815_);
  and (_26871_, _26843_, _05617_);
  or (_26872_, _26784_, _07795_);
  or (_26873_, _26872_, _26871_);
  and (_26874_, _26873_, _26870_);
  and (_26875_, _26874_, _26865_);
  nor (_26876_, _26793_, _04246_);
  or (_26878_, _26876_, _03453_);
  nor (_26879_, _26878_, _26875_);
  nor (_26880_, _26814_, _03823_);
  or (_26881_, _26880_, _03447_);
  nor (_26882_, _26881_, _26879_);
  nor (_26883_, _26792_, _26780_);
  and (_26884_, _26883_, _03447_);
  nor (_26885_, _26884_, _26882_);
  or (_26886_, _26885_, _43004_);
  or (_26887_, _43000_, \oc8051_golden_model_1.SCON [1]);
  and (_26889_, _26887_, _41806_);
  and (_43599_, _26889_, _26886_);
  not (_26890_, \oc8051_golden_model_1.SCON [2]);
  nor (_26891_, _05275_, _26890_);
  and (_26892_, _05275_, _06332_);
  nor (_26893_, _26892_, _26891_);
  and (_26894_, _26893_, _03601_);
  nor (_26895_, _10539_, _04875_);
  nor (_26896_, _26895_, _26891_);
  and (_26897_, _26896_, _07390_);
  nor (_26899_, _26896_, _03996_);
  nor (_26900_, _05922_, _26890_);
  and (_26901_, _12411_, _05922_);
  nor (_26902_, _26901_, _26900_);
  and (_26903_, _26902_, _03715_);
  nor (_26904_, _12416_, _10539_);
  nor (_26905_, _26904_, _26891_);
  nor (_26906_, _26905_, _04081_);
  nor (_26907_, _04409_, _26890_);
  and (_26908_, _05275_, \oc8051_golden_model_1.ACC [2]);
  nor (_26910_, _26908_, _26891_);
  nor (_26911_, _26910_, _09029_);
  nor (_26912_, _26911_, _26907_);
  nor (_26913_, _26912_, _03610_);
  or (_26914_, _26913_, _03715_);
  nor (_26915_, _26914_, _26906_);
  nor (_26916_, _26915_, _26903_);
  and (_26917_, _26916_, _03996_);
  or (_26918_, _26917_, _26899_);
  and (_26919_, _26918_, _03737_);
  nor (_26921_, _26910_, _03737_);
  or (_26922_, _26921_, _26919_);
  and (_26923_, _26922_, _03736_);
  and (_26924_, _12409_, _05922_);
  nor (_26925_, _26924_, _26900_);
  nor (_26926_, _26925_, _03736_);
  or (_26927_, _26926_, _26923_);
  and (_26928_, _26927_, _06840_);
  nor (_26929_, _26900_, _12443_);
  nor (_26930_, _26929_, _26902_);
  and (_26931_, _26930_, _03719_);
  or (_26932_, _26931_, _26928_);
  and (_26933_, _26932_, _03710_);
  nor (_26934_, _12461_, _10576_);
  nor (_26935_, _26934_, _26900_);
  nor (_26936_, _26935_, _03710_);
  nor (_26937_, _26936_, _07390_);
  not (_26938_, _26937_);
  nor (_26939_, _26938_, _26933_);
  nor (_26940_, _26939_, _26897_);
  nor (_26943_, _26940_, _04481_);
  and (_26944_, _06637_, _05275_);
  nor (_26945_, _26891_, _07400_);
  not (_26946_, _26945_);
  nor (_26947_, _26946_, _26944_);
  or (_26948_, _26947_, _03222_);
  nor (_26949_, _26948_, _26943_);
  nor (_26950_, _12519_, _10539_);
  nor (_26951_, _26891_, _26950_);
  nor (_26952_, _26951_, _03589_);
  or (_26954_, _26952_, _03601_);
  nor (_26955_, _26954_, _26949_);
  nor (_26956_, _26955_, _26894_);
  or (_26957_, _26956_, _03600_);
  and (_26958_, _12533_, _05275_);
  or (_26959_, _26958_, _26891_);
  or (_26960_, _26959_, _07766_);
  and (_26961_, _26960_, _07778_);
  and (_26962_, _26961_, _26957_);
  and (_26963_, _12539_, _05275_);
  nor (_26965_, _26963_, _26891_);
  nor (_26966_, _26965_, _07778_);
  nor (_26967_, _26966_, _26962_);
  nor (_26968_, _26967_, _03622_);
  nor (_26969_, _26891_, _05718_);
  not (_26970_, _26969_);
  nor (_26971_, _26893_, _07777_);
  and (_26972_, _26971_, _26970_);
  nor (_26973_, _26972_, _26968_);
  nor (_26974_, _26973_, _03790_);
  nor (_26976_, _26910_, _06828_);
  and (_26977_, _26976_, _26970_);
  or (_26978_, _26977_, _26974_);
  and (_26979_, _26978_, _07795_);
  nor (_26980_, _12532_, _10539_);
  nor (_26981_, _26980_, _26891_);
  nor (_26982_, _26981_, _07795_);
  or (_26983_, _26982_, _26979_);
  and (_26984_, _26983_, _07793_);
  nor (_26985_, _12538_, _10539_);
  nor (_26987_, _26985_, _26891_);
  nor (_26988_, _26987_, _07793_);
  or (_26989_, _26988_, _26984_);
  and (_26990_, _26989_, _04246_);
  nor (_26991_, _26905_, _04246_);
  or (_26992_, _26991_, _26990_);
  and (_26993_, _26992_, _03823_);
  nor (_26994_, _26925_, _03823_);
  or (_26995_, _26994_, _26993_);
  and (_26996_, _26995_, _03514_);
  and (_26998_, _12592_, _05275_);
  nor (_26999_, _26998_, _26891_);
  nor (_27000_, _26999_, _03514_);
  or (_27001_, _27000_, _26996_);
  or (_27002_, _27001_, _43004_);
  or (_27003_, _43000_, \oc8051_golden_model_1.SCON [2]);
  and (_27004_, _27003_, _41806_);
  and (_43600_, _27004_, _27002_);
  not (_27005_, \oc8051_golden_model_1.SCON [3]);
  nor (_27006_, _05275_, _27005_);
  and (_27008_, _05275_, _06276_);
  nor (_27009_, _27008_, _27006_);
  and (_27010_, _27009_, _03601_);
  nor (_27011_, _10539_, _05005_);
  nor (_27012_, _27011_, _27006_);
  and (_27013_, _27012_, _07390_);
  and (_27014_, _05275_, \oc8051_golden_model_1.ACC [3]);
  nor (_27015_, _27014_, _27006_);
  nor (_27016_, _27015_, _09029_);
  nor (_27017_, _04409_, _27005_);
  or (_27019_, _27017_, _27016_);
  and (_27020_, _27019_, _04081_);
  nor (_27021_, _12627_, _10539_);
  nor (_27022_, _27021_, _27006_);
  nor (_27023_, _27022_, _04081_);
  or (_27024_, _27023_, _27020_);
  and (_27025_, _27024_, _04055_);
  nor (_27026_, _05922_, _27005_);
  and (_27027_, _12631_, _05922_);
  nor (_27028_, _27027_, _27026_);
  nor (_27030_, _27028_, _04055_);
  or (_27031_, _27030_, _03723_);
  or (_27032_, _27031_, _27025_);
  nand (_27033_, _27012_, _03723_);
  and (_27034_, _27033_, _27032_);
  and (_27035_, _27034_, _03737_);
  nor (_27036_, _27015_, _03737_);
  or (_27037_, _27036_, _27035_);
  and (_27038_, _27037_, _03736_);
  and (_27039_, _12641_, _05922_);
  nor (_27040_, _27039_, _27026_);
  nor (_27041_, _27040_, _03736_);
  or (_27042_, _27041_, _03719_);
  or (_27043_, _27042_, _27038_);
  nor (_27044_, _27026_, _12648_);
  nor (_27045_, _27044_, _27028_);
  or (_27046_, _27045_, _06840_);
  and (_27047_, _27046_, _03710_);
  and (_27048_, _27047_, _27043_);
  nor (_27049_, _12612_, _10576_);
  nor (_27052_, _27049_, _27026_);
  nor (_27053_, _27052_, _03710_);
  nor (_27054_, _27053_, _07390_);
  not (_27055_, _27054_);
  nor (_27056_, _27055_, _27048_);
  nor (_27057_, _27056_, _27013_);
  nor (_27058_, _27057_, _04481_);
  and (_27059_, _06592_, _05275_);
  nor (_27060_, _27006_, _07400_);
  not (_27061_, _27060_);
  nor (_27063_, _27061_, _27059_);
  or (_27064_, _27063_, _03222_);
  nor (_27065_, _27064_, _27058_);
  nor (_27066_, _12718_, _10539_);
  nor (_27067_, _27006_, _27066_);
  nor (_27068_, _27067_, _03589_);
  or (_27069_, _27068_, _03601_);
  nor (_27070_, _27069_, _27065_);
  nor (_27071_, _27070_, _27010_);
  or (_27072_, _27071_, _03600_);
  and (_27074_, _12733_, _05275_);
  or (_27075_, _27074_, _27006_);
  or (_27076_, _27075_, _07766_);
  and (_27077_, _27076_, _07778_);
  and (_27078_, _27077_, _27072_);
  and (_27079_, _12739_, _05275_);
  nor (_27080_, _27079_, _27006_);
  nor (_27081_, _27080_, _07778_);
  nor (_27082_, _27081_, _27078_);
  nor (_27083_, _27082_, _03622_);
  nor (_27085_, _27006_, _05567_);
  not (_27086_, _27085_);
  nor (_27087_, _27009_, _07777_);
  and (_27088_, _27087_, _27086_);
  nor (_27089_, _27088_, _27083_);
  nor (_27090_, _27089_, _03790_);
  nor (_27091_, _27015_, _06828_);
  and (_27092_, _27091_, _27086_);
  nor (_27093_, _27092_, _03624_);
  not (_27094_, _27093_);
  nor (_27096_, _27094_, _27090_);
  nor (_27097_, _12732_, _10539_);
  or (_27098_, _27006_, _07795_);
  nor (_27099_, _27098_, _27097_);
  or (_27100_, _27099_, _03785_);
  nor (_27101_, _27100_, _27096_);
  nor (_27102_, _12738_, _10539_);
  nor (_27103_, _27102_, _27006_);
  nor (_27104_, _27103_, _07793_);
  or (_27105_, _27104_, _27101_);
  and (_27107_, _27105_, _04246_);
  nor (_27108_, _27022_, _04246_);
  or (_27109_, _27108_, _27107_);
  and (_27110_, _27109_, _03823_);
  nor (_27111_, _27040_, _03823_);
  or (_27112_, _27111_, _27110_);
  and (_27113_, _27112_, _03514_);
  and (_27114_, _12794_, _05275_);
  nor (_27115_, _27114_, _27006_);
  nor (_27116_, _27115_, _03514_);
  or (_27118_, _27116_, _27113_);
  or (_27119_, _27118_, _43004_);
  or (_27120_, _43000_, \oc8051_golden_model_1.SCON [3]);
  and (_27121_, _27120_, _41806_);
  and (_43601_, _27121_, _27119_);
  not (_27122_, \oc8051_golden_model_1.SCON [4]);
  nor (_27123_, _05275_, _27122_);
  nor (_27124_, _05777_, _10539_);
  nor (_27125_, _27124_, _27123_);
  and (_27126_, _27125_, _07390_);
  nor (_27128_, _05922_, _27122_);
  and (_27129_, _12827_, _05922_);
  nor (_27130_, _27129_, _27128_);
  nor (_27131_, _27130_, _03736_);
  and (_27132_, _05275_, \oc8051_golden_model_1.ACC [4]);
  nor (_27133_, _27132_, _27123_);
  nor (_27134_, _27133_, _09029_);
  nor (_27135_, _04409_, _27122_);
  or (_27136_, _27135_, _27134_);
  and (_27137_, _27136_, _04081_);
  nor (_27139_, _12841_, _10539_);
  nor (_27140_, _27139_, _27123_);
  nor (_27141_, _27140_, _04081_);
  or (_27142_, _27141_, _27137_);
  and (_27143_, _27142_, _04055_);
  and (_27144_, _12845_, _05922_);
  nor (_27145_, _27144_, _27128_);
  nor (_27146_, _27145_, _04055_);
  or (_27147_, _27146_, _03723_);
  or (_27148_, _27147_, _27143_);
  nand (_27150_, _27125_, _03723_);
  and (_27151_, _27150_, _27148_);
  and (_27152_, _27151_, _03737_);
  nor (_27153_, _27133_, _03737_);
  or (_27154_, _27153_, _27152_);
  and (_27155_, _27154_, _03736_);
  nor (_27156_, _27155_, _27131_);
  nor (_27157_, _27156_, _03719_);
  nor (_27158_, _27128_, _12860_);
  or (_27159_, _27145_, _06840_);
  nor (_27161_, _27159_, _27158_);
  nor (_27162_, _27161_, _27157_);
  nor (_27163_, _27162_, _03505_);
  nor (_27164_, _12825_, _10576_);
  nor (_27165_, _27164_, _27128_);
  nor (_27166_, _27165_, _03710_);
  nor (_27167_, _27166_, _07390_);
  not (_27168_, _27167_);
  nor (_27169_, _27168_, _27163_);
  nor (_27170_, _27169_, _27126_);
  nor (_27172_, _27170_, _04481_);
  and (_27173_, _06730_, _05275_);
  nor (_27174_, _27123_, _07400_);
  not (_27175_, _27174_);
  nor (_27176_, _27175_, _27173_);
  nor (_27177_, _27176_, _03222_);
  not (_27178_, _27177_);
  nor (_27179_, _27178_, _27172_);
  nor (_27180_, _12933_, _10539_);
  nor (_27181_, _27180_, _27123_);
  nor (_27183_, _27181_, _03589_);
  or (_27184_, _27183_, _08828_);
  or (_27185_, _27184_, _27179_);
  and (_27186_, _12821_, _05275_);
  or (_27187_, _27123_, _07766_);
  or (_27188_, _27187_, _27186_);
  and (_27189_, _06298_, _05275_);
  nor (_27190_, _27189_, _27123_);
  and (_27191_, _27190_, _03601_);
  nor (_27192_, _27191_, _03780_);
  and (_27194_, _27192_, _27188_);
  and (_27195_, _27194_, _27185_);
  and (_27196_, _12817_, _05275_);
  nor (_27197_, _27196_, _27123_);
  nor (_27198_, _27197_, _07778_);
  nor (_27199_, _27198_, _27195_);
  nor (_27200_, _27199_, _03622_);
  nor (_27201_, _27123_, _05825_);
  not (_27202_, _27201_);
  nor (_27203_, _27190_, _07777_);
  and (_27205_, _27203_, _27202_);
  nor (_27206_, _27205_, _27200_);
  nor (_27207_, _27206_, _03790_);
  nor (_27208_, _27133_, _06828_);
  and (_27209_, _27208_, _27202_);
  nor (_27210_, _27209_, _03624_);
  not (_27211_, _27210_);
  nor (_27212_, _27211_, _27207_);
  nor (_27213_, _12819_, _10539_);
  or (_27214_, _27123_, _07795_);
  nor (_27216_, _27214_, _27213_);
  or (_27217_, _27216_, _03785_);
  nor (_27218_, _27217_, _27212_);
  nor (_27219_, _12816_, _10539_);
  nor (_27220_, _27219_, _27123_);
  nor (_27221_, _27220_, _07793_);
  or (_27222_, _27221_, _27218_);
  and (_27223_, _27222_, _04246_);
  nor (_27224_, _27140_, _04246_);
  or (_27225_, _27224_, _27223_);
  and (_27227_, _27225_, _03823_);
  nor (_27228_, _27130_, _03823_);
  or (_27229_, _27228_, _27227_);
  and (_27230_, _27229_, _03514_);
  and (_27231_, _13003_, _05275_);
  nor (_27232_, _27231_, _27123_);
  nor (_27233_, _27232_, _03514_);
  or (_27234_, _27233_, _27230_);
  or (_27235_, _27234_, _43004_);
  or (_27236_, _43000_, \oc8051_golden_model_1.SCON [4]);
  and (_27238_, _27236_, _41806_);
  and (_43602_, _27238_, _27235_);
  not (_27239_, \oc8051_golden_model_1.SCON [5]);
  nor (_27240_, _05275_, _27239_);
  and (_27241_, _06684_, _05275_);
  or (_27242_, _27241_, _27240_);
  and (_27243_, _27242_, _04481_);
  and (_27244_, _05275_, \oc8051_golden_model_1.ACC [5]);
  nor (_27245_, _27244_, _27240_);
  nor (_27246_, _27245_, _09029_);
  nor (_27248_, _04409_, _27239_);
  or (_27249_, _27248_, _27246_);
  and (_27250_, _27249_, _04081_);
  nor (_27251_, _13014_, _10539_);
  nor (_27252_, _27251_, _27240_);
  nor (_27253_, _27252_, _04081_);
  or (_27254_, _27253_, _27250_);
  and (_27255_, _27254_, _04055_);
  nor (_27256_, _05922_, _27239_);
  and (_27257_, _13037_, _05922_);
  nor (_27258_, _27257_, _27256_);
  nor (_27259_, _27258_, _04055_);
  or (_27260_, _27259_, _03723_);
  or (_27261_, _27260_, _27255_);
  nor (_27262_, _05469_, _10539_);
  nor (_27263_, _27262_, _27240_);
  nand (_27264_, _27263_, _03723_);
  and (_27265_, _27264_, _27261_);
  and (_27266_, _27265_, _03737_);
  nor (_27267_, _27245_, _03737_);
  or (_27270_, _27267_, _27266_);
  and (_27271_, _27270_, _03736_);
  and (_27272_, _13047_, _05922_);
  nor (_27273_, _27272_, _27256_);
  nor (_27274_, _27273_, _03736_);
  or (_27275_, _27274_, _27271_);
  and (_27276_, _27275_, _06840_);
  nor (_27277_, _27256_, _13054_);
  nor (_27278_, _27277_, _27258_);
  and (_27279_, _27278_, _03719_);
  or (_27281_, _27279_, _27276_);
  and (_27282_, _27281_, _03710_);
  nor (_27283_, _13020_, _10576_);
  nor (_27284_, _27283_, _27256_);
  nor (_27285_, _27284_, _03710_);
  nor (_27286_, _27285_, _07390_);
  not (_27287_, _27286_);
  nor (_27288_, _27287_, _27282_);
  and (_27289_, _27263_, _07390_);
  or (_27290_, _27289_, _04481_);
  nor (_27292_, _27290_, _27288_);
  or (_27293_, _27292_, _27243_);
  and (_27294_, _27293_, _03589_);
  nor (_27295_, _13127_, _10539_);
  nor (_27296_, _27295_, _27240_);
  nor (_27297_, _27296_, _03589_);
  or (_27298_, _27297_, _08828_);
  or (_27299_, _27298_, _27294_);
  and (_27300_, _13141_, _05275_);
  or (_27301_, _27240_, _07766_);
  or (_27303_, _27301_, _27300_);
  and (_27304_, _06306_, _05275_);
  nor (_27305_, _27304_, _27240_);
  and (_27306_, _27305_, _03601_);
  nor (_27307_, _27306_, _03780_);
  and (_27308_, _27307_, _27303_);
  and (_27309_, _27308_, _27299_);
  and (_27310_, _13147_, _05275_);
  nor (_27311_, _27310_, _27240_);
  nor (_27312_, _27311_, _07778_);
  nor (_27314_, _27312_, _27309_);
  nor (_27315_, _27314_, _03622_);
  nor (_27316_, _27240_, _05518_);
  not (_27317_, _27316_);
  nor (_27318_, _27305_, _07777_);
  and (_27319_, _27318_, _27317_);
  nor (_27320_, _27319_, _27315_);
  nor (_27321_, _27320_, _03790_);
  nor (_27322_, _27245_, _06828_);
  and (_27323_, _27322_, _27317_);
  nor (_27325_, _27323_, _03624_);
  not (_27326_, _27325_);
  nor (_27327_, _27326_, _27321_);
  nor (_27328_, _13140_, _10539_);
  or (_27329_, _27240_, _07795_);
  nor (_27330_, _27329_, _27328_);
  or (_27331_, _27330_, _03785_);
  nor (_27332_, _27331_, _27327_);
  nor (_27333_, _13146_, _10539_);
  nor (_27334_, _27333_, _27240_);
  nor (_27336_, _27334_, _07793_);
  or (_27337_, _27336_, _27332_);
  and (_27338_, _27337_, _04246_);
  nor (_27339_, _27252_, _04246_);
  or (_27340_, _27339_, _27338_);
  and (_27341_, _27340_, _03823_);
  nor (_27342_, _27273_, _03823_);
  or (_27343_, _27342_, _27341_);
  and (_27344_, _27343_, _03514_);
  and (_27345_, _13199_, _05275_);
  nor (_27347_, _27345_, _27240_);
  nor (_27348_, _27347_, _03514_);
  or (_27349_, _27348_, _27344_);
  or (_27350_, _27349_, _43004_);
  or (_27351_, _43000_, \oc8051_golden_model_1.SCON [5]);
  and (_27352_, _27351_, _41806_);
  and (_43603_, _27352_, _27350_);
  not (_27353_, \oc8051_golden_model_1.SCON [6]);
  nor (_27354_, _05275_, _27353_);
  and (_27355_, _06455_, _05275_);
  or (_27357_, _27355_, _27354_);
  and (_27358_, _27357_, _04481_);
  and (_27359_, _05275_, \oc8051_golden_model_1.ACC [6]);
  nor (_27360_, _27359_, _27354_);
  nor (_27361_, _27360_, _09029_);
  nor (_27362_, _04409_, _27353_);
  or (_27363_, _27362_, _27361_);
  and (_27364_, _27363_, _04081_);
  nor (_27365_, _13242_, _10539_);
  nor (_27366_, _27365_, _27354_);
  nor (_27368_, _27366_, _04081_);
  or (_27369_, _27368_, _27364_);
  and (_27370_, _27369_, _04055_);
  nor (_27371_, _05922_, _27353_);
  and (_27372_, _13229_, _05922_);
  nor (_27373_, _27372_, _27371_);
  nor (_27374_, _27373_, _04055_);
  or (_27375_, _27374_, _03723_);
  or (_27376_, _27375_, _27370_);
  nor (_27377_, _05363_, _10539_);
  nor (_27379_, _27377_, _27354_);
  nand (_27380_, _27379_, _03723_);
  and (_27381_, _27380_, _27376_);
  and (_27382_, _27381_, _03737_);
  nor (_27383_, _27360_, _03737_);
  or (_27384_, _27383_, _27382_);
  and (_27385_, _27384_, _03736_);
  and (_27386_, _13253_, _05922_);
  nor (_27387_, _27386_, _27371_);
  nor (_27388_, _27387_, _03736_);
  or (_27390_, _27388_, _03719_);
  or (_27391_, _27390_, _27385_);
  nor (_27392_, _27371_, _13260_);
  nor (_27393_, _27392_, _27373_);
  or (_27394_, _27393_, _06840_);
  and (_27395_, _27394_, _03710_);
  and (_27396_, _27395_, _27391_);
  nor (_27397_, _13226_, _10576_);
  nor (_27398_, _27397_, _27371_);
  nor (_27399_, _27398_, _03710_);
  nor (_27401_, _27399_, _07390_);
  not (_27402_, _27401_);
  nor (_27403_, _27402_, _27396_);
  and (_27404_, _27379_, _07390_);
  or (_27405_, _27404_, _04481_);
  nor (_27406_, _27405_, _27403_);
  or (_27407_, _27406_, _27358_);
  and (_27408_, _27407_, _03589_);
  nor (_27409_, _13332_, _10539_);
  nor (_27410_, _27409_, _27354_);
  nor (_27412_, _27410_, _03589_);
  or (_27413_, _27412_, _08828_);
  or (_27414_, _27413_, _27408_);
  and (_27415_, _13347_, _05275_);
  or (_27416_, _27354_, _07766_);
  or (_27417_, _27416_, _27415_);
  and (_27418_, _13339_, _05275_);
  nor (_27419_, _27418_, _27354_);
  and (_27420_, _27419_, _03601_);
  nor (_27421_, _27420_, _03780_);
  and (_27423_, _27421_, _27417_);
  and (_27424_, _27423_, _27414_);
  and (_27425_, _13353_, _05275_);
  nor (_27426_, _27425_, _27354_);
  nor (_27427_, _27426_, _07778_);
  nor (_27428_, _27427_, _27424_);
  nor (_27429_, _27428_, _03622_);
  nor (_27430_, _27354_, _05412_);
  not (_27431_, _27430_);
  nor (_27432_, _27419_, _07777_);
  and (_27434_, _27432_, _27431_);
  nor (_27435_, _27434_, _27429_);
  nor (_27436_, _27435_, _03790_);
  nor (_27437_, _27360_, _06828_);
  and (_27438_, _27437_, _27431_);
  nor (_27439_, _27438_, _03624_);
  not (_27440_, _27439_);
  nor (_27441_, _27440_, _27436_);
  nor (_27442_, _13346_, _10539_);
  or (_27443_, _27354_, _07795_);
  nor (_27445_, _27443_, _27442_);
  or (_27446_, _27445_, _03785_);
  nor (_27447_, _27446_, _27441_);
  nor (_27448_, _13352_, _10539_);
  nor (_27449_, _27448_, _27354_);
  nor (_27450_, _27449_, _07793_);
  or (_27451_, _27450_, _27447_);
  and (_27452_, _27451_, _04246_);
  nor (_27453_, _27366_, _04246_);
  or (_27454_, _27453_, _27452_);
  and (_27456_, _27454_, _03823_);
  nor (_27457_, _27387_, _03823_);
  or (_27458_, _27457_, _27456_);
  and (_27459_, _27458_, _03514_);
  and (_27460_, _13402_, _05275_);
  nor (_27461_, _27460_, _27354_);
  nor (_27462_, _27461_, _03514_);
  or (_27463_, _27462_, _27459_);
  or (_27464_, _27463_, _43004_);
  or (_27465_, _43000_, \oc8051_golden_model_1.SCON [6]);
  and (_27467_, _27465_, _41806_);
  and (_43604_, _27467_, _27464_);
  nor (_27468_, _05300_, _03498_);
  nor (_27469_, _05666_, _10706_);
  nor (_27470_, _27469_, _27468_);
  and (_27471_, _27470_, _17166_);
  and (_27472_, _05300_, \oc8051_golden_model_1.ACC [0]);
  nor (_27473_, _27472_, _27468_);
  nor (_27474_, _27473_, _09029_);
  nor (_27475_, _04409_, _03498_);
  or (_27477_, _27475_, _27474_);
  and (_27478_, _27477_, _04081_);
  nor (_27479_, _27470_, _04081_);
  or (_27480_, _27479_, _27478_);
  and (_27481_, _27480_, _03996_);
  nor (_27482_, _27481_, _04089_);
  and (_27483_, _27473_, _03729_);
  nor (_27484_, _27483_, _03508_);
  not (_27485_, _27484_);
  nor (_27486_, _27485_, _27482_);
  nor (_27488_, _07390_, _04657_);
  not (_27489_, _27488_);
  nor (_27490_, _27489_, _27486_);
  not (_27491_, _27468_);
  and (_27492_, _05300_, _04620_);
  nor (_27493_, _27492_, _06838_);
  and (_27494_, _27493_, _27491_);
  nor (_27495_, _27494_, _27490_);
  nor (_27496_, _27495_, _04481_);
  and (_27497_, _06546_, _05300_);
  nor (_27499_, _27468_, _07400_);
  not (_27500_, _27499_);
  nor (_27501_, _27500_, _27497_);
  nor (_27502_, _27501_, _27496_);
  nor (_27503_, _27502_, _03222_);
  nor (_27504_, _12109_, _10706_);
  or (_27505_, _27468_, _03589_);
  nor (_27506_, _27505_, _27504_);
  or (_27507_, _27506_, _03601_);
  nor (_27508_, _27507_, _27503_);
  and (_27510_, _05300_, _06274_);
  nor (_27511_, _27510_, _27468_);
  nand (_27512_, _27511_, _07766_);
  and (_27513_, _27512_, _08828_);
  nor (_27514_, _27513_, _27508_);
  and (_27515_, _12124_, _05300_);
  nor (_27516_, _27515_, _27468_);
  and (_27517_, _27516_, _03600_);
  nor (_27518_, _27517_, _27514_);
  nor (_27519_, _27518_, _03780_);
  and (_27520_, _12128_, _05300_);
  or (_27521_, _27468_, _07778_);
  nor (_27522_, _27521_, _27520_);
  or (_27523_, _27522_, _03622_);
  nor (_27524_, _27523_, _27519_);
  or (_27525_, _27511_, _07777_);
  nor (_27526_, _27525_, _27469_);
  nor (_27527_, _27526_, _27524_);
  nor (_27528_, _27527_, _03790_);
  and (_27529_, _12005_, _05300_);
  or (_27532_, _27529_, _27468_);
  and (_27533_, _27532_, _03790_);
  or (_27534_, _27533_, _27528_);
  and (_27535_, _27534_, _07795_);
  nor (_27536_, _12122_, _10706_);
  nor (_27537_, _27536_, _27468_);
  nor (_27538_, _27537_, _07795_);
  or (_27539_, _27538_, _27535_);
  and (_27540_, _27539_, _07793_);
  nor (_27541_, _12003_, _10706_);
  nor (_27543_, _27541_, _27468_);
  nor (_27544_, _27543_, _07793_);
  nor (_27545_, _27544_, _17166_);
  not (_27546_, _27545_);
  nor (_27547_, _27546_, _27540_);
  nor (_27548_, _27547_, _27471_);
  and (_27549_, _27548_, _43000_);
  nor (_27550_, \oc8051_golden_model_1.SP [0], rst);
  nor (_27551_, _27550_, _00000_);
  or (_43606_, _27551_, _27549_);
  nor (_27553_, _05300_, _03496_);
  and (_27554_, _12213_, _05300_);
  nor (_27555_, _27554_, _27553_);
  nor (_27556_, _27555_, _03514_);
  nor (_27557_, _10774_, _03496_);
  and (_27558_, _03178_, _03496_);
  nor (_27559_, _05300_, \oc8051_golden_model_1.SP [1]);
  and (_27560_, _05300_, _03274_);
  nor (_27561_, _27560_, _27559_);
  and (_27562_, _27561_, _04409_);
  nor (_27564_, _04409_, _03496_);
  or (_27565_, _27564_, _27562_);
  and (_27566_, _27565_, _04763_);
  and (_27567_, _03980_, _03496_);
  or (_27568_, _27567_, _27566_);
  and (_27569_, _27568_, _04081_);
  nor (_27570_, _27559_, _27554_);
  and (_27571_, _27570_, _03610_);
  or (_27572_, _27571_, _27569_);
  and (_27573_, _27572_, _03230_);
  nor (_27575_, _03230_, \oc8051_golden_model_1.SP [1]);
  or (_27576_, _27575_, _03723_);
  or (_27577_, _27576_, _27573_);
  nand (_27578_, _03501_, _03723_);
  and (_27579_, _27578_, _27577_);
  and (_27580_, _27579_, _03737_);
  and (_27581_, _27561_, _03729_);
  or (_27582_, _27581_, _27580_);
  and (_27583_, _27582_, _03510_);
  or (_27584_, _27583_, _10694_);
  nor (_27586_, _27584_, _03509_);
  nor (_27587_, _04767_, _03496_);
  or (_27588_, _27587_, _07390_);
  nor (_27589_, _27588_, _27586_);
  or (_27590_, _10706_, _06764_);
  nor (_27591_, _27559_, _06838_);
  and (_27592_, _27591_, _27590_);
  nor (_27593_, _27592_, _04481_);
  not (_27594_, _27593_);
  nor (_27595_, _27594_, _27589_);
  and (_27597_, _06501_, _05300_);
  nor (_27598_, _27553_, _07400_);
  not (_27599_, _27598_);
  nor (_27600_, _27599_, _27597_);
  nor (_27601_, _27600_, _03222_);
  not (_27602_, _27601_);
  nor (_27603_, _27602_, _27595_);
  nor (_27604_, _12313_, _10706_);
  or (_27605_, _27604_, _27553_);
  and (_27606_, _27605_, _03222_);
  nor (_27608_, _27606_, _27603_);
  nor (_27609_, _27608_, _03601_);
  and (_27610_, _05300_, _06282_);
  or (_27611_, _27610_, _27553_);
  and (_27612_, _27611_, _03601_);
  or (_27613_, _27612_, _27609_);
  and (_27614_, _27613_, _10736_);
  or (_27615_, _27614_, _27558_);
  and (_27616_, _27615_, _07766_);
  nor (_27617_, _12327_, _10706_);
  or (_27619_, _27617_, _07766_);
  nor (_27620_, _27619_, _27559_);
  nor (_27621_, _27620_, _27616_);
  nor (_27622_, _27621_, _03780_);
  nor (_27623_, _12333_, _10706_);
  or (_27624_, _27623_, _07778_);
  nor (_27625_, _27624_, _27559_);
  nor (_27626_, _27625_, _27622_);
  nor (_27627_, _27626_, _03622_);
  nor (_27628_, _12207_, _10706_);
  or (_27630_, _27628_, _07777_);
  nor (_27631_, _27630_, _27559_);
  nor (_27632_, _27631_, _27627_);
  nor (_27633_, _27632_, _10754_);
  and (_27634_, _03192_, _03496_);
  nor (_27635_, _27553_, _05618_);
  nor (_27636_, _27635_, _06828_);
  and (_27637_, _27636_, _27561_);
  nor (_27638_, _27637_, _27634_);
  not (_27639_, _27638_);
  nor (_27641_, _27639_, _27633_);
  or (_27642_, _27641_, _18499_);
  nor (_27643_, _12332_, _10706_);
  or (_27644_, _27643_, _27553_);
  and (_27645_, _27644_, _03785_);
  not (_27646_, _10774_);
  nor (_27647_, _12326_, _10706_);
  or (_27648_, _27647_, _27553_);
  and (_27649_, _27648_, _03624_);
  or (_27650_, _27649_, _27646_);
  nor (_27652_, _27650_, _27645_);
  and (_27653_, _27652_, _27642_);
  nor (_27654_, _27653_, _27557_);
  and (_27655_, _27654_, _03516_);
  and (_27656_, _03515_, _03496_);
  or (_27657_, _27656_, _27655_);
  and (_27658_, _27657_, _04246_);
  and (_27659_, _27570_, _03815_);
  nor (_27660_, _27659_, _05103_);
  not (_27661_, _27660_);
  nor (_27663_, _27661_, _27658_);
  nor (_27664_, _04540_, _03496_);
  nor (_27665_, _27664_, _03447_);
  not (_27666_, _27665_);
  nor (_27667_, _27666_, _27663_);
  nor (_27668_, _27667_, _27556_);
  nor (_27669_, _27668_, _43004_);
  nor (_27670_, \oc8051_golden_model_1.SP [1], rst);
  nor (_27671_, _27670_, _00000_);
  or (_43607_, _27671_, _27669_);
  and (_27673_, _05129_, _03188_);
  nor (_27674_, _05300_, _03995_);
  and (_27675_, _12539_, _05300_);
  nor (_27676_, _27675_, _27674_);
  nor (_27677_, _27676_, _07778_);
  and (_27678_, _12192_, _03178_);
  not (_27679_, _27674_);
  nor (_27680_, _10706_, _04875_);
  nor (_27681_, _27680_, _06838_);
  and (_27682_, _27681_, _27679_);
  nor (_27684_, _12416_, _10706_);
  nor (_27685_, _27684_, _27674_);
  nor (_27686_, _27685_, _04081_);
  nor (_27687_, _04409_, _03995_);
  and (_27688_, _05300_, \oc8051_golden_model_1.ACC [2]);
  nor (_27689_, _27688_, _27674_);
  nor (_27690_, _27689_, _09029_);
  nor (_27691_, _27690_, _27687_);
  nor (_27692_, _27691_, _03980_);
  and (_27693_, _05129_, _03980_);
  nor (_27695_, _27693_, _27692_);
  nor (_27696_, _27695_, _03610_);
  or (_27697_, _27696_, _04768_);
  nor (_27698_, _27697_, _27686_);
  nor (_27699_, _05129_, _03230_);
  or (_27700_, _27699_, _03723_);
  nor (_27701_, _27700_, _27698_);
  nor (_27702_, _05984_, _03996_);
  or (_27703_, _27702_, _27701_);
  and (_27704_, _27703_, _03737_);
  nor (_27706_, _27689_, _03737_);
  or (_27707_, _27706_, _27704_);
  and (_27708_, _27707_, _03510_);
  nor (_27709_, _27708_, _04811_);
  nor (_27710_, _27709_, _10694_);
  nor (_27711_, _12192_, _04767_);
  nor (_27712_, _27711_, _07390_);
  not (_27713_, _27712_);
  nor (_27714_, _27713_, _27710_);
  nor (_27715_, _27714_, _27682_);
  nor (_27717_, _27715_, _04481_);
  and (_27718_, _06637_, _05300_);
  nor (_27719_, _27674_, _07400_);
  not (_27720_, _27719_);
  nor (_27721_, _27720_, _27718_);
  or (_27722_, _27721_, _03222_);
  nor (_27723_, _27722_, _27717_);
  nor (_27724_, _12519_, _10706_);
  nor (_27725_, _27724_, _27674_);
  nor (_27726_, _27725_, _03589_);
  or (_27728_, _27726_, _03601_);
  or (_27729_, _27728_, _27723_);
  and (_27730_, _05300_, _06332_);
  nor (_27731_, _27730_, _27674_);
  nand (_27732_, _27731_, _03601_);
  and (_27733_, _27732_, _27729_);
  nor (_27734_, _27733_, _03178_);
  nor (_27735_, _27734_, _27678_);
  nor (_27736_, _27735_, _03600_);
  and (_27737_, _12533_, _05300_);
  or (_27739_, _27674_, _07766_);
  nor (_27740_, _27739_, _27737_);
  or (_27741_, _27740_, _03780_);
  nor (_27742_, _27741_, _27736_);
  nor (_27743_, _27742_, _27677_);
  nor (_27744_, _27743_, _03622_);
  and (_27745_, _27679_, _05717_);
  not (_27746_, _27745_);
  nor (_27747_, _27731_, _07777_);
  and (_27748_, _27747_, _27746_);
  nor (_27750_, _27748_, _27744_);
  nor (_27751_, _27750_, _10754_);
  nor (_27752_, _27689_, _06828_);
  and (_27753_, _27752_, _27746_);
  and (_27754_, _05129_, _03192_);
  nor (_27755_, _27754_, _27753_);
  and (_27756_, _27755_, _07795_);
  not (_27757_, _27756_);
  nor (_27758_, _27757_, _27751_);
  nor (_27759_, _12532_, _10706_);
  nor (_27761_, _27759_, _27674_);
  and (_27762_, _27761_, _03624_);
  nor (_27763_, _27762_, _27758_);
  nor (_27764_, _27763_, _03785_);
  nor (_27765_, _12538_, _10706_);
  or (_27766_, _27674_, _07793_);
  nor (_27767_, _27766_, _27765_);
  or (_27768_, _27767_, _03798_);
  nor (_27769_, _27768_, _27764_);
  and (_27770_, _12192_, _03798_);
  or (_27772_, _27770_, _27769_);
  and (_27773_, _27772_, _06399_);
  or (_27774_, _27773_, _27673_);
  and (_27775_, _27774_, _03516_);
  and (_27776_, _12192_, _03515_);
  or (_27777_, _27776_, _03815_);
  nor (_27778_, _27777_, _27775_);
  and (_27779_, _27685_, _03815_);
  or (_27780_, _27779_, _05103_);
  nor (_27781_, _27780_, _27778_);
  nor (_27783_, _12192_, _04540_);
  nor (_27784_, _27783_, _03447_);
  not (_27785_, _27784_);
  nor (_27786_, _27785_, _27781_);
  and (_27787_, _12592_, _05300_);
  nor (_27788_, _27787_, _27674_);
  and (_27789_, _27788_, _03447_);
  nor (_27790_, _27789_, _27786_);
  and (_27791_, _27790_, _43000_);
  nor (_27792_, \oc8051_golden_model_1.SP [2], rst);
  nor (_27794_, _27792_, _00000_);
  or (_43608_, _27794_, _27791_);
  nor (_27795_, _05133_, _04540_);
  and (_27796_, _05133_, _03188_);
  and (_27797_, _05133_, _03192_);
  nor (_27798_, _27797_, _03624_);
  nor (_27799_, _05300_, _03722_);
  and (_27800_, _12739_, _05300_);
  nor (_27801_, _27800_, _27799_);
  nor (_27802_, _27801_, _07778_);
  and (_27803_, _05132_, _03178_);
  nor (_27804_, _04409_, _03722_);
  and (_27805_, _05300_, \oc8051_golden_model_1.ACC [3]);
  nor (_27806_, _27805_, _27799_);
  nor (_27807_, _27806_, _09029_);
  or (_27808_, _27807_, _27804_);
  and (_27809_, _27808_, _04763_);
  and (_27810_, _05133_, _03980_);
  nor (_27811_, _27810_, _27809_);
  nor (_27812_, _27811_, _03610_);
  nor (_27815_, _12627_, _10706_);
  nor (_27816_, _27815_, _27799_);
  nor (_27817_, _27816_, _04081_);
  or (_27818_, _27817_, _27812_);
  and (_27819_, _27818_, _03230_);
  nor (_27820_, _05132_, _03230_);
  or (_27821_, _27820_, _03723_);
  or (_27822_, _27821_, _27819_);
  nand (_27823_, _05973_, _03723_);
  and (_27824_, _27823_, _27822_);
  and (_27826_, _27824_, _03737_);
  nor (_27827_, _27806_, _03737_);
  or (_27828_, _27827_, _27826_);
  and (_27829_, _27828_, _03510_);
  or (_27830_, _27829_, _10694_);
  nor (_27831_, _27830_, _05053_);
  nor (_27832_, _05133_, _04767_);
  or (_27833_, _27832_, _07390_);
  nor (_27834_, _27833_, _27831_);
  nor (_27835_, _10706_, _05005_);
  nor (_27837_, _27835_, _27799_);
  nor (_27838_, _27837_, _06838_);
  nor (_27839_, _27838_, _04481_);
  not (_27840_, _27839_);
  nor (_27841_, _27840_, _27834_);
  and (_27842_, _06592_, _05300_);
  nor (_27843_, _27799_, _07400_);
  not (_27844_, _27843_);
  nor (_27845_, _27844_, _27842_);
  or (_27846_, _27845_, _03222_);
  nor (_27848_, _27846_, _27841_);
  nor (_27849_, _12718_, _10706_);
  nor (_27850_, _27849_, _27799_);
  nor (_27851_, _27850_, _03589_);
  or (_27852_, _27851_, _03601_);
  or (_27853_, _27852_, _27848_);
  and (_27854_, _05300_, _06276_);
  nor (_27855_, _27854_, _27799_);
  nand (_27856_, _27855_, _03601_);
  and (_27857_, _27856_, _27853_);
  nor (_27859_, _27857_, _03178_);
  nor (_27860_, _27859_, _27803_);
  nor (_27861_, _27860_, _03600_);
  and (_27862_, _12733_, _05300_);
  or (_27863_, _27799_, _07766_);
  nor (_27864_, _27863_, _27862_);
  or (_27865_, _27864_, _03780_);
  nor (_27866_, _27865_, _27861_);
  nor (_27867_, _27866_, _27802_);
  nor (_27868_, _27867_, _03622_);
  nor (_27870_, _27799_, _05567_);
  not (_27871_, _27870_);
  nor (_27872_, _27855_, _07777_);
  and (_27873_, _27872_, _27871_);
  nor (_27874_, _27873_, _27868_);
  nor (_27875_, _27874_, _10754_);
  nor (_27876_, _27806_, _06828_);
  and (_27877_, _27876_, _27871_);
  nor (_27878_, _27877_, _27875_);
  and (_27879_, _27878_, _27798_);
  nor (_27881_, _12732_, _10706_);
  nor (_27882_, _27881_, _27799_);
  and (_27883_, _27882_, _03624_);
  nor (_27884_, _27883_, _27879_);
  nor (_27885_, _27884_, _03785_);
  nor (_27886_, _12738_, _10706_);
  or (_27887_, _27799_, _07793_);
  nor (_27888_, _27887_, _27886_);
  or (_27889_, _27888_, _03798_);
  nor (_27890_, _27889_, _27885_);
  nor (_27892_, _05970_, _03722_);
  nor (_27893_, _27892_, _05971_);
  nor (_27894_, _27893_, _10652_);
  or (_27895_, _27894_, _27890_);
  and (_27896_, _27895_, _06399_);
  or (_27897_, _27896_, _27796_);
  and (_27898_, _27897_, _03516_);
  nor (_27899_, _27893_, _03516_);
  or (_27900_, _27899_, _27898_);
  and (_27901_, _27900_, _04246_);
  nor (_27903_, _27816_, _04246_);
  nor (_27904_, _27903_, _05103_);
  not (_27905_, _27904_);
  nor (_27906_, _27905_, _27901_);
  nor (_27907_, _27906_, _27795_);
  and (_27908_, _27907_, _03514_);
  and (_27909_, _12794_, _05300_);
  nor (_27910_, _27909_, _27799_);
  nor (_27911_, _27910_, _03514_);
  or (_27912_, _27911_, _27908_);
  or (_27914_, _27912_, _43004_);
  or (_27915_, _43000_, \oc8051_golden_model_1.SP [3]);
  and (_27916_, _27915_, _41806_);
  and (_43609_, _27916_, _27914_);
  nor (_27917_, _05010_, \oc8051_golden_model_1.SP [4]);
  nor (_27918_, _27917_, _10645_);
  nor (_27919_, _27918_, _04540_);
  and (_27920_, _27918_, _03192_);
  nor (_27921_, _27920_, _03624_);
  nor (_27922_, _05300_, _10679_);
  and (_27924_, _12817_, _05300_);
  nor (_27925_, _27924_, _27922_);
  nor (_27926_, _27925_, _07778_);
  and (_27927_, _05011_, \oc8051_golden_model_1.SP [4]);
  nor (_27928_, _05011_, \oc8051_golden_model_1.SP [4]);
  nor (_27929_, _27928_, _27927_);
  and (_27930_, _27929_, _03508_);
  nor (_27931_, _04409_, _10679_);
  and (_27932_, _05300_, \oc8051_golden_model_1.ACC [4]);
  nor (_27933_, _27932_, _27922_);
  nor (_27935_, _27933_, _09029_);
  or (_27936_, _27935_, _27931_);
  and (_27937_, _27936_, _04763_);
  and (_27938_, _27918_, _03980_);
  nor (_27939_, _27938_, _27937_);
  nor (_27940_, _27939_, _03610_);
  nor (_27941_, _12841_, _10706_);
  nor (_27942_, _27941_, _27922_);
  nor (_27943_, _27942_, _04081_);
  or (_27944_, _27943_, _27940_);
  and (_27946_, _27944_, _03230_);
  and (_27947_, _27918_, _04768_);
  or (_27948_, _27947_, _27946_);
  and (_27949_, _27948_, _03996_);
  and (_27950_, _10680_, _03498_);
  nor (_27951_, _05972_, _10679_);
  nor (_27952_, _27951_, _27950_);
  nor (_27953_, _27952_, _03996_);
  or (_27954_, _27953_, _27949_);
  and (_27955_, _27954_, _03737_);
  nor (_27957_, _27933_, _03737_);
  or (_27958_, _27957_, _27955_);
  and (_27959_, _27958_, _03510_);
  or (_27960_, _27959_, _10694_);
  nor (_27961_, _27960_, _27930_);
  nor (_27962_, _27918_, _04767_);
  or (_27963_, _27962_, _07390_);
  nor (_27964_, _27963_, _27961_);
  nor (_27965_, _05777_, _10706_);
  nor (_27966_, _27965_, _27922_);
  nor (_27968_, _27966_, _06838_);
  nor (_27969_, _27968_, _04481_);
  not (_27970_, _27969_);
  nor (_27971_, _27970_, _27964_);
  and (_27972_, _06730_, _05300_);
  nor (_27973_, _27922_, _07400_);
  not (_27974_, _27973_);
  nor (_27975_, _27974_, _27972_);
  nor (_27976_, _27975_, _03222_);
  not (_27977_, _27976_);
  nor (_27979_, _27977_, _27971_);
  nor (_27980_, _12933_, _10706_);
  nor (_27981_, _27980_, _27922_);
  nor (_27982_, _27981_, _03589_);
  or (_27983_, _27982_, _27979_);
  and (_27984_, _27983_, _05886_);
  and (_27985_, _06298_, _05300_);
  nor (_27986_, _27985_, _27922_);
  nor (_27987_, _27986_, _05886_);
  or (_27988_, _27987_, _27984_);
  and (_27990_, _27988_, _10736_);
  and (_27991_, _27918_, _03178_);
  or (_27992_, _27991_, _03600_);
  nor (_27993_, _27992_, _27990_);
  and (_27994_, _12821_, _05300_);
  or (_27995_, _27922_, _07766_);
  nor (_27996_, _27995_, _27994_);
  or (_27997_, _27996_, _03780_);
  nor (_27998_, _27997_, _27993_);
  nor (_27999_, _27998_, _27926_);
  nor (_28001_, _27999_, _03622_);
  nor (_28002_, _27922_, _05825_);
  not (_28003_, _28002_);
  nor (_28004_, _27986_, _07777_);
  and (_28005_, _28004_, _28003_);
  nor (_28006_, _28005_, _28001_);
  nor (_28007_, _28006_, _10754_);
  nor (_28008_, _27933_, _06828_);
  and (_28009_, _28008_, _28003_);
  nor (_28010_, _28009_, _28007_);
  and (_28012_, _28010_, _27921_);
  nor (_28013_, _12819_, _10706_);
  nor (_28014_, _28013_, _27922_);
  and (_28015_, _28014_, _03624_);
  nor (_28016_, _28015_, _28012_);
  nor (_28017_, _28016_, _03785_);
  nor (_28018_, _12816_, _10706_);
  or (_28019_, _27922_, _07793_);
  nor (_28020_, _28019_, _28018_);
  or (_28021_, _28020_, _03798_);
  nor (_28023_, _28021_, _28017_);
  nor (_28024_, _05971_, _10679_);
  nor (_28025_, _28024_, _10680_);
  nor (_28026_, _28025_, _10652_);
  or (_28027_, _28026_, _28023_);
  and (_28028_, _28027_, _06399_);
  and (_28029_, _27918_, _03188_);
  or (_28030_, _28029_, _28028_);
  and (_28031_, _28030_, _03516_);
  nor (_28032_, _28025_, _03516_);
  or (_28034_, _28032_, _28031_);
  and (_28035_, _28034_, _04246_);
  nor (_28036_, _27942_, _04246_);
  nor (_28037_, _28036_, _05103_);
  not (_28038_, _28037_);
  nor (_28039_, _28038_, _28035_);
  nor (_28040_, _28039_, _27919_);
  and (_28041_, _28040_, _03514_);
  and (_28042_, _13003_, _05300_);
  nor (_28043_, _28042_, _27922_);
  nor (_28045_, _28043_, _03514_);
  or (_28046_, _28045_, _28041_);
  or (_28047_, _28046_, _43004_);
  or (_28048_, _43000_, \oc8051_golden_model_1.SP [4]);
  and (_28049_, _28048_, _41806_);
  and (_43610_, _28049_, _28047_);
  nor (_28050_, _10645_, \oc8051_golden_model_1.SP [5]);
  nor (_28051_, _28050_, _10646_);
  nor (_28052_, _28051_, _04540_);
  nor (_28053_, _05300_, _10678_);
  and (_28055_, _13147_, _05300_);
  nor (_28056_, _28055_, _28053_);
  nor (_28057_, _28056_, _07778_);
  nor (_28058_, _04409_, _10678_);
  and (_28059_, _05300_, \oc8051_golden_model_1.ACC [5]);
  nor (_28060_, _28059_, _28053_);
  nor (_28061_, _28060_, _09029_);
  or (_28062_, _28061_, _28058_);
  and (_28063_, _28062_, _04763_);
  and (_28064_, _28051_, _03980_);
  nor (_28066_, _28064_, _28063_);
  nor (_28067_, _28066_, _03610_);
  nor (_28068_, _13014_, _10706_);
  nor (_28069_, _28068_, _28053_);
  nor (_28070_, _28069_, _04081_);
  or (_28071_, _28070_, _28067_);
  and (_28072_, _28071_, _03230_);
  and (_28073_, _28051_, _04768_);
  or (_28074_, _28073_, _28072_);
  and (_28075_, _28074_, _03996_);
  and (_28077_, _10681_, _03498_);
  nor (_28078_, _27950_, _10678_);
  nor (_28079_, _28078_, _28077_);
  nor (_28080_, _28079_, _03996_);
  or (_28081_, _28080_, _28075_);
  and (_28082_, _28081_, _03737_);
  nor (_28083_, _28060_, _03737_);
  or (_28084_, _28083_, _28082_);
  and (_28085_, _28084_, _03510_);
  and (_28086_, _10646_, \oc8051_golden_model_1.SP [0]);
  nor (_28088_, _27927_, \oc8051_golden_model_1.SP [5]);
  nor (_28089_, _28088_, _28086_);
  and (_28090_, _28089_, _03508_);
  nor (_28091_, _28090_, _10694_);
  not (_28092_, _28091_);
  nor (_28093_, _28092_, _28085_);
  nor (_28094_, _28051_, _04767_);
  or (_28095_, _28094_, _07390_);
  nor (_28096_, _28095_, _28093_);
  nor (_28097_, _05469_, _10706_);
  nor (_28099_, _28097_, _28053_);
  nor (_28100_, _28099_, _06838_);
  nor (_28101_, _28100_, _04481_);
  not (_28102_, _28101_);
  nor (_28103_, _28102_, _28096_);
  and (_28104_, _06684_, _05300_);
  nor (_28105_, _28053_, _07400_);
  not (_28106_, _28105_);
  nor (_28107_, _28106_, _28104_);
  nor (_28108_, _28107_, _03222_);
  not (_28110_, _28108_);
  nor (_28111_, _28110_, _28103_);
  nor (_28112_, _13127_, _10706_);
  nor (_28113_, _28112_, _28053_);
  nor (_28114_, _28113_, _03589_);
  or (_28115_, _28114_, _28111_);
  and (_28116_, _28115_, _05886_);
  and (_28117_, _06306_, _05300_);
  nor (_28118_, _28117_, _28053_);
  nor (_28119_, _28118_, _05886_);
  or (_28121_, _28119_, _28116_);
  and (_28122_, _28121_, _10736_);
  and (_28123_, _28051_, _03178_);
  or (_28124_, _28123_, _03600_);
  nor (_28125_, _28124_, _28122_);
  and (_28126_, _13141_, _05300_);
  or (_28127_, _28053_, _07766_);
  nor (_28128_, _28127_, _28126_);
  or (_28129_, _28128_, _03780_);
  nor (_28130_, _28129_, _28125_);
  nor (_28132_, _28130_, _28057_);
  nor (_28133_, _28132_, _03622_);
  nor (_28134_, _28053_, _05518_);
  not (_28135_, _28134_);
  nor (_28136_, _28118_, _07777_);
  and (_28137_, _28136_, _28135_);
  nor (_28138_, _28137_, _28133_);
  nor (_28139_, _28138_, _10754_);
  nor (_28140_, _28060_, _06828_);
  and (_28141_, _28140_, _28135_);
  and (_28143_, _28051_, _03192_);
  nor (_28144_, _28143_, _28141_);
  and (_28145_, _28144_, _07795_);
  not (_28146_, _28145_);
  nor (_28147_, _28146_, _28139_);
  nor (_28148_, _13140_, _10706_);
  nor (_28149_, _28148_, _28053_);
  and (_28150_, _28149_, _03624_);
  nor (_28151_, _28150_, _28147_);
  nor (_28152_, _28151_, _03785_);
  nor (_28154_, _13146_, _10706_);
  or (_28155_, _28053_, _07793_);
  nor (_28156_, _28155_, _28154_);
  or (_28157_, _28156_, _03798_);
  nor (_28158_, _28157_, _28152_);
  nor (_28159_, _10680_, _10678_);
  nor (_28160_, _28159_, _10681_);
  nor (_28161_, _28160_, _10652_);
  or (_28162_, _28161_, _28158_);
  and (_28163_, _28162_, _06399_);
  and (_28165_, _28051_, _03188_);
  or (_28166_, _28165_, _28163_);
  and (_28167_, _28166_, _03516_);
  nor (_28168_, _28160_, _03516_);
  or (_28169_, _28168_, _28167_);
  and (_28170_, _28169_, _04246_);
  nor (_28171_, _28069_, _04246_);
  nor (_28172_, _28171_, _05103_);
  not (_28173_, _28172_);
  nor (_28174_, _28173_, _28170_);
  nor (_28176_, _28174_, _28052_);
  nor (_28177_, _28176_, _03447_);
  and (_28178_, _13199_, _05300_);
  nor (_28179_, _28178_, _28053_);
  and (_28180_, _28179_, _03447_);
  nor (_28181_, _28180_, _28177_);
  or (_28182_, _28181_, _43004_);
  or (_28183_, _43000_, \oc8051_golden_model_1.SP [5]);
  and (_28184_, _28183_, _41806_);
  and (_43611_, _28184_, _28182_);
  nor (_28186_, _05300_, _10677_);
  and (_28187_, _13353_, _05300_);
  nor (_28188_, _28187_, _28186_);
  nor (_28189_, _28188_, _07778_);
  and (_28190_, _06455_, _05300_);
  or (_28191_, _28190_, _28186_);
  and (_28192_, _28191_, _04481_);
  and (_28193_, _05300_, \oc8051_golden_model_1.ACC [6]);
  nor (_28194_, _28193_, _28186_);
  nor (_28195_, _28194_, _09029_);
  nor (_28197_, _04409_, _10677_);
  or (_28198_, _28197_, _03980_);
  nor (_28199_, _28198_, _28195_);
  nor (_28200_, _10646_, \oc8051_golden_model_1.SP [6]);
  nor (_28201_, _28200_, _10647_);
  not (_28202_, _28201_);
  and (_28203_, _28202_, _03980_);
  nor (_28204_, _28203_, _28199_);
  and (_28205_, _28204_, _04081_);
  nor (_28206_, _13242_, _10706_);
  nor (_28208_, _28206_, _28186_);
  nor (_28209_, _28208_, _04081_);
  or (_28210_, _28209_, _28205_);
  and (_28211_, _28210_, _03230_);
  nor (_28212_, _28202_, _03230_);
  or (_28213_, _28212_, _28211_);
  and (_28214_, _28213_, _03996_);
  nor (_28215_, _28077_, _10677_);
  nor (_28216_, _28215_, _10683_);
  nor (_28217_, _28216_, _03996_);
  or (_28219_, _28217_, _28214_);
  and (_28220_, _28219_, _03737_);
  nor (_28221_, _28194_, _03737_);
  or (_28222_, _28221_, _28220_);
  and (_28223_, _28222_, _03510_);
  nor (_28224_, _28086_, \oc8051_golden_model_1.SP [6]);
  nor (_28225_, _28224_, _10695_);
  and (_28226_, _28225_, _03508_);
  nor (_28227_, _28226_, _28223_);
  nor (_28228_, _28227_, _10694_);
  nor (_28230_, _28202_, _04767_);
  nor (_28231_, _28230_, _07390_);
  not (_28232_, _28231_);
  nor (_28233_, _28232_, _28228_);
  not (_28234_, _28186_);
  nor (_28235_, _05363_, _10706_);
  nor (_28236_, _28235_, _06838_);
  and (_28237_, _28236_, _28234_);
  or (_28238_, _28237_, _04481_);
  nor (_28239_, _28238_, _28233_);
  or (_28240_, _28239_, _28192_);
  and (_28241_, _28240_, _03589_);
  nor (_28242_, _13332_, _10706_);
  nor (_28243_, _28242_, _28186_);
  nor (_28244_, _28243_, _03589_);
  or (_28245_, _28244_, _03601_);
  or (_28246_, _28245_, _28241_);
  and (_28247_, _13339_, _05300_);
  nor (_28248_, _28247_, _28186_);
  nand (_28249_, _28248_, _03601_);
  and (_28252_, _28249_, _28246_);
  nor (_28253_, _28252_, _03178_);
  and (_28254_, _28202_, _03178_);
  nor (_28255_, _28254_, _28253_);
  nor (_28256_, _28255_, _03600_);
  and (_28257_, _13347_, _05300_);
  or (_28258_, _28186_, _07766_);
  nor (_28259_, _28258_, _28257_);
  or (_28260_, _28259_, _03780_);
  nor (_28261_, _28260_, _28256_);
  nor (_28263_, _28261_, _28189_);
  nor (_28264_, _28263_, _03622_);
  and (_28265_, _28234_, _05411_);
  not (_28266_, _28265_);
  nor (_28267_, _28248_, _07777_);
  and (_28268_, _28267_, _28266_);
  nor (_28269_, _28268_, _28264_);
  nor (_28270_, _28269_, _10754_);
  and (_28271_, _28201_, _03192_);
  or (_28272_, _28265_, _06828_);
  nor (_28274_, _28272_, _28194_);
  nor (_28275_, _28274_, _28271_);
  and (_28276_, _28275_, _07795_);
  not (_28277_, _28276_);
  nor (_28278_, _28277_, _28270_);
  nor (_28279_, _13346_, _10706_);
  nor (_28280_, _28279_, _28186_);
  and (_28281_, _28280_, _03624_);
  nor (_28282_, _28281_, _28278_);
  and (_28283_, _28282_, _07793_);
  nor (_28285_, _13352_, _10706_);
  nor (_28286_, _28285_, _28186_);
  nor (_28287_, _28286_, _07793_);
  or (_28288_, _28287_, _28283_);
  and (_28289_, _28288_, _10652_);
  nor (_28290_, _10681_, _10677_);
  nor (_28291_, _28290_, _10682_);
  not (_28292_, _28291_);
  nor (_28293_, _28292_, _03188_);
  nor (_28294_, _28293_, _10774_);
  nor (_28296_, _28294_, _28289_);
  and (_28297_, _28202_, _03188_);
  or (_28298_, _28297_, _03515_);
  nor (_28299_, _28298_, _28296_);
  and (_28300_, _28292_, _03515_);
  or (_28301_, _28300_, _03815_);
  nor (_28302_, _28301_, _28299_);
  and (_28303_, _28208_, _03815_);
  nor (_28304_, _28303_, _05103_);
  not (_28305_, _28304_);
  nor (_28307_, _28305_, _28302_);
  nor (_28308_, _28202_, _04540_);
  nor (_28309_, _28308_, _03447_);
  not (_28310_, _28309_);
  nor (_28311_, _28310_, _28307_);
  and (_28312_, _13402_, _05300_);
  or (_28313_, _28186_, _03514_);
  nor (_28314_, _28313_, _28312_);
  nor (_28315_, _28314_, _28311_);
  or (_28316_, _28315_, _43004_);
  or (_28318_, _43000_, \oc8051_golden_model_1.SP [6]);
  and (_28319_, _28318_, _41806_);
  and (_43612_, _28319_, _28316_);
  not (_28320_, \oc8051_golden_model_1.TCON [0]);
  nor (_28321_, _05258_, _28320_);
  and (_28322_, _12128_, _05258_);
  nor (_28323_, _28322_, _28321_);
  nor (_28324_, _28323_, _07778_);
  and (_28325_, _05258_, _06274_);
  nor (_28326_, _28325_, _28321_);
  and (_28328_, _28326_, _03601_);
  and (_28329_, _05258_, _04620_);
  nor (_28330_, _28329_, _28321_);
  and (_28331_, _28330_, _07390_);
  and (_28332_, _05258_, \oc8051_golden_model_1.ACC [0]);
  nor (_28333_, _28332_, _28321_);
  nor (_28334_, _28333_, _09029_);
  nor (_28335_, _04409_, _28320_);
  or (_28336_, _28335_, _28334_);
  and (_28337_, _28336_, _04081_);
  nor (_28339_, _05666_, _10802_);
  nor (_28340_, _28339_, _28321_);
  nor (_28341_, _28340_, _04081_);
  or (_28342_, _28341_, _28337_);
  and (_28343_, _28342_, _04055_);
  nor (_28344_, _05927_, _28320_);
  and (_28345_, _12021_, _05927_);
  nor (_28346_, _28345_, _28344_);
  nor (_28347_, _28346_, _04055_);
  nor (_28348_, _28347_, _28343_);
  nor (_28350_, _28348_, _03723_);
  nor (_28351_, _28330_, _03996_);
  or (_28352_, _28351_, _28350_);
  and (_28353_, _28352_, _03737_);
  nor (_28354_, _28333_, _03737_);
  or (_28355_, _28354_, _28353_);
  and (_28356_, _28355_, _03736_);
  and (_28357_, _28321_, _03714_);
  or (_28358_, _28357_, _28356_);
  and (_28359_, _28358_, _06840_);
  nor (_28361_, _28340_, _06840_);
  or (_28362_, _28361_, _28359_);
  and (_28363_, _28362_, _03710_);
  nor (_28364_, _12052_, _10839_);
  nor (_28365_, _28364_, _28344_);
  nor (_28366_, _28365_, _03710_);
  or (_28367_, _28366_, _07390_);
  nor (_28368_, _28367_, _28363_);
  nor (_28369_, _28368_, _28331_);
  nor (_28370_, _28369_, _04481_);
  and (_28372_, _06546_, _05258_);
  nor (_28373_, _28321_, _07400_);
  not (_28374_, _28373_);
  nor (_28375_, _28374_, _28372_);
  or (_28376_, _28375_, _03222_);
  nor (_28377_, _28376_, _28370_);
  nor (_28378_, _12109_, _10802_);
  nor (_28379_, _28378_, _28321_);
  nor (_28380_, _28379_, _03589_);
  or (_28381_, _28380_, _03601_);
  nor (_28383_, _28381_, _28377_);
  nor (_28384_, _28383_, _28328_);
  or (_28385_, _28384_, _03600_);
  and (_28386_, _12124_, _05258_);
  or (_28387_, _28386_, _28321_);
  or (_28388_, _28387_, _07766_);
  and (_28389_, _28388_, _07778_);
  and (_28390_, _28389_, _28385_);
  nor (_28391_, _28390_, _28324_);
  nor (_28392_, _28391_, _03622_);
  or (_28394_, _28326_, _07777_);
  nor (_28395_, _28394_, _28339_);
  nor (_28396_, _28395_, _28392_);
  nor (_28397_, _28396_, _03790_);
  and (_28398_, _12005_, _05258_);
  or (_28399_, _28398_, _28321_);
  and (_28400_, _28399_, _03790_);
  or (_28401_, _28400_, _28397_);
  and (_28402_, _28401_, _07795_);
  nor (_28403_, _12122_, _10802_);
  nor (_28405_, _28403_, _28321_);
  nor (_28406_, _28405_, _07795_);
  or (_28407_, _28406_, _28402_);
  and (_28408_, _28407_, _07793_);
  nor (_28409_, _12003_, _10802_);
  nor (_28410_, _28409_, _28321_);
  nor (_28411_, _28410_, _07793_);
  or (_28412_, _28411_, _28408_);
  and (_28413_, _28412_, _04246_);
  nor (_28414_, _28340_, _04246_);
  or (_28416_, _28414_, _28413_);
  and (_28417_, _28416_, _03823_);
  and (_28418_, _28321_, _03453_);
  nor (_28419_, _28418_, _03447_);
  not (_28420_, _28419_);
  nor (_28421_, _28420_, _28417_);
  and (_28422_, _28340_, _03447_);
  or (_28423_, _28422_, _28421_);
  nand (_28424_, _28423_, _43000_);
  or (_28425_, _43000_, \oc8051_golden_model_1.TCON [0]);
  and (_28426_, _28425_, _41806_);
  and (_43613_, _28426_, _28424_);
  or (_28427_, _05258_, \oc8051_golden_model_1.TCON [1]);
  and (_28428_, _12213_, _05258_);
  not (_28429_, _28428_);
  and (_28430_, _28429_, _28427_);
  or (_28431_, _28430_, _04081_);
  nand (_28432_, _05258_, _03274_);
  and (_28433_, _28432_, _28427_);
  and (_28434_, _28433_, _04409_);
  not (_28437_, \oc8051_golden_model_1.TCON [1]);
  nor (_28438_, _04409_, _28437_);
  or (_28439_, _28438_, _03610_);
  or (_28440_, _28439_, _28434_);
  and (_28441_, _28440_, _04055_);
  and (_28442_, _28441_, _28431_);
  and (_28443_, _12224_, _05927_);
  nor (_28444_, _05927_, _28437_);
  or (_28445_, _28444_, _03723_);
  or (_28446_, _28445_, _28443_);
  and (_28448_, _28446_, _14265_);
  or (_28449_, _28448_, _28442_);
  nor (_28450_, _05258_, _28437_);
  and (_28451_, _05258_, _06764_);
  or (_28452_, _28451_, _28450_);
  or (_28453_, _28452_, _03996_);
  and (_28454_, _28453_, _28449_);
  or (_28455_, _28454_, _03729_);
  or (_28456_, _28433_, _03737_);
  and (_28457_, _28456_, _03736_);
  and (_28459_, _28457_, _28455_);
  and (_28460_, _12211_, _05927_);
  or (_28461_, _28460_, _28444_);
  and (_28462_, _28461_, _03714_);
  or (_28463_, _28462_, _03719_);
  or (_28464_, _28463_, _28459_);
  and (_28465_, _28443_, _12239_);
  or (_28466_, _28444_, _06840_);
  or (_28467_, _28466_, _28465_);
  and (_28468_, _28467_, _28464_);
  and (_28470_, _28468_, _03710_);
  nor (_28471_, _12256_, _10839_);
  or (_28472_, _28444_, _28471_);
  and (_28473_, _28472_, _03505_);
  or (_28474_, _28473_, _07390_);
  or (_28475_, _28474_, _28470_);
  or (_28476_, _28452_, _06838_);
  and (_28477_, _28476_, _28475_);
  or (_28478_, _28477_, _04481_);
  and (_28479_, _06501_, _05258_);
  or (_28481_, _28450_, _07400_);
  or (_28482_, _28481_, _28479_);
  and (_28483_, _28482_, _03589_);
  and (_28484_, _28483_, _28478_);
  nor (_28485_, _12313_, _10802_);
  or (_28486_, _28485_, _28450_);
  and (_28487_, _28486_, _03222_);
  or (_28488_, _28487_, _28484_);
  and (_28489_, _28488_, _03602_);
  or (_28490_, _12327_, _10802_);
  and (_28492_, _28490_, _03600_);
  nand (_28493_, _05258_, _04303_);
  and (_28494_, _28493_, _03601_);
  or (_28495_, _28494_, _28492_);
  and (_28496_, _28495_, _28427_);
  or (_28497_, _28496_, _28489_);
  and (_28498_, _28497_, _07778_);
  or (_28499_, _12333_, _10802_);
  and (_28500_, _28427_, _03780_);
  and (_28501_, _28500_, _28499_);
  or (_28503_, _28501_, _28498_);
  and (_28504_, _28503_, _07777_);
  or (_28505_, _12207_, _10802_);
  and (_28506_, _28427_, _03622_);
  and (_28507_, _28506_, _28505_);
  or (_28508_, _28507_, _28504_);
  and (_28509_, _28508_, _06828_);
  or (_28510_, _28450_, _05618_);
  and (_28511_, _28433_, _03790_);
  and (_28512_, _28511_, _28510_);
  or (_28514_, _28512_, _28509_);
  and (_28515_, _28514_, _03786_);
  or (_28516_, _28493_, _05618_);
  and (_28517_, _28427_, _03624_);
  and (_28518_, _28517_, _28516_);
  or (_28519_, _28432_, _05618_);
  and (_28520_, _28427_, _03785_);
  and (_28521_, _28520_, _28519_);
  or (_28522_, _28521_, _03815_);
  or (_28523_, _28522_, _28518_);
  or (_28525_, _28523_, _28515_);
  or (_28526_, _28430_, _04246_);
  and (_28527_, _28526_, _03823_);
  and (_28528_, _28527_, _28525_);
  and (_28529_, _28461_, _03453_);
  or (_28530_, _28529_, _03447_);
  or (_28531_, _28530_, _28528_);
  or (_28532_, _28450_, _03514_);
  or (_28533_, _28532_, _28428_);
  and (_28534_, _28533_, _28531_);
  and (_28536_, _28534_, _43000_);
  nor (_28537_, \oc8051_golden_model_1.TCON [1], rst);
  nor (_28538_, _28537_, _00000_);
  or (_43614_, _28538_, _28536_);
  not (_28539_, \oc8051_golden_model_1.TCON [2]);
  nor (_28540_, _05258_, _28539_);
  and (_28541_, _05258_, _06332_);
  nor (_28542_, _28541_, _28540_);
  and (_28543_, _28542_, _03601_);
  nor (_28544_, _10802_, _04875_);
  nor (_28546_, _28544_, _28540_);
  and (_28547_, _28546_, _07390_);
  and (_28548_, _05258_, \oc8051_golden_model_1.ACC [2]);
  nor (_28549_, _28548_, _28540_);
  nor (_28550_, _28549_, _09029_);
  nor (_28551_, _04409_, _28539_);
  or (_28552_, _28551_, _28550_);
  and (_28553_, _28552_, _04081_);
  nor (_28554_, _12416_, _10802_);
  nor (_28555_, _28554_, _28540_);
  nor (_28557_, _28555_, _04081_);
  or (_28558_, _28557_, _28553_);
  and (_28559_, _28558_, _04055_);
  nor (_28560_, _05927_, _28539_);
  and (_28561_, _12411_, _05927_);
  nor (_28562_, _28561_, _28560_);
  nor (_28563_, _28562_, _04055_);
  or (_28564_, _28563_, _28559_);
  and (_28565_, _28564_, _03996_);
  nor (_28566_, _28546_, _03996_);
  or (_28568_, _28566_, _28565_);
  and (_28569_, _28568_, _03737_);
  nor (_28570_, _28549_, _03737_);
  or (_28571_, _28570_, _28569_);
  and (_28572_, _28571_, _03736_);
  and (_28573_, _12409_, _05927_);
  nor (_28574_, _28573_, _28560_);
  nor (_28575_, _28574_, _03736_);
  or (_28576_, _28575_, _03719_);
  or (_28577_, _28576_, _28572_);
  and (_28579_, _28561_, _12443_);
  or (_28580_, _28560_, _06840_);
  or (_28581_, _28580_, _28579_);
  and (_28582_, _28581_, _03710_);
  and (_28583_, _28582_, _28577_);
  nor (_28584_, _12461_, _10839_);
  nor (_28585_, _28584_, _28560_);
  nor (_28586_, _28585_, _03710_);
  nor (_28587_, _28586_, _07390_);
  not (_28588_, _28587_);
  nor (_28590_, _28588_, _28583_);
  nor (_28591_, _28590_, _28547_);
  nor (_28592_, _28591_, _04481_);
  and (_28593_, _06637_, _05258_);
  nor (_28594_, _28540_, _07400_);
  not (_28595_, _28594_);
  nor (_28596_, _28595_, _28593_);
  or (_28597_, _28596_, _03222_);
  nor (_28598_, _28597_, _28592_);
  nor (_28599_, _12519_, _10802_);
  nor (_28601_, _28540_, _28599_);
  nor (_28602_, _28601_, _03589_);
  or (_28603_, _28602_, _03601_);
  nor (_28604_, _28603_, _28598_);
  nor (_28605_, _28604_, _28543_);
  or (_28606_, _28605_, _03600_);
  and (_28607_, _12533_, _05258_);
  or (_28608_, _28607_, _28540_);
  or (_28609_, _28608_, _07766_);
  and (_28610_, _28609_, _07778_);
  and (_28612_, _28610_, _28606_);
  and (_28613_, _12539_, _05258_);
  nor (_28614_, _28613_, _28540_);
  nor (_28615_, _28614_, _07778_);
  nor (_28616_, _28615_, _28612_);
  nor (_28617_, _28616_, _03622_);
  nor (_28618_, _28540_, _05718_);
  not (_28619_, _28618_);
  nor (_28620_, _28542_, _07777_);
  and (_28621_, _28620_, _28619_);
  nor (_28623_, _28621_, _28617_);
  nor (_28624_, _28623_, _03790_);
  nor (_28625_, _28549_, _06828_);
  and (_28626_, _28625_, _28619_);
  or (_28627_, _28626_, _28624_);
  and (_28628_, _28627_, _07795_);
  nor (_28629_, _12532_, _10802_);
  nor (_28630_, _28629_, _28540_);
  nor (_28631_, _28630_, _07795_);
  or (_28632_, _28631_, _28628_);
  and (_28634_, _28632_, _07793_);
  nor (_28635_, _12538_, _10802_);
  nor (_28636_, _28635_, _28540_);
  nor (_28637_, _28636_, _07793_);
  or (_28638_, _28637_, _28634_);
  and (_28639_, _28638_, _04246_);
  nor (_28640_, _28555_, _04246_);
  or (_28641_, _28640_, _28639_);
  and (_28642_, _28641_, _03823_);
  nor (_28643_, _28574_, _03823_);
  or (_28645_, _28643_, _28642_);
  and (_28646_, _28645_, _03514_);
  and (_28647_, _12592_, _05258_);
  nor (_28648_, _28647_, _28540_);
  nor (_28649_, _28648_, _03514_);
  or (_28650_, _28649_, _28646_);
  or (_28651_, _28650_, _43004_);
  or (_28652_, _43000_, \oc8051_golden_model_1.TCON [2]);
  and (_28653_, _28652_, _41806_);
  and (_43615_, _28653_, _28651_);
  not (_28655_, \oc8051_golden_model_1.TCON [3]);
  nor (_28656_, _05258_, _28655_);
  and (_28657_, _05258_, _06276_);
  nor (_28658_, _28657_, _28656_);
  and (_28659_, _28658_, _03601_);
  nor (_28660_, _10802_, _05005_);
  nor (_28661_, _28660_, _28656_);
  and (_28662_, _28661_, _07390_);
  and (_28663_, _05258_, \oc8051_golden_model_1.ACC [3]);
  nor (_28664_, _28663_, _28656_);
  nor (_28666_, _28664_, _09029_);
  nor (_28667_, _04409_, _28655_);
  or (_28668_, _28667_, _28666_);
  and (_28669_, _28668_, _04081_);
  nor (_28670_, _12627_, _10802_);
  nor (_28671_, _28670_, _28656_);
  nor (_28672_, _28671_, _04081_);
  or (_28673_, _28672_, _28669_);
  and (_28674_, _28673_, _04055_);
  nor (_28675_, _05927_, _28655_);
  and (_28677_, _12631_, _05927_);
  nor (_28678_, _28677_, _28675_);
  nor (_28679_, _28678_, _04055_);
  or (_28680_, _28679_, _03723_);
  or (_28681_, _28680_, _28674_);
  nand (_28682_, _28661_, _03723_);
  and (_28683_, _28682_, _28681_);
  and (_28684_, _28683_, _03737_);
  nor (_28685_, _28664_, _03737_);
  or (_28686_, _28685_, _28684_);
  and (_28688_, _28686_, _03736_);
  and (_28689_, _12641_, _05927_);
  nor (_28690_, _28689_, _28675_);
  nor (_28691_, _28690_, _03736_);
  or (_28692_, _28691_, _28688_);
  and (_28693_, _28692_, _06840_);
  nor (_28694_, _28675_, _12648_);
  nor (_28695_, _28694_, _28678_);
  and (_28696_, _28695_, _03719_);
  or (_28697_, _28696_, _28693_);
  and (_28699_, _28697_, _03710_);
  nor (_28700_, _12612_, _10839_);
  nor (_28701_, _28700_, _28675_);
  nor (_28702_, _28701_, _03710_);
  nor (_28703_, _28702_, _07390_);
  not (_28704_, _28703_);
  nor (_28705_, _28704_, _28699_);
  nor (_28706_, _28705_, _28662_);
  nor (_28707_, _28706_, _04481_);
  and (_28708_, _06592_, _05258_);
  nor (_28710_, _28656_, _07400_);
  not (_28711_, _28710_);
  nor (_28712_, _28711_, _28708_);
  or (_28713_, _28712_, _03222_);
  nor (_28714_, _28713_, _28707_);
  nor (_28715_, _12718_, _10802_);
  nor (_28716_, _28656_, _28715_);
  nor (_28717_, _28716_, _03589_);
  or (_28718_, _28717_, _03601_);
  nor (_28719_, _28718_, _28714_);
  nor (_28721_, _28719_, _28659_);
  or (_28722_, _28721_, _03600_);
  and (_28723_, _12733_, _05258_);
  or (_28724_, _28723_, _28656_);
  or (_28725_, _28724_, _07766_);
  and (_28726_, _28725_, _07778_);
  and (_28727_, _28726_, _28722_);
  and (_28728_, _12739_, _05258_);
  nor (_28729_, _28728_, _28656_);
  nor (_28730_, _28729_, _07778_);
  nor (_28732_, _28730_, _28727_);
  nor (_28733_, _28732_, _03622_);
  nor (_28734_, _28656_, _05567_);
  not (_28735_, _28734_);
  nor (_28736_, _28658_, _07777_);
  and (_28737_, _28736_, _28735_);
  nor (_28738_, _28737_, _28733_);
  nor (_28739_, _28738_, _03790_);
  nor (_28740_, _28664_, _06828_);
  and (_28741_, _28740_, _28735_);
  or (_28743_, _28741_, _28739_);
  and (_28744_, _28743_, _07795_);
  nor (_28745_, _12732_, _10802_);
  nor (_28746_, _28745_, _28656_);
  nor (_28747_, _28746_, _07795_);
  or (_28748_, _28747_, _28744_);
  and (_28749_, _28748_, _07793_);
  nor (_28750_, _12738_, _10802_);
  nor (_28751_, _28750_, _28656_);
  nor (_28752_, _28751_, _07793_);
  or (_28754_, _28752_, _28749_);
  and (_28755_, _28754_, _04246_);
  nor (_28756_, _28671_, _04246_);
  or (_28757_, _28756_, _28755_);
  and (_28758_, _28757_, _03823_);
  nor (_28759_, _28690_, _03823_);
  nor (_28760_, _28759_, _03447_);
  not (_28761_, _28760_);
  nor (_28762_, _28761_, _28758_);
  and (_28763_, _12794_, _05258_);
  or (_28765_, _28656_, _03514_);
  nor (_28766_, _28765_, _28763_);
  nor (_28767_, _28766_, _28762_);
  or (_28768_, _28767_, _43004_);
  or (_28769_, _43000_, \oc8051_golden_model_1.TCON [3]);
  and (_28770_, _28769_, _41806_);
  and (_43618_, _28770_, _28768_);
  not (_28771_, \oc8051_golden_model_1.TCON [4]);
  nor (_28772_, _05258_, _28771_);
  nor (_28773_, _05777_, _10802_);
  nor (_28775_, _28773_, _28772_);
  and (_28776_, _28775_, _07390_);
  nor (_28777_, _05927_, _28771_);
  and (_28778_, _12827_, _05927_);
  nor (_28779_, _28778_, _28777_);
  nor (_28780_, _28779_, _03736_);
  and (_28781_, _05258_, \oc8051_golden_model_1.ACC [4]);
  nor (_28782_, _28781_, _28772_);
  nor (_28783_, _28782_, _09029_);
  nor (_28784_, _04409_, _28771_);
  or (_28786_, _28784_, _28783_);
  and (_28787_, _28786_, _04081_);
  nor (_28788_, _12841_, _10802_);
  nor (_28789_, _28788_, _28772_);
  nor (_28790_, _28789_, _04081_);
  or (_28791_, _28790_, _28787_);
  and (_28792_, _28791_, _04055_);
  and (_28793_, _12845_, _05927_);
  nor (_28794_, _28793_, _28777_);
  nor (_28795_, _28794_, _04055_);
  or (_28797_, _28795_, _03723_);
  or (_28798_, _28797_, _28792_);
  nand (_28799_, _28775_, _03723_);
  and (_28800_, _28799_, _28798_);
  and (_28801_, _28800_, _03737_);
  nor (_28802_, _28782_, _03737_);
  or (_28803_, _28802_, _28801_);
  and (_28804_, _28803_, _03736_);
  nor (_28805_, _28804_, _28780_);
  nor (_28806_, _28805_, _03719_);
  nor (_28807_, _28777_, _12860_);
  or (_28808_, _28794_, _06840_);
  nor (_28809_, _28808_, _28807_);
  nor (_28810_, _28809_, _28806_);
  nor (_28811_, _28810_, _03505_);
  nor (_28812_, _12825_, _10839_);
  nor (_28813_, _28812_, _28777_);
  nor (_28814_, _28813_, _03710_);
  nor (_28815_, _28814_, _07390_);
  not (_28816_, _28815_);
  nor (_28818_, _28816_, _28811_);
  nor (_28819_, _28818_, _28776_);
  nor (_28820_, _28819_, _04481_);
  and (_28821_, _06730_, _05258_);
  nor (_28822_, _28772_, _07400_);
  not (_28823_, _28822_);
  nor (_28824_, _28823_, _28821_);
  nor (_28825_, _28824_, _03222_);
  not (_28826_, _28825_);
  nor (_28827_, _28826_, _28820_);
  nor (_28829_, _12933_, _10802_);
  nor (_28830_, _28829_, _28772_);
  nor (_28831_, _28830_, _03589_);
  or (_28832_, _28831_, _08828_);
  or (_28833_, _28832_, _28827_);
  and (_28834_, _12821_, _05258_);
  or (_28835_, _28772_, _07766_);
  or (_28836_, _28835_, _28834_);
  and (_28837_, _06298_, _05258_);
  nor (_28838_, _28837_, _28772_);
  and (_28840_, _28838_, _03601_);
  nor (_28841_, _28840_, _03780_);
  and (_28842_, _28841_, _28836_);
  and (_28843_, _28842_, _28833_);
  and (_28844_, _12817_, _05258_);
  nor (_28845_, _28844_, _28772_);
  nor (_28846_, _28845_, _07778_);
  nor (_28847_, _28846_, _28843_);
  nor (_28848_, _28847_, _03622_);
  nor (_28849_, _28772_, _05825_);
  not (_28851_, _28849_);
  nor (_28852_, _28838_, _07777_);
  and (_28853_, _28852_, _28851_);
  nor (_28854_, _28853_, _28848_);
  nor (_28855_, _28854_, _03790_);
  nor (_28856_, _28782_, _06828_);
  and (_28857_, _28856_, _28851_);
  or (_28858_, _28857_, _28855_);
  and (_28859_, _28858_, _07795_);
  nor (_28860_, _12819_, _10802_);
  nor (_28862_, _28860_, _28772_);
  nor (_28863_, _28862_, _07795_);
  or (_28864_, _28863_, _28859_);
  and (_28865_, _28864_, _07793_);
  nor (_28866_, _12816_, _10802_);
  nor (_28867_, _28866_, _28772_);
  nor (_28868_, _28867_, _07793_);
  or (_28869_, _28868_, _28865_);
  and (_28870_, _28869_, _04246_);
  nor (_28871_, _28789_, _04246_);
  or (_28873_, _28871_, _28870_);
  and (_28874_, _28873_, _03823_);
  nor (_28875_, _28779_, _03823_);
  nor (_28876_, _28875_, _03447_);
  not (_28877_, _28876_);
  nor (_28878_, _28877_, _28874_);
  and (_28879_, _13003_, _05258_);
  or (_28880_, _28772_, _03514_);
  nor (_28881_, _28880_, _28879_);
  nor (_28882_, _28881_, _28878_);
  or (_28884_, _28882_, _43004_);
  or (_28885_, _43000_, \oc8051_golden_model_1.TCON [4]);
  and (_28886_, _28885_, _41806_);
  and (_43619_, _28886_, _28884_);
  not (_28887_, \oc8051_golden_model_1.TCON [5]);
  nor (_28888_, _05258_, _28887_);
  and (_28889_, _06684_, _05258_);
  or (_28890_, _28889_, _28888_);
  and (_28891_, _28890_, _04481_);
  and (_28892_, _05258_, \oc8051_golden_model_1.ACC [5]);
  nor (_28894_, _28892_, _28888_);
  nor (_28895_, _28894_, _09029_);
  nor (_28896_, _04409_, _28887_);
  or (_28897_, _28896_, _28895_);
  and (_28898_, _28897_, _04081_);
  nor (_28899_, _13014_, _10802_);
  nor (_28900_, _28899_, _28888_);
  nor (_28901_, _28900_, _04081_);
  or (_28902_, _28901_, _28898_);
  and (_28903_, _28902_, _04055_);
  nor (_28905_, _05927_, _28887_);
  and (_28906_, _13037_, _05927_);
  nor (_28907_, _28906_, _28905_);
  nor (_28908_, _28907_, _04055_);
  or (_28909_, _28908_, _03723_);
  or (_28910_, _28909_, _28903_);
  nor (_28911_, _05469_, _10802_);
  nor (_28912_, _28911_, _28888_);
  nand (_28913_, _28912_, _03723_);
  and (_28914_, _28913_, _28910_);
  and (_28916_, _28914_, _03737_);
  nor (_28917_, _28894_, _03737_);
  or (_28918_, _28917_, _28916_);
  and (_28919_, _28918_, _03736_);
  and (_28920_, _13047_, _05927_);
  nor (_28921_, _28920_, _28905_);
  nor (_28922_, _28921_, _03736_);
  or (_28923_, _28922_, _03719_);
  or (_28924_, _28923_, _28919_);
  nor (_28925_, _28905_, _13054_);
  nor (_28927_, _28925_, _28907_);
  or (_28928_, _28927_, _06840_);
  and (_28929_, _28928_, _03710_);
  and (_28930_, _28929_, _28924_);
  nor (_28931_, _13020_, _10839_);
  nor (_28932_, _28931_, _28905_);
  nor (_28933_, _28932_, _03710_);
  nor (_28934_, _28933_, _07390_);
  not (_28935_, _28934_);
  nor (_28936_, _28935_, _28930_);
  and (_28938_, _28912_, _07390_);
  or (_28939_, _28938_, _04481_);
  nor (_28940_, _28939_, _28936_);
  or (_28941_, _28940_, _28891_);
  and (_28942_, _28941_, _03589_);
  nor (_28943_, _13127_, _10802_);
  nor (_28944_, _28943_, _28888_);
  nor (_28945_, _28944_, _03589_);
  or (_28946_, _28945_, _08828_);
  or (_28947_, _28946_, _28942_);
  and (_28949_, _13141_, _05258_);
  or (_28950_, _28888_, _07766_);
  or (_28951_, _28950_, _28949_);
  and (_28952_, _06306_, _05258_);
  nor (_28953_, _28952_, _28888_);
  and (_28954_, _28953_, _03601_);
  nor (_28955_, _28954_, _03780_);
  and (_28956_, _28955_, _28951_);
  and (_28957_, _28956_, _28947_);
  and (_28958_, _13147_, _05258_);
  nor (_28959_, _28958_, _28888_);
  nor (_28960_, _28959_, _07778_);
  nor (_28961_, _28960_, _28957_);
  nor (_28962_, _28961_, _03622_);
  nor (_28963_, _28888_, _05518_);
  not (_28964_, _28963_);
  nor (_28965_, _28953_, _07777_);
  and (_28966_, _28965_, _28964_);
  nor (_28967_, _28966_, _28962_);
  nor (_28968_, _28967_, _03790_);
  nor (_28971_, _28894_, _06828_);
  and (_28972_, _28971_, _28964_);
  nor (_28973_, _28972_, _03624_);
  not (_28974_, _28973_);
  nor (_28975_, _28974_, _28968_);
  nor (_28976_, _13140_, _10802_);
  or (_28977_, _28888_, _07795_);
  nor (_28978_, _28977_, _28976_);
  or (_28979_, _28978_, _03785_);
  nor (_28980_, _28979_, _28975_);
  nor (_28982_, _13146_, _10802_);
  nor (_28983_, _28982_, _28888_);
  nor (_28984_, _28983_, _07793_);
  or (_28985_, _28984_, _28980_);
  and (_28986_, _28985_, _04246_);
  nor (_28987_, _28900_, _04246_);
  or (_28988_, _28987_, _28986_);
  and (_28989_, _28988_, _03823_);
  nor (_28990_, _28921_, _03823_);
  or (_28991_, _28990_, _28989_);
  and (_28993_, _28991_, _03514_);
  and (_28994_, _13199_, _05258_);
  nor (_28995_, _28994_, _28888_);
  nor (_28996_, _28995_, _03514_);
  or (_28997_, _28996_, _28993_);
  or (_28998_, _28997_, _43004_);
  or (_28999_, _43000_, \oc8051_golden_model_1.TCON [5]);
  and (_29000_, _28999_, _41806_);
  and (_43620_, _29000_, _28998_);
  not (_29001_, \oc8051_golden_model_1.TCON [6]);
  nor (_29003_, _05258_, _29001_);
  and (_29004_, _06455_, _05258_);
  or (_29005_, _29004_, _29003_);
  and (_29006_, _29005_, _04481_);
  and (_29007_, _05258_, \oc8051_golden_model_1.ACC [6]);
  nor (_29008_, _29007_, _29003_);
  nor (_29009_, _29008_, _09029_);
  nor (_29010_, _04409_, _29001_);
  or (_29011_, _29010_, _29009_);
  and (_29012_, _29011_, _04081_);
  nor (_29014_, _13242_, _10802_);
  nor (_29015_, _29014_, _29003_);
  nor (_29016_, _29015_, _04081_);
  or (_29017_, _29016_, _29012_);
  and (_29018_, _29017_, _04055_);
  nor (_29019_, _05927_, _29001_);
  and (_29020_, _13229_, _05927_);
  nor (_29021_, _29020_, _29019_);
  nor (_29022_, _29021_, _04055_);
  or (_29023_, _29022_, _03723_);
  or (_29025_, _29023_, _29018_);
  nor (_29026_, _05363_, _10802_);
  nor (_29027_, _29026_, _29003_);
  nand (_29028_, _29027_, _03723_);
  and (_29029_, _29028_, _29025_);
  and (_29030_, _29029_, _03737_);
  nor (_29031_, _29008_, _03737_);
  or (_29032_, _29031_, _29030_);
  and (_29033_, _29032_, _03736_);
  and (_29034_, _13253_, _05927_);
  nor (_29036_, _29034_, _29019_);
  nor (_29037_, _29036_, _03736_);
  or (_29038_, _29037_, _29033_);
  and (_29039_, _29038_, _06840_);
  nor (_29040_, _29019_, _13260_);
  nor (_29041_, _29040_, _29021_);
  and (_29042_, _29041_, _03719_);
  or (_29043_, _29042_, _29039_);
  and (_29044_, _29043_, _03710_);
  nor (_29045_, _13226_, _10839_);
  nor (_29047_, _29045_, _29019_);
  nor (_29048_, _29047_, _03710_);
  nor (_29049_, _29048_, _07390_);
  not (_29050_, _29049_);
  nor (_29051_, _29050_, _29044_);
  and (_29052_, _29027_, _07390_);
  or (_29053_, _29052_, _04481_);
  nor (_29054_, _29053_, _29051_);
  or (_29055_, _29054_, _29006_);
  and (_29056_, _29055_, _03589_);
  nor (_29058_, _13332_, _10802_);
  nor (_29059_, _29058_, _29003_);
  nor (_29060_, _29059_, _03589_);
  or (_29061_, _29060_, _08828_);
  or (_29062_, _29061_, _29056_);
  and (_29063_, _13347_, _05258_);
  or (_29064_, _29003_, _07766_);
  or (_29065_, _29064_, _29063_);
  and (_29066_, _13339_, _05258_);
  nor (_29067_, _29066_, _29003_);
  and (_29069_, _29067_, _03601_);
  nor (_29070_, _29069_, _03780_);
  and (_29071_, _29070_, _29065_);
  and (_29072_, _29071_, _29062_);
  and (_29073_, _13353_, _05258_);
  nor (_29074_, _29073_, _29003_);
  nor (_29075_, _29074_, _07778_);
  nor (_29076_, _29075_, _29072_);
  nor (_29077_, _29076_, _03622_);
  nor (_29078_, _29003_, _05412_);
  not (_29080_, _29078_);
  nor (_29081_, _29067_, _07777_);
  and (_29082_, _29081_, _29080_);
  nor (_29083_, _29082_, _29077_);
  nor (_29084_, _29083_, _03790_);
  nor (_29085_, _29008_, _06828_);
  and (_29086_, _29085_, _29080_);
  nor (_29087_, _29086_, _03624_);
  not (_29088_, _29087_);
  nor (_29089_, _29088_, _29084_);
  nor (_29091_, _13346_, _10802_);
  or (_29092_, _29003_, _07795_);
  nor (_29093_, _29092_, _29091_);
  or (_29094_, _29093_, _03785_);
  nor (_29095_, _29094_, _29089_);
  nor (_29096_, _13352_, _10802_);
  nor (_29097_, _29096_, _29003_);
  nor (_29098_, _29097_, _07793_);
  or (_29099_, _29098_, _29095_);
  and (_29100_, _29099_, _04246_);
  nor (_29102_, _29015_, _04246_);
  or (_29103_, _29102_, _29100_);
  and (_29104_, _29103_, _03823_);
  nor (_29105_, _29036_, _03823_);
  or (_29106_, _29105_, _29104_);
  and (_29107_, _29106_, _03514_);
  and (_29108_, _13402_, _05258_);
  nor (_29109_, _29108_, _29003_);
  nor (_29110_, _29109_, _03514_);
  or (_29111_, _29110_, _29107_);
  or (_29113_, _29111_, _43004_);
  or (_29114_, _43000_, \oc8051_golden_model_1.TCON [6]);
  and (_29115_, _29114_, _41806_);
  and (_43621_, _29115_, _29113_);
  not (_29116_, \oc8051_golden_model_1.TH0 [0]);
  nor (_29117_, _05263_, _29116_);
  nor (_29118_, _05666_, _10909_);
  nor (_29119_, _29118_, _29117_);
  and (_29120_, _29119_, _17166_);
  and (_29121_, _05263_, \oc8051_golden_model_1.ACC [0]);
  nor (_29123_, _29121_, _29117_);
  nor (_29124_, _29123_, _03737_);
  nor (_29125_, _29124_, _07390_);
  nor (_29126_, _29119_, _04081_);
  nor (_29127_, _04409_, _29116_);
  nor (_29128_, _29123_, _09029_);
  nor (_29129_, _29128_, _29127_);
  nor (_29130_, _29129_, _03610_);
  or (_29131_, _29130_, _03723_);
  nor (_29132_, _29131_, _29126_);
  or (_29134_, _29132_, _03729_);
  and (_29135_, _29134_, _29125_);
  and (_29136_, _05263_, _04620_);
  or (_29137_, _29117_, _25480_);
  nor (_29138_, _29137_, _29136_);
  nor (_29139_, _29138_, _29135_);
  nor (_29140_, _29139_, _04481_);
  and (_29141_, _06546_, _05263_);
  nor (_29142_, _29117_, _07400_);
  not (_29143_, _29142_);
  nor (_29145_, _29143_, _29141_);
  nor (_29146_, _29145_, _29140_);
  nor (_29147_, _29146_, _03222_);
  nor (_29148_, _12109_, _10909_);
  or (_29149_, _29117_, _03589_);
  nor (_29150_, _29149_, _29148_);
  or (_29151_, _29150_, _03601_);
  nor (_29152_, _29151_, _29147_);
  and (_29153_, _05263_, _06274_);
  nor (_29154_, _29153_, _29117_);
  nand (_29156_, _29154_, _07766_);
  and (_29157_, _29156_, _08828_);
  nor (_29158_, _29157_, _29152_);
  and (_29159_, _12124_, _05263_);
  nor (_29160_, _29159_, _29117_);
  and (_29161_, _29160_, _03600_);
  nor (_29162_, _29161_, _29158_);
  nor (_29163_, _29162_, _03780_);
  and (_29164_, _12128_, _05263_);
  or (_29165_, _29117_, _07778_);
  nor (_29167_, _29165_, _29164_);
  or (_29168_, _29167_, _03622_);
  nor (_29169_, _29168_, _29163_);
  or (_29170_, _29154_, _07777_);
  nor (_29171_, _29170_, _29118_);
  nor (_29172_, _29171_, _29169_);
  nor (_29173_, _29172_, _03790_);
  and (_29174_, _12005_, _05263_);
  or (_29175_, _29174_, _29117_);
  and (_29176_, _29175_, _03790_);
  or (_29178_, _29176_, _29173_);
  and (_29179_, _29178_, _07795_);
  nor (_29180_, _12122_, _10909_);
  nor (_29181_, _29180_, _29117_);
  nor (_29182_, _29181_, _07795_);
  or (_29183_, _29182_, _29179_);
  and (_29184_, _29183_, _07793_);
  nor (_29185_, _12003_, _10909_);
  nor (_29186_, _29185_, _29117_);
  nor (_29187_, _29186_, _07793_);
  nor (_29189_, _29187_, _17166_);
  not (_29190_, _29189_);
  nor (_29191_, _29190_, _29184_);
  nor (_29192_, _29191_, _29120_);
  or (_29193_, _29192_, _43004_);
  or (_29194_, _43000_, \oc8051_golden_model_1.TH0 [0]);
  and (_29195_, _29194_, _41806_);
  and (_43624_, _29195_, _29193_);
  and (_29196_, _06501_, _05263_);
  not (_29197_, \oc8051_golden_model_1.TH0 [1]);
  nor (_29199_, _05263_, _29197_);
  nor (_29200_, _29199_, _07400_);
  not (_29201_, _29200_);
  nor (_29202_, _29201_, _29196_);
  not (_29203_, _29202_);
  nor (_29204_, _05263_, \oc8051_golden_model_1.TH0 [1]);
  and (_29205_, _05263_, _03274_);
  nor (_29206_, _29205_, _29204_);
  and (_29207_, _29206_, _03729_);
  and (_29208_, _29206_, _04409_);
  nor (_29210_, _04409_, _29197_);
  or (_29211_, _29210_, _29208_);
  and (_29212_, _29211_, _04081_);
  and (_29213_, _12213_, _05263_);
  nor (_29214_, _29213_, _29204_);
  and (_29215_, _29214_, _03610_);
  or (_29216_, _29215_, _29212_);
  and (_29217_, _29216_, _03996_);
  and (_29218_, _05263_, _06764_);
  nor (_29219_, _29218_, _29199_);
  nor (_29221_, _29219_, _03996_);
  nor (_29222_, _29221_, _29217_);
  nor (_29223_, _29222_, _03729_);
  or (_29224_, _29223_, _07390_);
  nor (_29225_, _29224_, _29207_);
  and (_29226_, _29219_, _07390_);
  nor (_29227_, _29226_, _29225_);
  nor (_29228_, _29227_, _04481_);
  nor (_29229_, _29228_, _03222_);
  and (_29230_, _29229_, _29203_);
  not (_29232_, _29204_);
  and (_29233_, _12313_, _05263_);
  nor (_29234_, _29233_, _03589_);
  and (_29235_, _29234_, _29232_);
  nor (_29236_, _29235_, _29230_);
  nor (_29237_, _29236_, _08828_);
  nor (_29238_, _12327_, _10909_);
  nor (_29239_, _29238_, _07766_);
  and (_29240_, _05263_, _04303_);
  nor (_29241_, _29240_, _05886_);
  nor (_29243_, _29241_, _29239_);
  nor (_29244_, _29243_, _29204_);
  nor (_29245_, _29244_, _29237_);
  nor (_29246_, _29245_, _03780_);
  nor (_29247_, _12333_, _10909_);
  nor (_29248_, _29247_, _07778_);
  and (_29249_, _29248_, _29232_);
  nor (_29250_, _29249_, _29246_);
  nor (_29251_, _29250_, _03622_);
  nor (_29252_, _12207_, _10909_);
  nor (_29254_, _29252_, _07777_);
  and (_29255_, _29254_, _29232_);
  nor (_29256_, _29255_, _29251_);
  nor (_29257_, _29256_, _03790_);
  nor (_29258_, _29199_, _05618_);
  nor (_29259_, _29258_, _06828_);
  and (_29260_, _29259_, _29206_);
  nor (_29261_, _29260_, _29257_);
  or (_29262_, _29261_, _18499_);
  and (_29263_, _29240_, _05617_);
  nor (_29265_, _29263_, _07795_);
  and (_29266_, _29265_, _29232_);
  nand (_29267_, _29205_, _05617_);
  nor (_29268_, _29204_, _07793_);
  and (_29269_, _29268_, _29267_);
  or (_29270_, _29269_, _03815_);
  nor (_29271_, _29270_, _29266_);
  and (_29272_, _29271_, _29262_);
  nor (_29273_, _29214_, _04246_);
  nor (_29274_, _29273_, _29272_);
  and (_29276_, _29274_, _03514_);
  nor (_29277_, _29213_, _29199_);
  nor (_29278_, _29277_, _03514_);
  or (_29279_, _29278_, _29276_);
  or (_29280_, _29279_, _43004_);
  or (_29281_, _43000_, \oc8051_golden_model_1.TH0 [1]);
  and (_29282_, _29281_, _41806_);
  and (_43625_, _29282_, _29280_);
  not (_29283_, \oc8051_golden_model_1.TH0 [2]);
  nor (_29284_, _05263_, _29283_);
  nor (_29286_, _12538_, _10909_);
  nor (_29287_, _29286_, _29284_);
  nor (_29288_, _29287_, _07793_);
  nor (_29289_, _10909_, _04875_);
  nor (_29290_, _29289_, _29284_);
  and (_29291_, _29290_, _07390_);
  nor (_29292_, _12416_, _10909_);
  nor (_29293_, _29292_, _29284_);
  nor (_29294_, _29293_, _04081_);
  nor (_29295_, _04409_, _29283_);
  and (_29297_, _05263_, \oc8051_golden_model_1.ACC [2]);
  nor (_29298_, _29297_, _29284_);
  nor (_29299_, _29298_, _09029_);
  nor (_29300_, _29299_, _29295_);
  nor (_29301_, _29300_, _03610_);
  or (_29302_, _29301_, _29294_);
  and (_29303_, _29302_, _03996_);
  nor (_29304_, _29290_, _03996_);
  or (_29305_, _29304_, _29303_);
  and (_29306_, _29305_, _03737_);
  nor (_29308_, _29298_, _03737_);
  nor (_29309_, _29308_, _07390_);
  not (_29310_, _29309_);
  nor (_29311_, _29310_, _29306_);
  nor (_29312_, _29311_, _29291_);
  nor (_29313_, _29312_, _04481_);
  and (_29314_, _06637_, _05263_);
  nor (_29315_, _29284_, _07400_);
  not (_29316_, _29315_);
  nor (_29317_, _29316_, _29314_);
  nor (_29319_, _29317_, _29313_);
  nor (_29320_, _29319_, _03222_);
  nor (_29321_, _12519_, _10909_);
  or (_29322_, _29284_, _03589_);
  nor (_29323_, _29322_, _29321_);
  or (_29324_, _29323_, _03601_);
  nor (_29325_, _29324_, _29320_);
  and (_29326_, _05263_, _06332_);
  nor (_29327_, _29326_, _29284_);
  nand (_29328_, _29327_, _07766_);
  and (_29330_, _29328_, _08828_);
  nor (_29331_, _29330_, _29325_);
  and (_29332_, _12533_, _05263_);
  nor (_29333_, _29332_, _29284_);
  and (_29334_, _29333_, _03600_);
  nor (_29335_, _29334_, _29331_);
  nor (_29336_, _29335_, _03780_);
  and (_29337_, _12539_, _05263_);
  or (_29338_, _29284_, _07778_);
  nor (_29339_, _29338_, _29337_);
  or (_29341_, _29339_, _03622_);
  nor (_29342_, _29341_, _29336_);
  nor (_29343_, _29284_, _05718_);
  not (_29344_, _29343_);
  nor (_29345_, _29327_, _07777_);
  and (_29346_, _29345_, _29344_);
  nor (_29347_, _29346_, _29342_);
  nor (_29348_, _29347_, _03790_);
  nor (_29349_, _29298_, _06828_);
  and (_29350_, _29349_, _29344_);
  or (_29352_, _29350_, _29348_);
  and (_29353_, _29352_, _07795_);
  nor (_29354_, _12532_, _10909_);
  nor (_29355_, _29354_, _29284_);
  nor (_29356_, _29355_, _07795_);
  or (_29357_, _29356_, _29353_);
  and (_29358_, _29357_, _07793_);
  nor (_29359_, _29358_, _29288_);
  nor (_29360_, _29359_, _03815_);
  nor (_29361_, _29293_, _04246_);
  or (_29363_, _29361_, _03447_);
  nor (_29364_, _29363_, _29360_);
  and (_29365_, _12592_, _05263_);
  or (_29366_, _29284_, _03514_);
  nor (_29367_, _29366_, _29365_);
  nor (_29368_, _29367_, _29364_);
  or (_29369_, _29368_, _43004_);
  or (_29370_, _43000_, \oc8051_golden_model_1.TH0 [2]);
  and (_29371_, _29370_, _41806_);
  and (_43626_, _29371_, _29369_);
  not (_29373_, \oc8051_golden_model_1.TH0 [3]);
  nor (_29374_, _05263_, _29373_);
  nor (_29375_, _12738_, _10909_);
  nor (_29376_, _29375_, _29374_);
  nor (_29377_, _29376_, _07793_);
  and (_29378_, _12739_, _05263_);
  nor (_29379_, _29378_, _29374_);
  nor (_29380_, _29379_, _07778_);
  and (_29381_, _06592_, _05263_);
  or (_29382_, _29381_, _29374_);
  and (_29383_, _29382_, _04481_);
  and (_29384_, _05263_, \oc8051_golden_model_1.ACC [3]);
  nor (_29385_, _29384_, _29374_);
  nor (_29386_, _29385_, _03737_);
  nor (_29387_, _29385_, _09029_);
  nor (_29388_, _04409_, _29373_);
  or (_29389_, _29388_, _29387_);
  and (_29390_, _29389_, _04081_);
  nor (_29391_, _12627_, _10909_);
  nor (_29392_, _29391_, _29374_);
  nor (_29394_, _29392_, _04081_);
  or (_29395_, _29394_, _29390_);
  and (_29396_, _29395_, _03996_);
  nor (_29397_, _10909_, _05005_);
  nor (_29398_, _29397_, _29374_);
  nor (_29399_, _29398_, _03996_);
  nor (_29400_, _29399_, _29396_);
  nor (_29401_, _29400_, _03729_);
  or (_29402_, _29401_, _07390_);
  nor (_29403_, _29402_, _29386_);
  and (_29405_, _29398_, _07390_);
  or (_29406_, _29405_, _04481_);
  nor (_29407_, _29406_, _29403_);
  or (_29408_, _29407_, _29383_);
  and (_29409_, _29408_, _03589_);
  nor (_29410_, _12718_, _10909_);
  nor (_29411_, _29410_, _29374_);
  nor (_29412_, _29411_, _03589_);
  or (_29413_, _29412_, _08828_);
  or (_29414_, _29413_, _29409_);
  and (_29416_, _12733_, _05263_);
  or (_29417_, _29374_, _07766_);
  or (_29418_, _29417_, _29416_);
  and (_29419_, _05263_, _06276_);
  nor (_29420_, _29419_, _29374_);
  and (_29421_, _29420_, _03601_);
  nor (_29422_, _29421_, _03780_);
  and (_29423_, _29422_, _29418_);
  and (_29424_, _29423_, _29414_);
  nor (_29425_, _29424_, _29380_);
  nor (_29427_, _29425_, _03622_);
  nor (_29428_, _29374_, _05567_);
  not (_29429_, _29428_);
  nor (_29430_, _29420_, _07777_);
  and (_29431_, _29430_, _29429_);
  nor (_29432_, _29431_, _29427_);
  nor (_29433_, _29432_, _03790_);
  nor (_29434_, _29385_, _06828_);
  and (_29435_, _29434_, _29429_);
  nor (_29436_, _29435_, _03624_);
  not (_29438_, _29436_);
  nor (_29439_, _29438_, _29433_);
  nor (_29440_, _12732_, _10909_);
  or (_29441_, _29374_, _07795_);
  nor (_29442_, _29441_, _29440_);
  or (_29443_, _29442_, _03785_);
  nor (_29444_, _29443_, _29439_);
  nor (_29445_, _29444_, _29377_);
  nor (_29446_, _29445_, _03815_);
  nor (_29447_, _29392_, _04246_);
  or (_29449_, _29447_, _03447_);
  nor (_29450_, _29449_, _29446_);
  and (_29451_, _12794_, _05263_);
  or (_29452_, _29374_, _03514_);
  nor (_29453_, _29452_, _29451_);
  nor (_29454_, _29453_, _29450_);
  or (_29455_, _29454_, _43004_);
  or (_29456_, _43000_, \oc8051_golden_model_1.TH0 [3]);
  and (_29457_, _29456_, _41806_);
  and (_43627_, _29457_, _29455_);
  not (_29459_, \oc8051_golden_model_1.TH0 [4]);
  nor (_29460_, _05263_, _29459_);
  nor (_29461_, _12816_, _10909_);
  nor (_29462_, _29461_, _29460_);
  nor (_29463_, _29462_, _07793_);
  and (_29464_, _12817_, _05263_);
  nor (_29465_, _29464_, _29460_);
  nor (_29466_, _29465_, _07778_);
  and (_29467_, _06298_, _05263_);
  nor (_29468_, _29467_, _29460_);
  and (_29470_, _29468_, _03601_);
  and (_29471_, _05263_, \oc8051_golden_model_1.ACC [4]);
  nor (_29472_, _29471_, _29460_);
  nor (_29473_, _29472_, _03737_);
  nor (_29474_, _29472_, _09029_);
  nor (_29475_, _04409_, _29459_);
  or (_29476_, _29475_, _29474_);
  and (_29477_, _29476_, _04081_);
  nor (_29478_, _12841_, _10909_);
  nor (_29479_, _29478_, _29460_);
  nor (_29481_, _29479_, _04081_);
  or (_29482_, _29481_, _29477_);
  and (_29483_, _29482_, _03996_);
  nor (_29484_, _05777_, _10909_);
  nor (_29485_, _29484_, _29460_);
  nor (_29486_, _29485_, _03996_);
  nor (_29487_, _29486_, _29483_);
  nor (_29488_, _29487_, _03729_);
  or (_29489_, _29488_, _07390_);
  nor (_29490_, _29489_, _29473_);
  and (_29492_, _29485_, _07390_);
  nor (_29493_, _29492_, _29490_);
  nor (_29494_, _29493_, _04481_);
  and (_29495_, _06730_, _05263_);
  nor (_29496_, _29460_, _07400_);
  not (_29497_, _29496_);
  nor (_29498_, _29497_, _29495_);
  or (_29499_, _29498_, _03222_);
  nor (_29500_, _29499_, _29494_);
  nor (_29501_, _12933_, _10909_);
  nor (_29502_, _29501_, _29460_);
  nor (_29503_, _29502_, _03589_);
  or (_29504_, _29503_, _03601_);
  nor (_29505_, _29504_, _29500_);
  nor (_29506_, _29505_, _29470_);
  or (_29507_, _29506_, _03600_);
  and (_29508_, _12821_, _05263_);
  or (_29509_, _29508_, _29460_);
  or (_29510_, _29509_, _07766_);
  and (_29511_, _29510_, _07778_);
  and (_29514_, _29511_, _29507_);
  nor (_29515_, _29514_, _29466_);
  nor (_29516_, _29515_, _03622_);
  nor (_29517_, _29460_, _05825_);
  not (_29518_, _29517_);
  nor (_29519_, _29468_, _07777_);
  and (_29520_, _29519_, _29518_);
  nor (_29521_, _29520_, _29516_);
  nor (_29522_, _29521_, _03790_);
  nor (_29523_, _29472_, _06828_);
  and (_29525_, _29523_, _29518_);
  nor (_29526_, _29525_, _03624_);
  not (_29527_, _29526_);
  nor (_29528_, _29527_, _29522_);
  nor (_29529_, _12819_, _10909_);
  or (_29530_, _29460_, _07795_);
  nor (_29531_, _29530_, _29529_);
  or (_29532_, _29531_, _03785_);
  nor (_29533_, _29532_, _29528_);
  nor (_29534_, _29533_, _29463_);
  nor (_29536_, _29534_, _03815_);
  nor (_29537_, _29479_, _04246_);
  or (_29538_, _29537_, _03447_);
  nor (_29539_, _29538_, _29536_);
  and (_29540_, _13003_, _05263_);
  or (_29541_, _29460_, _03514_);
  nor (_29542_, _29541_, _29540_);
  nor (_29543_, _29542_, _29539_);
  or (_29544_, _29543_, _43004_);
  or (_29545_, _43000_, \oc8051_golden_model_1.TH0 [4]);
  and (_29547_, _29545_, _41806_);
  and (_43628_, _29547_, _29544_);
  not (_29548_, \oc8051_golden_model_1.TH0 [5]);
  nor (_29549_, _05263_, _29548_);
  nor (_29550_, _13146_, _10909_);
  nor (_29551_, _29550_, _29549_);
  nor (_29552_, _29551_, _07793_);
  and (_29553_, _13147_, _05263_);
  nor (_29554_, _29553_, _29549_);
  nor (_29555_, _29554_, _07778_);
  and (_29557_, _06684_, _05263_);
  or (_29558_, _29557_, _29549_);
  and (_29559_, _29558_, _04481_);
  and (_29560_, _05263_, \oc8051_golden_model_1.ACC [5]);
  nor (_29561_, _29560_, _29549_);
  nor (_29562_, _29561_, _03737_);
  nor (_29563_, _29561_, _09029_);
  nor (_29564_, _04409_, _29548_);
  or (_29565_, _29564_, _29563_);
  and (_29566_, _29565_, _04081_);
  nor (_29568_, _13014_, _10909_);
  nor (_29569_, _29568_, _29549_);
  nor (_29570_, _29569_, _04081_);
  or (_29571_, _29570_, _29566_);
  and (_29572_, _29571_, _03996_);
  nor (_29573_, _05469_, _10909_);
  nor (_29574_, _29573_, _29549_);
  nor (_29575_, _29574_, _03996_);
  nor (_29576_, _29575_, _29572_);
  nor (_29577_, _29576_, _03729_);
  or (_29579_, _29577_, _07390_);
  nor (_29580_, _29579_, _29562_);
  and (_29581_, _29574_, _07390_);
  or (_29582_, _29581_, _04481_);
  nor (_29583_, _29582_, _29580_);
  or (_29584_, _29583_, _29559_);
  and (_29585_, _29584_, _03589_);
  nor (_29586_, _13127_, _10909_);
  nor (_29587_, _29586_, _29549_);
  nor (_29588_, _29587_, _03589_);
  or (_29590_, _29588_, _08828_);
  or (_29591_, _29590_, _29585_);
  and (_29592_, _13141_, _05263_);
  or (_29593_, _29549_, _07766_);
  or (_29594_, _29593_, _29592_);
  and (_29595_, _06306_, _05263_);
  nor (_29596_, _29595_, _29549_);
  and (_29597_, _29596_, _03601_);
  nor (_29598_, _29597_, _03780_);
  and (_29599_, _29598_, _29594_);
  and (_29601_, _29599_, _29591_);
  nor (_29602_, _29601_, _29555_);
  nor (_29603_, _29602_, _03622_);
  nor (_29604_, _29549_, _05518_);
  not (_29605_, _29604_);
  nor (_29606_, _29596_, _07777_);
  and (_29607_, _29606_, _29605_);
  nor (_29608_, _29607_, _29603_);
  nor (_29609_, _29608_, _03790_);
  nor (_29610_, _29561_, _06828_);
  and (_29612_, _29610_, _29605_);
  or (_29613_, _29612_, _29609_);
  and (_29614_, _29613_, _07795_);
  nor (_29615_, _13140_, _10909_);
  nor (_29616_, _29615_, _29549_);
  nor (_29617_, _29616_, _07795_);
  or (_29618_, _29617_, _29614_);
  and (_29619_, _29618_, _07793_);
  nor (_29620_, _29619_, _29552_);
  nor (_29621_, _29620_, _03815_);
  nor (_29623_, _29569_, _04246_);
  or (_29624_, _29623_, _03447_);
  nor (_29625_, _29624_, _29621_);
  and (_29626_, _13199_, _05263_);
  or (_29627_, _29549_, _03514_);
  nor (_29628_, _29627_, _29626_);
  nor (_29629_, _29628_, _29625_);
  or (_29630_, _29629_, _43004_);
  or (_29631_, _43000_, \oc8051_golden_model_1.TH0 [5]);
  and (_29632_, _29631_, _41806_);
  and (_43629_, _29632_, _29630_);
  not (_29634_, \oc8051_golden_model_1.TH0 [6]);
  nor (_29635_, _05263_, _29634_);
  nor (_29636_, _13352_, _10909_);
  nor (_29637_, _29636_, _29635_);
  nor (_29638_, _29637_, _07793_);
  and (_29639_, _13353_, _05263_);
  nor (_29640_, _29639_, _29635_);
  nor (_29641_, _29640_, _07778_);
  and (_29642_, _06455_, _05263_);
  or (_29644_, _29642_, _29635_);
  and (_29645_, _29644_, _04481_);
  and (_29646_, _05263_, \oc8051_golden_model_1.ACC [6]);
  nor (_29647_, _29646_, _29635_);
  nor (_29648_, _29647_, _03737_);
  nor (_29649_, _29647_, _09029_);
  nor (_29650_, _04409_, _29634_);
  or (_29651_, _29650_, _29649_);
  and (_29652_, _29651_, _04081_);
  nor (_29653_, _13242_, _10909_);
  nor (_29655_, _29653_, _29635_);
  nor (_29656_, _29655_, _04081_);
  or (_29657_, _29656_, _29652_);
  and (_29658_, _29657_, _03996_);
  nor (_29659_, _05363_, _10909_);
  nor (_29660_, _29659_, _29635_);
  nor (_29661_, _29660_, _03996_);
  nor (_29662_, _29661_, _29658_);
  nor (_29663_, _29662_, _03729_);
  or (_29664_, _29663_, _07390_);
  nor (_29666_, _29664_, _29648_);
  and (_29667_, _29660_, _07390_);
  or (_29668_, _29667_, _04481_);
  nor (_29669_, _29668_, _29666_);
  or (_29670_, _29669_, _29645_);
  and (_29671_, _29670_, _03589_);
  nor (_29672_, _13332_, _10909_);
  nor (_29673_, _29672_, _29635_);
  nor (_29674_, _29673_, _03589_);
  or (_29675_, _29674_, _08828_);
  or (_29677_, _29675_, _29671_);
  and (_29678_, _13347_, _05263_);
  or (_29679_, _29635_, _07766_);
  or (_29680_, _29679_, _29678_);
  and (_29681_, _13339_, _05263_);
  nor (_29682_, _29681_, _29635_);
  and (_29683_, _29682_, _03601_);
  nor (_29684_, _29683_, _03780_);
  and (_29685_, _29684_, _29680_);
  and (_29686_, _29685_, _29677_);
  nor (_29688_, _29686_, _29641_);
  nor (_29689_, _29688_, _03622_);
  nor (_29690_, _29635_, _05412_);
  not (_29691_, _29690_);
  nor (_29692_, _29682_, _07777_);
  and (_29693_, _29692_, _29691_);
  nor (_29694_, _29693_, _29689_);
  nor (_29695_, _29694_, _03790_);
  nor (_29696_, _29647_, _06828_);
  and (_29697_, _29696_, _29691_);
  nor (_29699_, _29697_, _03624_);
  not (_29700_, _29699_);
  nor (_29701_, _29700_, _29695_);
  nor (_29702_, _13346_, _10909_);
  or (_29703_, _29635_, _07795_);
  nor (_29704_, _29703_, _29702_);
  or (_29705_, _29704_, _03785_);
  nor (_29706_, _29705_, _29701_);
  nor (_29707_, _29706_, _29638_);
  nor (_29708_, _29707_, _03815_);
  nor (_29710_, _29655_, _04246_);
  or (_29711_, _29710_, _03447_);
  nor (_29712_, _29711_, _29708_);
  and (_29713_, _13402_, _05263_);
  or (_29714_, _29635_, _03514_);
  nor (_29715_, _29714_, _29713_);
  nor (_29716_, _29715_, _29712_);
  or (_29717_, _29716_, _43004_);
  or (_29718_, _43000_, \oc8051_golden_model_1.TH0 [6]);
  and (_29719_, _29718_, _41806_);
  and (_43630_, _29719_, _29717_);
  not (_29721_, \oc8051_golden_model_1.TH1 [0]);
  nor (_29722_, _05278_, _29721_);
  nor (_29723_, _05666_, _10991_);
  nor (_29724_, _29723_, _29722_);
  and (_29725_, _29724_, _17166_);
  and (_29726_, _05278_, \oc8051_golden_model_1.ACC [0]);
  nor (_29727_, _29726_, _29722_);
  nor (_29728_, _29727_, _03737_);
  nor (_29729_, _29727_, _09029_);
  nor (_29731_, _04409_, _29721_);
  or (_29732_, _29731_, _29729_);
  and (_29733_, _29732_, _04081_);
  nor (_29734_, _29724_, _04081_);
  or (_29735_, _29734_, _29733_);
  and (_29736_, _29735_, _03996_);
  and (_29737_, _05278_, _04620_);
  nor (_29738_, _29737_, _29722_);
  nor (_29739_, _29738_, _03996_);
  nor (_29740_, _29739_, _29736_);
  nor (_29742_, _29740_, _03729_);
  or (_29743_, _29742_, _07390_);
  nor (_29744_, _29743_, _29728_);
  and (_29745_, _29738_, _07390_);
  nor (_29746_, _29745_, _29744_);
  nor (_29747_, _29746_, _04481_);
  and (_29748_, _06546_, _05278_);
  nor (_29749_, _29722_, _07400_);
  not (_29750_, _29749_);
  nor (_29751_, _29750_, _29748_);
  nor (_29753_, _29751_, _29747_);
  nor (_29754_, _29753_, _03222_);
  nor (_29755_, _12109_, _10991_);
  or (_29756_, _29722_, _03589_);
  nor (_29757_, _29756_, _29755_);
  or (_29758_, _29757_, _03601_);
  nor (_29759_, _29758_, _29754_);
  and (_29760_, _05278_, _06274_);
  nor (_29761_, _29760_, _29722_);
  nand (_29762_, _29761_, _07766_);
  and (_29763_, _29762_, _08828_);
  nor (_29764_, _29763_, _29759_);
  and (_29765_, _12124_, _05278_);
  nor (_29766_, _29765_, _29722_);
  and (_29767_, _29766_, _03600_);
  nor (_29768_, _29767_, _29764_);
  nor (_29769_, _29768_, _03780_);
  and (_29770_, _12128_, _05278_);
  or (_29771_, _29722_, _07778_);
  nor (_29772_, _29771_, _29770_);
  or (_29775_, _29772_, _03622_);
  nor (_29776_, _29775_, _29769_);
  or (_29777_, _29761_, _07777_);
  nor (_29778_, _29777_, _29723_);
  nor (_29779_, _29778_, _29776_);
  nor (_29780_, _29779_, _03790_);
  nor (_29781_, _29722_, _05666_);
  or (_29782_, _29781_, _06828_);
  nor (_29783_, _29782_, _29727_);
  or (_29784_, _29783_, _29780_);
  and (_29786_, _29784_, _07795_);
  nor (_29787_, _12122_, _10991_);
  nor (_29788_, _29787_, _29722_);
  nor (_29789_, _29788_, _07795_);
  or (_29790_, _29789_, _29786_);
  and (_29791_, _29790_, _07793_);
  nor (_29792_, _12003_, _10991_);
  nor (_29793_, _29792_, _29722_);
  nor (_29794_, _29793_, _07793_);
  nor (_29795_, _29794_, _17166_);
  not (_29797_, _29795_);
  nor (_29798_, _29797_, _29791_);
  nor (_29799_, _29798_, _29725_);
  or (_29800_, _29799_, _43004_);
  or (_29801_, _43000_, \oc8051_golden_model_1.TH1 [0]);
  and (_29802_, _29801_, _41806_);
  and (_43631_, _29802_, _29800_);
  and (_29803_, _06501_, _05278_);
  not (_29804_, \oc8051_golden_model_1.TH1 [1]);
  nor (_29805_, _05278_, _29804_);
  nor (_29807_, _29805_, _07400_);
  not (_29808_, _29807_);
  nor (_29809_, _29808_, _29803_);
  not (_29810_, _29809_);
  and (_29811_, _05278_, _06764_);
  or (_29812_, _29805_, _25480_);
  nor (_29813_, _29812_, _29811_);
  nor (_29814_, _05278_, \oc8051_golden_model_1.TH1 [1]);
  and (_29815_, _05278_, _03274_);
  nor (_29816_, _29815_, _29814_);
  and (_29818_, _29816_, _03729_);
  nor (_29819_, _29818_, _07390_);
  and (_29820_, _12213_, _05278_);
  nor (_29821_, _29820_, _29814_);
  and (_29822_, _29821_, _03610_);
  and (_29823_, _29816_, _04409_);
  nor (_29824_, _04409_, _29804_);
  nor (_29825_, _29824_, _29823_);
  nor (_29826_, _29825_, _03610_);
  or (_29827_, _29826_, _03723_);
  nor (_29829_, _29827_, _29822_);
  or (_29830_, _29829_, _03729_);
  and (_29831_, _29830_, _29819_);
  nor (_29832_, _29831_, _29813_);
  nor (_29833_, _29832_, _04481_);
  nor (_29834_, _29833_, _03222_);
  and (_29835_, _29834_, _29810_);
  not (_29836_, _29814_);
  and (_29837_, _12313_, _05278_);
  nor (_29838_, _29837_, _03589_);
  and (_29840_, _29838_, _29836_);
  nor (_29841_, _29840_, _29835_);
  nor (_29842_, _29841_, _08828_);
  nor (_29843_, _12327_, _10991_);
  nor (_29844_, _29843_, _07766_);
  and (_29845_, _05278_, _04303_);
  nor (_29846_, _29845_, _05886_);
  nor (_29847_, _29846_, _29844_);
  nor (_29848_, _29847_, _29814_);
  nor (_29849_, _29848_, _29842_);
  nor (_29851_, _29849_, _03780_);
  nor (_29852_, _12333_, _10991_);
  nor (_29853_, _29852_, _07778_);
  and (_29854_, _29853_, _29836_);
  nor (_29855_, _29854_, _29851_);
  nor (_29856_, _29855_, _03622_);
  nor (_29857_, _12207_, _10991_);
  nor (_29858_, _29857_, _07777_);
  and (_29859_, _29858_, _29836_);
  nor (_29860_, _29859_, _29856_);
  nor (_29862_, _29860_, _03790_);
  nor (_29863_, _29805_, _05618_);
  nor (_29864_, _29863_, _06828_);
  and (_29865_, _29864_, _29816_);
  nor (_29866_, _29865_, _29862_);
  or (_29867_, _29866_, _18499_);
  nand (_29868_, _29815_, _05617_);
  nor (_29869_, _29814_, _07793_);
  and (_29870_, _29869_, _29868_);
  nor (_29871_, _29870_, _03815_);
  and (_29873_, _29845_, _05617_);
  or (_29874_, _29814_, _07795_);
  or (_29875_, _29874_, _29873_);
  and (_29876_, _29875_, _29871_);
  and (_29877_, _29876_, _29867_);
  nor (_29878_, _29821_, _04246_);
  nor (_29879_, _29878_, _29877_);
  and (_29880_, _29879_, _03514_);
  nor (_29881_, _29820_, _29805_);
  nor (_29882_, _29881_, _03514_);
  or (_29884_, _29882_, _29880_);
  or (_29885_, _29884_, _43004_);
  or (_29886_, _43000_, \oc8051_golden_model_1.TH1 [1]);
  and (_29887_, _29886_, _41806_);
  and (_43632_, _29887_, _29885_);
  not (_29888_, \oc8051_golden_model_1.TH1 [2]);
  nor (_29889_, _05278_, _29888_);
  nor (_29890_, _12538_, _10991_);
  nor (_29891_, _29890_, _29889_);
  nor (_29892_, _29891_, _07793_);
  and (_29894_, _12539_, _05278_);
  nor (_29895_, _29894_, _29889_);
  nor (_29896_, _29895_, _07778_);
  and (_29897_, _05278_, \oc8051_golden_model_1.ACC [2]);
  nor (_29898_, _29897_, _29889_);
  nor (_29899_, _29898_, _03737_);
  nor (_29900_, _29898_, _09029_);
  nor (_29901_, _04409_, _29888_);
  or (_29902_, _29901_, _29900_);
  and (_29903_, _29902_, _04081_);
  nor (_29905_, _12416_, _10991_);
  nor (_29906_, _29905_, _29889_);
  nor (_29907_, _29906_, _04081_);
  or (_29908_, _29907_, _29903_);
  and (_29909_, _29908_, _03996_);
  nor (_29910_, _10991_, _04875_);
  nor (_29911_, _29910_, _29889_);
  nor (_29912_, _29911_, _03996_);
  nor (_29913_, _29912_, _29909_);
  nor (_29914_, _29913_, _03729_);
  or (_29916_, _29914_, _07390_);
  nor (_29917_, _29916_, _29899_);
  and (_29918_, _29911_, _07390_);
  nor (_29919_, _29918_, _29917_);
  nor (_29920_, _29919_, _04481_);
  and (_29921_, _06637_, _05278_);
  nor (_29922_, _29889_, _07400_);
  not (_29923_, _29922_);
  nor (_29924_, _29923_, _29921_);
  nor (_29925_, _29924_, _03222_);
  not (_29927_, _29925_);
  nor (_29928_, _29927_, _29920_);
  nor (_29929_, _12519_, _10991_);
  nor (_29930_, _29929_, _29889_);
  nor (_29931_, _29930_, _03589_);
  or (_29932_, _29931_, _08828_);
  or (_29933_, _29932_, _29928_);
  and (_29934_, _12533_, _05278_);
  or (_29935_, _29889_, _07766_);
  or (_29936_, _29935_, _29934_);
  and (_29938_, _05278_, _06332_);
  nor (_29939_, _29938_, _29889_);
  and (_29940_, _29939_, _03601_);
  nor (_29941_, _29940_, _03780_);
  and (_29942_, _29941_, _29936_);
  and (_29943_, _29942_, _29933_);
  nor (_29944_, _29943_, _29896_);
  nor (_29945_, _29944_, _03622_);
  nor (_29946_, _29889_, _05718_);
  not (_29947_, _29946_);
  nor (_29949_, _29939_, _07777_);
  and (_29950_, _29949_, _29947_);
  nor (_29951_, _29950_, _29945_);
  nor (_29952_, _29951_, _03790_);
  nor (_29953_, _29898_, _06828_);
  and (_29954_, _29953_, _29947_);
  or (_29955_, _29954_, _29952_);
  and (_29956_, _29955_, _07795_);
  nor (_29957_, _12532_, _10991_);
  nor (_29958_, _29957_, _29889_);
  nor (_29960_, _29958_, _07795_);
  or (_29961_, _29960_, _29956_);
  and (_29962_, _29961_, _07793_);
  nor (_29963_, _29962_, _29892_);
  nor (_29964_, _29963_, _03815_);
  nor (_29965_, _29906_, _04246_);
  or (_29966_, _29965_, _03447_);
  nor (_29967_, _29966_, _29964_);
  and (_29968_, _12592_, _05278_);
  or (_29969_, _29889_, _03514_);
  nor (_29971_, _29969_, _29968_);
  nor (_29972_, _29971_, _29967_);
  or (_29973_, _29972_, _43004_);
  or (_29974_, _43000_, \oc8051_golden_model_1.TH1 [2]);
  and (_29975_, _29974_, _41806_);
  and (_43633_, _29975_, _29973_);
  not (_29976_, \oc8051_golden_model_1.TH1 [3]);
  nor (_29977_, _05278_, _29976_);
  nor (_29978_, _12738_, _10991_);
  nor (_29979_, _29978_, _29977_);
  nor (_29981_, _29979_, _07793_);
  and (_29982_, _12739_, _05278_);
  nor (_29983_, _29982_, _29977_);
  nor (_29984_, _29983_, _07778_);
  and (_29985_, _06592_, _05278_);
  or (_29986_, _29985_, _29977_);
  and (_29987_, _29986_, _04481_);
  and (_29988_, _05278_, \oc8051_golden_model_1.ACC [3]);
  nor (_29989_, _29988_, _29977_);
  nor (_29990_, _29989_, _03737_);
  nor (_29992_, _29989_, _09029_);
  nor (_29993_, _04409_, _29976_);
  or (_29994_, _29993_, _29992_);
  and (_29995_, _29994_, _04081_);
  nor (_29996_, _12627_, _10991_);
  nor (_29997_, _29996_, _29977_);
  nor (_29998_, _29997_, _04081_);
  or (_29999_, _29998_, _29995_);
  and (_30000_, _29999_, _03996_);
  nor (_30001_, _10991_, _05005_);
  nor (_30003_, _30001_, _29977_);
  nor (_30004_, _30003_, _03996_);
  nor (_30005_, _30004_, _30000_);
  nor (_30006_, _30005_, _03729_);
  or (_30007_, _30006_, _07390_);
  nor (_30008_, _30007_, _29990_);
  and (_30009_, _30003_, _07390_);
  or (_30010_, _30009_, _04481_);
  nor (_30011_, _30010_, _30008_);
  or (_30012_, _30011_, _29987_);
  and (_30014_, _30012_, _03589_);
  nor (_30015_, _12718_, _10991_);
  nor (_30016_, _30015_, _29977_);
  nor (_30017_, _30016_, _03589_);
  or (_30018_, _30017_, _08828_);
  or (_30019_, _30018_, _30014_);
  and (_30020_, _12733_, _05278_);
  or (_30021_, _29977_, _07766_);
  or (_30022_, _30021_, _30020_);
  and (_30023_, _05278_, _06276_);
  nor (_30025_, _30023_, _29977_);
  and (_30026_, _30025_, _03601_);
  nor (_30027_, _30026_, _03780_);
  and (_30028_, _30027_, _30022_);
  and (_30029_, _30028_, _30019_);
  nor (_30030_, _30029_, _29984_);
  nor (_30031_, _30030_, _03622_);
  nor (_30032_, _29977_, _05567_);
  not (_30033_, _30032_);
  nor (_30034_, _30025_, _07777_);
  and (_30036_, _30034_, _30033_);
  nor (_30037_, _30036_, _30031_);
  nor (_30038_, _30037_, _03790_);
  nor (_30039_, _29989_, _06828_);
  and (_30040_, _30039_, _30033_);
  or (_30041_, _30040_, _30038_);
  and (_30042_, _30041_, _07795_);
  nor (_30043_, _12732_, _10991_);
  nor (_30044_, _30043_, _29977_);
  nor (_30045_, _30044_, _07795_);
  or (_30047_, _30045_, _30042_);
  and (_30048_, _30047_, _07793_);
  nor (_30049_, _30048_, _29981_);
  nor (_30050_, _30049_, _03815_);
  nor (_30051_, _29997_, _04246_);
  or (_30052_, _30051_, _03447_);
  nor (_30053_, _30052_, _30050_);
  and (_30054_, _12794_, _05278_);
  or (_30055_, _29977_, _03514_);
  nor (_30056_, _30055_, _30054_);
  nor (_30058_, _30056_, _30053_);
  or (_30059_, _30058_, _43004_);
  or (_30060_, _43000_, \oc8051_golden_model_1.TH1 [3]);
  and (_30061_, _30060_, _41806_);
  and (_43634_, _30061_, _30059_);
  not (_30062_, \oc8051_golden_model_1.TH1 [4]);
  nor (_30063_, _05278_, _30062_);
  nor (_30064_, _12816_, _10991_);
  nor (_30065_, _30064_, _30063_);
  nor (_30066_, _30065_, _07793_);
  and (_30067_, _12817_, _05278_);
  nor (_30068_, _30067_, _30063_);
  nor (_30069_, _30068_, _07778_);
  and (_30070_, _06298_, _05278_);
  nor (_30071_, _30070_, _30063_);
  and (_30072_, _30071_, _03601_);
  nor (_30073_, _05777_, _10991_);
  nor (_30074_, _30073_, _30063_);
  and (_30075_, _30074_, _07390_);
  and (_30076_, _05278_, \oc8051_golden_model_1.ACC [4]);
  nor (_30079_, _30076_, _30063_);
  nor (_30080_, _30079_, _03737_);
  nor (_30081_, _30079_, _09029_);
  nor (_30082_, _04409_, _30062_);
  or (_30083_, _30082_, _30081_);
  and (_30084_, _30083_, _04081_);
  nor (_30085_, _12841_, _10991_);
  nor (_30086_, _30085_, _30063_);
  nor (_30087_, _30086_, _04081_);
  or (_30088_, _30087_, _30084_);
  and (_30089_, _30088_, _03996_);
  nor (_30090_, _30074_, _03996_);
  nor (_30091_, _30090_, _30089_);
  nor (_30092_, _30091_, _03729_);
  or (_30093_, _30092_, _07390_);
  nor (_30094_, _30093_, _30080_);
  nor (_30095_, _30094_, _30075_);
  nor (_30096_, _30095_, _04481_);
  and (_30097_, _06730_, _05278_);
  nor (_30098_, _30063_, _07400_);
  not (_30100_, _30098_);
  nor (_30101_, _30100_, _30097_);
  or (_30102_, _30101_, _03222_);
  nor (_30103_, _30102_, _30096_);
  nor (_30104_, _12933_, _10991_);
  nor (_30105_, _30104_, _30063_);
  nor (_30106_, _30105_, _03589_);
  or (_30107_, _30106_, _03601_);
  nor (_30108_, _30107_, _30103_);
  nor (_30109_, _30108_, _30072_);
  or (_30111_, _30109_, _03600_);
  and (_30112_, _12821_, _05278_);
  or (_30113_, _30112_, _30063_);
  or (_30114_, _30113_, _07766_);
  and (_30115_, _30114_, _07778_);
  and (_30116_, _30115_, _30111_);
  nor (_30117_, _30116_, _30069_);
  nor (_30118_, _30117_, _03622_);
  nor (_30119_, _30063_, _05825_);
  not (_30120_, _30119_);
  nor (_30122_, _30071_, _07777_);
  and (_30123_, _30122_, _30120_);
  nor (_30124_, _30123_, _30118_);
  nor (_30125_, _30124_, _03790_);
  nor (_30126_, _30079_, _06828_);
  and (_30127_, _30126_, _30120_);
  nor (_30128_, _30127_, _03624_);
  not (_30129_, _30128_);
  nor (_30130_, _30129_, _30125_);
  nor (_30131_, _12819_, _10991_);
  or (_30133_, _30063_, _07795_);
  nor (_30134_, _30133_, _30131_);
  or (_30135_, _30134_, _03785_);
  nor (_30136_, _30135_, _30130_);
  nor (_30137_, _30136_, _30066_);
  nor (_30138_, _30137_, _03815_);
  nor (_30139_, _30086_, _04246_);
  or (_30140_, _30139_, _03447_);
  nor (_30141_, _30140_, _30138_);
  and (_30142_, _13003_, _05278_);
  or (_30144_, _30063_, _03514_);
  nor (_30145_, _30144_, _30142_);
  nor (_30146_, _30145_, _30141_);
  or (_30147_, _30146_, _43004_);
  or (_30148_, _43000_, \oc8051_golden_model_1.TH1 [4]);
  and (_30149_, _30148_, _41806_);
  and (_43635_, _30149_, _30147_);
  not (_30150_, \oc8051_golden_model_1.TH1 [5]);
  nor (_30151_, _05278_, _30150_);
  nor (_30152_, _13146_, _10991_);
  nor (_30154_, _30152_, _30151_);
  nor (_30155_, _30154_, _07793_);
  and (_30156_, _13147_, _05278_);
  nor (_30157_, _30156_, _30151_);
  nor (_30158_, _30157_, _07778_);
  and (_30159_, _06684_, _05278_);
  or (_30160_, _30159_, _30151_);
  and (_30161_, _30160_, _04481_);
  and (_30162_, _05278_, \oc8051_golden_model_1.ACC [5]);
  nor (_30163_, _30162_, _30151_);
  nor (_30165_, _30163_, _03737_);
  nor (_30166_, _30163_, _09029_);
  nor (_30167_, _04409_, _30150_);
  or (_30168_, _30167_, _30166_);
  and (_30169_, _30168_, _04081_);
  nor (_30170_, _13014_, _10991_);
  nor (_30171_, _30170_, _30151_);
  nor (_30172_, _30171_, _04081_);
  or (_30173_, _30172_, _30169_);
  and (_30174_, _30173_, _03996_);
  nor (_30176_, _05469_, _10991_);
  nor (_30177_, _30176_, _30151_);
  nor (_30178_, _30177_, _03996_);
  nor (_30179_, _30178_, _30174_);
  nor (_30180_, _30179_, _03729_);
  or (_30181_, _30180_, _07390_);
  nor (_30182_, _30181_, _30165_);
  and (_30183_, _30177_, _07390_);
  or (_30184_, _30183_, _04481_);
  nor (_30185_, _30184_, _30182_);
  or (_30187_, _30185_, _30161_);
  and (_30188_, _30187_, _03589_);
  nor (_30189_, _13127_, _10991_);
  nor (_30190_, _30189_, _30151_);
  nor (_30191_, _30190_, _03589_);
  or (_30192_, _30191_, _08828_);
  or (_30193_, _30192_, _30188_);
  and (_30194_, _13141_, _05278_);
  or (_30195_, _30151_, _07766_);
  or (_30196_, _30195_, _30194_);
  and (_30198_, _06306_, _05278_);
  nor (_30199_, _30198_, _30151_);
  and (_30200_, _30199_, _03601_);
  nor (_30201_, _30200_, _03780_);
  and (_30202_, _30201_, _30196_);
  and (_30203_, _30202_, _30193_);
  nor (_30204_, _30203_, _30158_);
  nor (_30205_, _30204_, _03622_);
  nor (_30206_, _30151_, _05518_);
  not (_30207_, _30206_);
  nor (_30209_, _30199_, _07777_);
  and (_30210_, _30209_, _30207_);
  nor (_30211_, _30210_, _30205_);
  nor (_30212_, _30211_, _03790_);
  nor (_30213_, _30163_, _06828_);
  and (_30214_, _30213_, _30207_);
  nor (_30215_, _30214_, _03624_);
  not (_30216_, _30215_);
  nor (_30217_, _30216_, _30212_);
  nor (_30218_, _13140_, _10991_);
  or (_30220_, _30151_, _07795_);
  nor (_30221_, _30220_, _30218_);
  or (_30222_, _30221_, _03785_);
  nor (_30223_, _30222_, _30217_);
  nor (_30224_, _30223_, _30155_);
  nor (_30225_, _30224_, _03815_);
  nor (_30226_, _30171_, _04246_);
  or (_30227_, _30226_, _03447_);
  nor (_30228_, _30227_, _30225_);
  and (_30229_, _13199_, _05278_);
  or (_30231_, _30151_, _03514_);
  nor (_30232_, _30231_, _30229_);
  nor (_30233_, _30232_, _30228_);
  or (_30234_, _30233_, _43004_);
  or (_30235_, _43000_, \oc8051_golden_model_1.TH1 [5]);
  and (_30236_, _30235_, _41806_);
  and (_43638_, _30236_, _30234_);
  not (_30237_, \oc8051_golden_model_1.TH1 [6]);
  nor (_30238_, _05278_, _30237_);
  nor (_30239_, _13352_, _10991_);
  nor (_30241_, _30239_, _30238_);
  nor (_30242_, _30241_, _07793_);
  and (_30243_, _13353_, _05278_);
  nor (_30244_, _30243_, _30238_);
  nor (_30245_, _30244_, _07778_);
  and (_30246_, _06455_, _05278_);
  or (_30247_, _30246_, _30238_);
  and (_30248_, _30247_, _04481_);
  and (_30249_, _05278_, \oc8051_golden_model_1.ACC [6]);
  nor (_30250_, _30249_, _30238_);
  nor (_30252_, _30250_, _03737_);
  nor (_30253_, _30250_, _09029_);
  nor (_30254_, _04409_, _30237_);
  or (_30255_, _30254_, _30253_);
  and (_30256_, _30255_, _04081_);
  nor (_30257_, _13242_, _10991_);
  nor (_30258_, _30257_, _30238_);
  nor (_30259_, _30258_, _04081_);
  or (_30260_, _30259_, _30256_);
  and (_30261_, _30260_, _03996_);
  nor (_30263_, _05363_, _10991_);
  nor (_30264_, _30263_, _30238_);
  nor (_30265_, _30264_, _03996_);
  nor (_30266_, _30265_, _30261_);
  nor (_30267_, _30266_, _03729_);
  or (_30268_, _30267_, _07390_);
  nor (_30269_, _30268_, _30252_);
  and (_30270_, _30264_, _07390_);
  or (_30271_, _30270_, _04481_);
  nor (_30272_, _30271_, _30269_);
  or (_30274_, _30272_, _30248_);
  and (_30275_, _30274_, _03589_);
  nor (_30276_, _13332_, _10991_);
  nor (_30277_, _30276_, _30238_);
  nor (_30278_, _30277_, _03589_);
  or (_30279_, _30278_, _08828_);
  or (_30280_, _30279_, _30275_);
  and (_30281_, _13347_, _05278_);
  or (_30282_, _30238_, _07766_);
  or (_30283_, _30282_, _30281_);
  and (_30285_, _13339_, _05278_);
  nor (_30286_, _30285_, _30238_);
  and (_30287_, _30286_, _03601_);
  nor (_30288_, _30287_, _03780_);
  and (_30289_, _30288_, _30283_);
  and (_30290_, _30289_, _30280_);
  nor (_30291_, _30290_, _30245_);
  nor (_30292_, _30291_, _03622_);
  nor (_30293_, _30238_, _05412_);
  not (_30294_, _30293_);
  nor (_30296_, _30286_, _07777_);
  and (_30297_, _30296_, _30294_);
  nor (_30298_, _30297_, _30292_);
  nor (_30299_, _30298_, _03790_);
  nor (_30300_, _30250_, _06828_);
  and (_30301_, _30300_, _30294_);
  or (_30302_, _30301_, _30299_);
  and (_30303_, _30302_, _07795_);
  nor (_30304_, _13346_, _10991_);
  nor (_30305_, _30304_, _30238_);
  nor (_30307_, _30305_, _07795_);
  or (_30308_, _30307_, _30303_);
  and (_30309_, _30308_, _07793_);
  nor (_30310_, _30309_, _30242_);
  nor (_30311_, _30310_, _03815_);
  nor (_30312_, _30258_, _04246_);
  or (_30313_, _30312_, _03447_);
  nor (_30314_, _30313_, _30311_);
  and (_30315_, _13402_, _05278_);
  or (_30316_, _30238_, _03514_);
  nor (_30318_, _30316_, _30315_);
  nor (_30319_, _30318_, _30314_);
  or (_30320_, _30319_, _43004_);
  or (_30321_, _43000_, \oc8051_golden_model_1.TH1 [6]);
  and (_30322_, _30321_, _41806_);
  and (_43639_, _30322_, _30320_);
  not (_30323_, \oc8051_golden_model_1.TL0 [0]);
  nor (_30324_, _05284_, _30323_);
  nor (_30325_, _05666_, _11072_);
  nor (_30326_, _30325_, _30324_);
  and (_30328_, _30326_, _17166_);
  and (_30329_, _05284_, \oc8051_golden_model_1.ACC [0]);
  nor (_30330_, _30329_, _30324_);
  nor (_30331_, _30330_, _03737_);
  nor (_30332_, _30331_, _07390_);
  nor (_30333_, _30326_, _04081_);
  nor (_30334_, _04409_, _30323_);
  nor (_30335_, _30330_, _09029_);
  nor (_30336_, _30335_, _30334_);
  nor (_30337_, _30336_, _03610_);
  or (_30339_, _30337_, _03723_);
  nor (_30340_, _30339_, _30333_);
  or (_30341_, _30340_, _03729_);
  and (_30342_, _30341_, _30332_);
  and (_30343_, _05284_, _04620_);
  or (_30344_, _30324_, _25480_);
  nor (_30345_, _30344_, _30343_);
  nor (_30346_, _30345_, _30342_);
  nor (_30347_, _30346_, _04481_);
  and (_30348_, _06546_, _05284_);
  nor (_30350_, _30324_, _07400_);
  not (_30351_, _30350_);
  nor (_30352_, _30351_, _30348_);
  nor (_30353_, _30352_, _30347_);
  nor (_30354_, _30353_, _03222_);
  nor (_30355_, _12109_, _11072_);
  or (_30356_, _30324_, _03589_);
  nor (_30357_, _30356_, _30355_);
  or (_30358_, _30357_, _03601_);
  nor (_30359_, _30358_, _30354_);
  and (_30361_, _05284_, _06274_);
  nor (_30362_, _30361_, _30324_);
  nor (_30363_, _30362_, _05886_);
  or (_30364_, _30363_, _30359_);
  and (_30365_, _30364_, _07766_);
  and (_30366_, _12124_, _05284_);
  nor (_30367_, _30366_, _30324_);
  nor (_30368_, _30367_, _07766_);
  or (_30369_, _30368_, _30365_);
  nor (_30370_, _30369_, _03780_);
  and (_30372_, _12128_, _05284_);
  or (_30373_, _30324_, _07778_);
  nor (_30374_, _30373_, _30372_);
  or (_30375_, _30374_, _03622_);
  nor (_30376_, _30375_, _30370_);
  or (_30377_, _30362_, _07777_);
  nor (_30378_, _30377_, _30325_);
  nor (_30379_, _30378_, _30376_);
  nor (_30380_, _30379_, _03790_);
  nor (_30381_, _30324_, _05666_);
  or (_30383_, _30381_, _06828_);
  nor (_30384_, _30383_, _30330_);
  or (_30385_, _30384_, _30380_);
  and (_30386_, _30385_, _07795_);
  nor (_30387_, _12122_, _11072_);
  nor (_30388_, _30387_, _30324_);
  nor (_30389_, _30388_, _07795_);
  or (_30390_, _30389_, _30386_);
  and (_30391_, _30390_, _07793_);
  nor (_30392_, _12003_, _11072_);
  nor (_30393_, _30392_, _30324_);
  nor (_30394_, _30393_, _07793_);
  nor (_30395_, _30394_, _17166_);
  not (_30396_, _30395_);
  nor (_30397_, _30396_, _30391_);
  nor (_30398_, _30397_, _30328_);
  or (_30399_, _30398_, _43004_);
  or (_30400_, _43000_, \oc8051_golden_model_1.TL0 [0]);
  and (_30401_, _30400_, _41806_);
  and (_43640_, _30401_, _30399_);
  and (_30404_, _06501_, _05284_);
  not (_30405_, \oc8051_golden_model_1.TL0 [1]);
  nor (_30406_, _05284_, _30405_);
  nor (_30407_, _30406_, _07400_);
  not (_30408_, _30407_);
  nor (_30409_, _30408_, _30404_);
  not (_30410_, _30409_);
  and (_30411_, _05284_, _06764_);
  nor (_30412_, _30411_, _30406_);
  and (_30413_, _30412_, _07390_);
  nor (_30415_, _05284_, \oc8051_golden_model_1.TL0 [1]);
  and (_30416_, _05284_, _03274_);
  nor (_30417_, _30416_, _30415_);
  and (_30418_, _30417_, _03729_);
  and (_30419_, _30417_, _04409_);
  nor (_30420_, _04409_, _30405_);
  or (_30421_, _30420_, _30419_);
  and (_30422_, _30421_, _04081_);
  and (_30423_, _12213_, _05284_);
  nor (_30424_, _30423_, _30415_);
  and (_30426_, _30424_, _03610_);
  or (_30427_, _30426_, _30422_);
  and (_30428_, _30427_, _03996_);
  nor (_30429_, _30412_, _03996_);
  nor (_30430_, _30429_, _30428_);
  nor (_30431_, _30430_, _03729_);
  or (_30432_, _30431_, _07390_);
  nor (_30433_, _30432_, _30418_);
  nor (_30434_, _30433_, _30413_);
  nor (_30435_, _30434_, _04481_);
  nor (_30437_, _30435_, _03222_);
  and (_30438_, _30437_, _30410_);
  not (_30439_, _30415_);
  and (_30440_, _12313_, _05284_);
  nor (_30441_, _30440_, _03589_);
  and (_30442_, _30441_, _30439_);
  nor (_30443_, _30442_, _30438_);
  nor (_30444_, _30443_, _08828_);
  nor (_30445_, _12327_, _11072_);
  nor (_30446_, _30445_, _07766_);
  and (_30448_, _05284_, _04303_);
  nor (_30449_, _30448_, _05886_);
  nor (_30450_, _30449_, _30446_);
  nor (_30451_, _30450_, _30415_);
  nor (_30452_, _30451_, _30444_);
  nor (_30453_, _30452_, _03780_);
  nor (_30454_, _12333_, _11072_);
  nor (_30455_, _30454_, _07778_);
  and (_30456_, _30455_, _30439_);
  nor (_30457_, _30456_, _30453_);
  nor (_30459_, _30457_, _03622_);
  nor (_30460_, _12207_, _11072_);
  nor (_30461_, _30460_, _07777_);
  and (_30462_, _30461_, _30439_);
  nor (_30463_, _30462_, _30459_);
  nor (_30464_, _30463_, _03790_);
  nor (_30465_, _30406_, _05618_);
  nor (_30466_, _30465_, _06828_);
  and (_30467_, _30466_, _30417_);
  nor (_30469_, _30467_, _30464_);
  or (_30472_, _30469_, _18499_);
  and (_30474_, _30416_, _05617_);
  nor (_30476_, _30474_, _07793_);
  and (_30478_, _30476_, _30439_);
  nor (_30480_, _30478_, _03815_);
  and (_30482_, _30448_, _05617_);
  or (_30484_, _30415_, _07795_);
  or (_30486_, _30484_, _30482_);
  and (_30488_, _30486_, _30480_);
  and (_30490_, _30488_, _30472_);
  nor (_30492_, _30424_, _04246_);
  nor (_30493_, _30492_, _30490_);
  and (_30494_, _30493_, _03514_);
  nor (_30495_, _30423_, _30406_);
  nor (_30496_, _30495_, _03514_);
  or (_30497_, _30496_, _30494_);
  or (_30498_, _30497_, _43004_);
  or (_30499_, _43000_, \oc8051_golden_model_1.TL0 [1]);
  and (_30500_, _30499_, _41806_);
  and (_43643_, _30500_, _30498_);
  not (_30502_, \oc8051_golden_model_1.TL0 [2]);
  nor (_30503_, _05284_, _30502_);
  nor (_30504_, _12538_, _11072_);
  nor (_30505_, _30504_, _30503_);
  nor (_30506_, _30505_, _07793_);
  nor (_30507_, _11072_, _04875_);
  nor (_30508_, _30507_, _30503_);
  and (_30509_, _30508_, _07390_);
  nor (_30510_, _12416_, _11072_);
  nor (_30511_, _30510_, _30503_);
  nor (_30513_, _30511_, _04081_);
  nor (_30514_, _04409_, _30502_);
  and (_30515_, _05284_, \oc8051_golden_model_1.ACC [2]);
  nor (_30516_, _30515_, _30503_);
  nor (_30517_, _30516_, _09029_);
  nor (_30518_, _30517_, _30514_);
  nor (_30519_, _30518_, _03610_);
  or (_30520_, _30519_, _30513_);
  and (_30521_, _30520_, _03996_);
  nor (_30522_, _30508_, _03996_);
  or (_30524_, _30522_, _30521_);
  and (_30525_, _30524_, _03737_);
  nor (_30526_, _30516_, _03737_);
  nor (_30527_, _30526_, _07390_);
  not (_30528_, _30527_);
  nor (_30529_, _30528_, _30525_);
  nor (_30530_, _30529_, _30509_);
  nor (_30531_, _30530_, _04481_);
  and (_30532_, _06637_, _05284_);
  nor (_30533_, _30503_, _07400_);
  not (_30535_, _30533_);
  nor (_30536_, _30535_, _30532_);
  nor (_30537_, _30536_, _30531_);
  nor (_30538_, _30537_, _03222_);
  nor (_30539_, _12519_, _11072_);
  or (_30540_, _30503_, _03589_);
  nor (_30541_, _30540_, _30539_);
  or (_30542_, _30541_, _03601_);
  nor (_30543_, _30542_, _30538_);
  and (_30544_, _05284_, _06332_);
  nor (_30546_, _30544_, _30503_);
  nor (_30547_, _30546_, _05886_);
  or (_30548_, _30547_, _30543_);
  and (_30549_, _30548_, _07766_);
  and (_30550_, _12533_, _05284_);
  nor (_30551_, _30550_, _30503_);
  nor (_30552_, _30551_, _07766_);
  or (_30553_, _30552_, _30549_);
  nor (_30554_, _30553_, _03780_);
  and (_30555_, _12539_, _05284_);
  or (_30557_, _30503_, _07778_);
  nor (_30558_, _30557_, _30555_);
  or (_30559_, _30558_, _03622_);
  nor (_30560_, _30559_, _30554_);
  nor (_30561_, _30503_, _05718_);
  or (_30562_, _30546_, _07777_);
  nor (_30563_, _30562_, _30561_);
  nor (_30564_, _30563_, _30560_);
  nor (_30565_, _30564_, _03790_);
  or (_30566_, _30561_, _06828_);
  or (_30568_, _30566_, _30516_);
  and (_30569_, _30568_, _07795_);
  not (_30570_, _30569_);
  nor (_30571_, _30570_, _30565_);
  nor (_30572_, _12532_, _11072_);
  or (_30573_, _30503_, _07795_);
  nor (_30574_, _30573_, _30572_);
  or (_30575_, _30574_, _03785_);
  nor (_30576_, _30575_, _30571_);
  nor (_30577_, _30576_, _30506_);
  nor (_30579_, _30577_, _03815_);
  nor (_30580_, _30511_, _04246_);
  or (_30581_, _30580_, _03447_);
  nor (_30582_, _30581_, _30579_);
  and (_30583_, _12592_, _05284_);
  or (_30584_, _30503_, _03514_);
  nor (_30585_, _30584_, _30583_);
  nor (_30586_, _30585_, _30582_);
  or (_30587_, _30586_, _43004_);
  or (_30588_, _43000_, \oc8051_golden_model_1.TL0 [2]);
  and (_30590_, _30588_, _41806_);
  and (_43644_, _30590_, _30587_);
  not (_30591_, \oc8051_golden_model_1.TL0 [3]);
  nor (_30592_, _05284_, _30591_);
  nor (_30593_, _12738_, _11072_);
  nor (_30594_, _30593_, _30592_);
  nor (_30595_, _30594_, _07793_);
  and (_30596_, _12739_, _05284_);
  nor (_30597_, _30596_, _30592_);
  nor (_30598_, _30597_, _07778_);
  and (_30600_, _06592_, _05284_);
  or (_30601_, _30600_, _30592_);
  and (_30602_, _30601_, _04481_);
  and (_30603_, _05284_, \oc8051_golden_model_1.ACC [3]);
  nor (_30604_, _30603_, _30592_);
  nor (_30605_, _30604_, _03737_);
  nor (_30606_, _30604_, _09029_);
  nor (_30607_, _04409_, _30591_);
  or (_30608_, _30607_, _30606_);
  and (_30609_, _30608_, _04081_);
  nor (_30611_, _12627_, _11072_);
  nor (_30612_, _30611_, _30592_);
  nor (_30613_, _30612_, _04081_);
  or (_30614_, _30613_, _30609_);
  and (_30615_, _30614_, _03996_);
  nor (_30616_, _11072_, _05005_);
  nor (_30617_, _30616_, _30592_);
  nor (_30618_, _30617_, _03996_);
  nor (_30619_, _30618_, _30615_);
  nor (_30620_, _30619_, _03729_);
  or (_30622_, _30620_, _07390_);
  nor (_30623_, _30622_, _30605_);
  and (_30624_, _30617_, _07390_);
  or (_30625_, _30624_, _04481_);
  nor (_30626_, _30625_, _30623_);
  or (_30627_, _30626_, _30602_);
  and (_30628_, _30627_, _03589_);
  nor (_30629_, _12718_, _11072_);
  nor (_30630_, _30629_, _30592_);
  nor (_30631_, _30630_, _03589_);
  or (_30633_, _30631_, _08828_);
  or (_30634_, _30633_, _30628_);
  and (_30635_, _12733_, _05284_);
  or (_30636_, _30592_, _07766_);
  or (_30637_, _30636_, _30635_);
  and (_30638_, _05284_, _06276_);
  nor (_30639_, _30638_, _30592_);
  and (_30640_, _30639_, _03601_);
  nor (_30641_, _30640_, _03780_);
  and (_30642_, _30641_, _30637_);
  and (_30644_, _30642_, _30634_);
  nor (_30645_, _30644_, _30598_);
  nor (_30646_, _30645_, _03622_);
  nor (_30647_, _30592_, _05567_);
  not (_30648_, _30647_);
  nor (_30649_, _30639_, _07777_);
  and (_30650_, _30649_, _30648_);
  nor (_30651_, _30650_, _30646_);
  nor (_30652_, _30651_, _03790_);
  nor (_30653_, _30604_, _06828_);
  and (_30655_, _30653_, _30648_);
  or (_30656_, _30655_, _30652_);
  and (_30657_, _30656_, _07795_);
  nor (_30658_, _12732_, _11072_);
  nor (_30659_, _30658_, _30592_);
  nor (_30660_, _30659_, _07795_);
  or (_30661_, _30660_, _30657_);
  and (_30662_, _30661_, _07793_);
  nor (_30663_, _30662_, _30595_);
  nor (_30664_, _30663_, _03815_);
  nor (_30666_, _30612_, _04246_);
  or (_30667_, _30666_, _03447_);
  nor (_30668_, _30667_, _30664_);
  and (_30669_, _12794_, _05284_);
  or (_30670_, _30592_, _03514_);
  nor (_30671_, _30670_, _30669_);
  nor (_30672_, _30671_, _30668_);
  or (_30673_, _30672_, _43004_);
  or (_30674_, _43000_, \oc8051_golden_model_1.TL0 [3]);
  and (_30675_, _30674_, _41806_);
  and (_43645_, _30675_, _30673_);
  not (_30677_, \oc8051_golden_model_1.TL0 [4]);
  nor (_30678_, _05284_, _30677_);
  nor (_30679_, _12816_, _11072_);
  nor (_30680_, _30679_, _30678_);
  nor (_30681_, _30680_, _07793_);
  and (_30682_, _12817_, _05284_);
  nor (_30683_, _30682_, _30678_);
  nor (_30684_, _30683_, _07778_);
  and (_30685_, _06298_, _05284_);
  nor (_30687_, _30685_, _30678_);
  and (_30688_, _30687_, _03601_);
  nor (_30689_, _05777_, _11072_);
  nor (_30690_, _30689_, _30678_);
  and (_30691_, _30690_, _07390_);
  and (_30692_, _05284_, \oc8051_golden_model_1.ACC [4]);
  nor (_30693_, _30692_, _30678_);
  nor (_30694_, _30693_, _03737_);
  nor (_30695_, _30693_, _09029_);
  nor (_30696_, _04409_, _30677_);
  or (_30698_, _30696_, _30695_);
  and (_30699_, _30698_, _04081_);
  nor (_30700_, _12841_, _11072_);
  nor (_30701_, _30700_, _30678_);
  nor (_30702_, _30701_, _04081_);
  or (_30703_, _30702_, _30699_);
  and (_30704_, _30703_, _03996_);
  nor (_30705_, _30690_, _03996_);
  nor (_30706_, _30705_, _30704_);
  nor (_30707_, _30706_, _03729_);
  or (_30709_, _30707_, _07390_);
  nor (_30710_, _30709_, _30694_);
  nor (_30711_, _30710_, _30691_);
  nor (_30712_, _30711_, _04481_);
  and (_30713_, _06730_, _05284_);
  nor (_30714_, _30678_, _07400_);
  not (_30715_, _30714_);
  nor (_30716_, _30715_, _30713_);
  or (_30717_, _30716_, _03222_);
  nor (_30718_, _30717_, _30712_);
  nor (_30720_, _12933_, _11072_);
  nor (_30721_, _30720_, _30678_);
  nor (_30722_, _30721_, _03589_);
  or (_30723_, _30722_, _03601_);
  nor (_30724_, _30723_, _30718_);
  nor (_30725_, _30724_, _30688_);
  or (_30726_, _30725_, _03600_);
  and (_30727_, _12821_, _05284_);
  or (_30728_, _30727_, _30678_);
  or (_30729_, _30728_, _07766_);
  and (_30731_, _30729_, _07778_);
  and (_30732_, _30731_, _30726_);
  nor (_30733_, _30732_, _30684_);
  nor (_30734_, _30733_, _03622_);
  nor (_30735_, _30678_, _05825_);
  not (_30736_, _30735_);
  nor (_30737_, _30687_, _07777_);
  and (_30738_, _30737_, _30736_);
  nor (_30739_, _30738_, _30734_);
  nor (_30740_, _30739_, _03790_);
  nor (_30742_, _30693_, _06828_);
  and (_30743_, _30742_, _30736_);
  or (_30744_, _30743_, _30740_);
  and (_30745_, _30744_, _07795_);
  nor (_30746_, _12819_, _11072_);
  nor (_30747_, _30746_, _30678_);
  nor (_30748_, _30747_, _07795_);
  or (_30749_, _30748_, _30745_);
  and (_30750_, _30749_, _07793_);
  nor (_30751_, _30750_, _30681_);
  nor (_30753_, _30751_, _03815_);
  nor (_30754_, _30701_, _04246_);
  or (_30755_, _30754_, _03447_);
  nor (_30756_, _30755_, _30753_);
  and (_30757_, _13003_, _05284_);
  or (_30758_, _30678_, _03514_);
  nor (_30759_, _30758_, _30757_);
  nor (_30760_, _30759_, _30756_);
  or (_30761_, _30760_, _43004_);
  or (_30762_, _43000_, \oc8051_golden_model_1.TL0 [4]);
  and (_30764_, _30762_, _41806_);
  and (_43646_, _30764_, _30761_);
  not (_30765_, \oc8051_golden_model_1.TL0 [5]);
  nor (_30766_, _05284_, _30765_);
  nor (_30767_, _13146_, _11072_);
  nor (_30768_, _30767_, _30766_);
  nor (_30769_, _30768_, _07793_);
  and (_30770_, _13147_, _05284_);
  nor (_30771_, _30770_, _30766_);
  nor (_30772_, _30771_, _07778_);
  and (_30774_, _06684_, _05284_);
  or (_30775_, _30774_, _30766_);
  and (_30776_, _30775_, _04481_);
  and (_30777_, _05284_, \oc8051_golden_model_1.ACC [5]);
  nor (_30778_, _30777_, _30766_);
  nor (_30779_, _30778_, _03737_);
  nor (_30780_, _30778_, _09029_);
  nor (_30781_, _04409_, _30765_);
  or (_30782_, _30781_, _30780_);
  and (_30783_, _30782_, _04081_);
  nor (_30785_, _13014_, _11072_);
  nor (_30786_, _30785_, _30766_);
  nor (_30787_, _30786_, _04081_);
  or (_30788_, _30787_, _30783_);
  and (_30789_, _30788_, _03996_);
  nor (_30790_, _05469_, _11072_);
  nor (_30791_, _30790_, _30766_);
  nor (_30792_, _30791_, _03996_);
  nor (_30793_, _30792_, _30789_);
  nor (_30794_, _30793_, _03729_);
  or (_30796_, _30794_, _07390_);
  nor (_30797_, _30796_, _30779_);
  and (_30798_, _30791_, _07390_);
  or (_30799_, _30798_, _04481_);
  nor (_30800_, _30799_, _30797_);
  or (_30801_, _30800_, _30776_);
  and (_30802_, _30801_, _03589_);
  nor (_30803_, _13127_, _11072_);
  nor (_30804_, _30803_, _30766_);
  nor (_30805_, _30804_, _03589_);
  or (_30807_, _30805_, _08828_);
  or (_30808_, _30807_, _30802_);
  and (_30809_, _13141_, _05284_);
  or (_30810_, _30766_, _07766_);
  or (_30811_, _30810_, _30809_);
  and (_30812_, _06306_, _05284_);
  nor (_30813_, _30812_, _30766_);
  and (_30814_, _30813_, _03601_);
  nor (_30815_, _30814_, _03780_);
  and (_30816_, _30815_, _30811_);
  and (_30817_, _30816_, _30808_);
  nor (_30818_, _30817_, _30772_);
  nor (_30819_, _30818_, _03622_);
  nor (_30820_, _30766_, _05518_);
  not (_30821_, _30820_);
  nor (_30822_, _30813_, _07777_);
  and (_30823_, _30822_, _30821_);
  nor (_30824_, _30823_, _30819_);
  nor (_30825_, _30824_, _03790_);
  nor (_30826_, _30778_, _06828_);
  and (_30828_, _30826_, _30821_);
  nor (_30829_, _30828_, _03624_);
  not (_30830_, _30829_);
  nor (_30831_, _30830_, _30825_);
  nor (_30832_, _13140_, _11072_);
  or (_30833_, _30766_, _07795_);
  nor (_30834_, _30833_, _30832_);
  or (_30835_, _30834_, _03785_);
  nor (_30836_, _30835_, _30831_);
  nor (_30837_, _30836_, _30769_);
  nor (_30839_, _30837_, _03815_);
  nor (_30840_, _30786_, _04246_);
  or (_30841_, _30840_, _03447_);
  nor (_30842_, _30841_, _30839_);
  and (_30843_, _13199_, _05284_);
  or (_30844_, _30766_, _03514_);
  nor (_30845_, _30844_, _30843_);
  nor (_30846_, _30845_, _30842_);
  or (_30847_, _30846_, _43004_);
  or (_30848_, _43000_, \oc8051_golden_model_1.TL0 [5]);
  and (_30850_, _30848_, _41806_);
  and (_43647_, _30850_, _30847_);
  not (_30851_, \oc8051_golden_model_1.TL0 [6]);
  nor (_30852_, _05284_, _30851_);
  nor (_30853_, _13352_, _11072_);
  nor (_30854_, _30853_, _30852_);
  nor (_30855_, _30854_, _07793_);
  and (_30856_, _13353_, _05284_);
  nor (_30857_, _30856_, _30852_);
  nor (_30858_, _30857_, _07778_);
  and (_30860_, _06455_, _05284_);
  or (_30861_, _30860_, _30852_);
  and (_30862_, _30861_, _04481_);
  and (_30863_, _05284_, \oc8051_golden_model_1.ACC [6]);
  nor (_30864_, _30863_, _30852_);
  nor (_30865_, _30864_, _03737_);
  nor (_30866_, _30864_, _09029_);
  nor (_30867_, _04409_, _30851_);
  or (_30868_, _30867_, _30866_);
  and (_30869_, _30868_, _04081_);
  nor (_30871_, _13242_, _11072_);
  nor (_30872_, _30871_, _30852_);
  nor (_30873_, _30872_, _04081_);
  or (_30874_, _30873_, _30869_);
  and (_30875_, _30874_, _03996_);
  nor (_30876_, _05363_, _11072_);
  nor (_30877_, _30876_, _30852_);
  nor (_30878_, _30877_, _03996_);
  nor (_30879_, _30878_, _30875_);
  nor (_30880_, _30879_, _03729_);
  or (_30881_, _30880_, _07390_);
  nor (_30882_, _30881_, _30865_);
  and (_30883_, _30877_, _07390_);
  or (_30884_, _30883_, _04481_);
  nor (_30885_, _30884_, _30882_);
  or (_30886_, _30885_, _30862_);
  and (_30887_, _30886_, _03589_);
  nor (_30888_, _13332_, _11072_);
  nor (_30889_, _30888_, _30852_);
  nor (_30890_, _30889_, _03589_);
  or (_30893_, _30890_, _08828_);
  or (_30894_, _30893_, _30887_);
  and (_30895_, _13347_, _05284_);
  or (_30896_, _30852_, _07766_);
  or (_30897_, _30896_, _30895_);
  and (_30898_, _13339_, _05284_);
  nor (_30899_, _30898_, _30852_);
  and (_30900_, _30899_, _03601_);
  nor (_30901_, _30900_, _03780_);
  and (_30902_, _30901_, _30897_);
  and (_30904_, _30902_, _30894_);
  nor (_30905_, _30904_, _30858_);
  nor (_30906_, _30905_, _03622_);
  nor (_30907_, _30852_, _05412_);
  not (_30908_, _30907_);
  nor (_30909_, _30899_, _07777_);
  and (_30910_, _30909_, _30908_);
  nor (_30911_, _30910_, _30906_);
  nor (_30912_, _30911_, _03790_);
  nor (_30913_, _30864_, _06828_);
  and (_30915_, _30913_, _30908_);
  nor (_30916_, _30915_, _03624_);
  not (_30917_, _30916_);
  nor (_30918_, _30917_, _30912_);
  nor (_30919_, _13346_, _11072_);
  or (_30920_, _30852_, _07795_);
  nor (_30921_, _30920_, _30919_);
  or (_30922_, _30921_, _03785_);
  nor (_30923_, _30922_, _30918_);
  nor (_30924_, _30923_, _30855_);
  nor (_30926_, _30924_, _03815_);
  nor (_30927_, _30872_, _04246_);
  or (_30928_, _30927_, _03447_);
  nor (_30929_, _30928_, _30926_);
  and (_30930_, _13402_, _05284_);
  or (_30931_, _30852_, _03514_);
  nor (_30932_, _30931_, _30930_);
  nor (_30933_, _30932_, _30929_);
  or (_30934_, _30933_, _43004_);
  or (_30935_, _43000_, \oc8051_golden_model_1.TL0 [6]);
  and (_30937_, _30935_, _41806_);
  and (_43648_, _30937_, _30934_);
  not (_30938_, \oc8051_golden_model_1.TL1 [0]);
  nor (_30939_, _05271_, _30938_);
  nor (_30940_, _05666_, _11154_);
  nor (_30941_, _30940_, _30939_);
  and (_30942_, _30941_, _17166_);
  and (_30943_, _05271_, \oc8051_golden_model_1.ACC [0]);
  nor (_30944_, _30943_, _30939_);
  nor (_30945_, _30944_, _03737_);
  nor (_30947_, _30944_, _09029_);
  nor (_30948_, _04409_, _30938_);
  or (_30949_, _30948_, _30947_);
  and (_30950_, _30949_, _04081_);
  nor (_30951_, _30941_, _04081_);
  or (_30952_, _30951_, _30950_);
  and (_30953_, _30952_, _03996_);
  and (_30954_, _05271_, _04620_);
  nor (_30955_, _30954_, _30939_);
  nor (_30956_, _30955_, _03996_);
  nor (_30958_, _30956_, _30953_);
  nor (_30959_, _30958_, _03729_);
  or (_30960_, _30959_, _07390_);
  nor (_30961_, _30960_, _30945_);
  and (_30962_, _30955_, _07390_);
  nor (_30963_, _30962_, _30961_);
  nor (_30964_, _30963_, _04481_);
  and (_30965_, _06546_, _05271_);
  nor (_30966_, _30939_, _07400_);
  not (_30967_, _30966_);
  nor (_30969_, _30967_, _30965_);
  nor (_30970_, _30969_, _30964_);
  nor (_30971_, _30970_, _03222_);
  nor (_30972_, _12109_, _11154_);
  or (_30973_, _30939_, _03589_);
  nor (_30974_, _30973_, _30972_);
  or (_30975_, _30974_, _03601_);
  nor (_30976_, _30975_, _30971_);
  and (_30977_, _05271_, _06274_);
  nor (_30978_, _30977_, _30939_);
  nor (_30980_, _30978_, _05886_);
  or (_30981_, _30980_, _30976_);
  and (_30982_, _30981_, _07766_);
  and (_30983_, _12124_, _05271_);
  nor (_30984_, _30983_, _30939_);
  nor (_30985_, _30984_, _07766_);
  or (_30986_, _30985_, _30982_);
  nor (_30987_, _30986_, _03780_);
  and (_30988_, _12128_, _05271_);
  or (_30989_, _30939_, _07778_);
  nor (_30991_, _30989_, _30988_);
  or (_30992_, _30991_, _03622_);
  nor (_30993_, _30992_, _30987_);
  or (_30994_, _30978_, _07777_);
  nor (_30995_, _30994_, _30940_);
  nor (_30996_, _30995_, _30993_);
  nor (_30997_, _30996_, _03790_);
  nor (_30998_, _30939_, _05666_);
  or (_30999_, _30998_, _06828_);
  nor (_31000_, _30999_, _30944_);
  or (_31002_, _31000_, _30997_);
  and (_31003_, _31002_, _07795_);
  nor (_31004_, _12122_, _11154_);
  nor (_31005_, _31004_, _30939_);
  nor (_31006_, _31005_, _07795_);
  or (_31007_, _31006_, _31003_);
  and (_31008_, _31007_, _07793_);
  nor (_31009_, _12003_, _11154_);
  nor (_31010_, _31009_, _30939_);
  nor (_31011_, _31010_, _07793_);
  nor (_31013_, _31011_, _17166_);
  not (_31014_, _31013_);
  nor (_31015_, _31014_, _31008_);
  nor (_31016_, _31015_, _30942_);
  or (_31017_, _31016_, _43004_);
  or (_31018_, _43000_, \oc8051_golden_model_1.TL1 [0]);
  and (_31019_, _31018_, _41806_);
  and (_43649_, _31019_, _31017_);
  and (_31020_, _06501_, _05271_);
  not (_31021_, \oc8051_golden_model_1.TL1 [1]);
  nor (_31023_, _05271_, _31021_);
  nor (_31024_, _31023_, _07400_);
  not (_31025_, _31024_);
  nor (_31026_, _31025_, _31020_);
  not (_31027_, _31026_);
  nor (_31028_, _05271_, \oc8051_golden_model_1.TL1 [1]);
  and (_31029_, _05271_, _03274_);
  nor (_31030_, _31029_, _31028_);
  and (_31031_, _31030_, _03729_);
  and (_31032_, _31030_, _04409_);
  nor (_31034_, _04409_, _31021_);
  or (_31035_, _31034_, _31032_);
  and (_31036_, _31035_, _04081_);
  and (_31037_, _12213_, _05271_);
  nor (_31038_, _31037_, _31028_);
  and (_31039_, _31038_, _03610_);
  or (_31040_, _31039_, _31036_);
  and (_31041_, _31040_, _03996_);
  and (_31042_, _05271_, _06764_);
  nor (_31043_, _31042_, _31023_);
  nor (_31045_, _31043_, _03996_);
  nor (_31046_, _31045_, _31041_);
  nor (_31047_, _31046_, _03729_);
  or (_31048_, _31047_, _07390_);
  nor (_31049_, _31048_, _31031_);
  and (_31050_, _31043_, _07390_);
  nor (_31051_, _31050_, _31049_);
  nor (_31052_, _31051_, _04481_);
  nor (_31053_, _31052_, _03222_);
  and (_31054_, _31053_, _31027_);
  not (_31056_, _31028_);
  and (_31057_, _12313_, _05271_);
  nor (_31058_, _31057_, _03589_);
  and (_31059_, _31058_, _31056_);
  nor (_31060_, _31059_, _31054_);
  nor (_31061_, _31060_, _08828_);
  nor (_31062_, _12327_, _11154_);
  nor (_31063_, _31062_, _07766_);
  and (_31064_, _05271_, _04303_);
  nor (_31065_, _31064_, _05886_);
  nor (_31067_, _31065_, _31063_);
  nor (_31068_, _31067_, _31028_);
  nor (_31069_, _31068_, _31061_);
  nor (_31070_, _31069_, _03780_);
  nor (_31071_, _12333_, _11154_);
  nor (_31072_, _31071_, _07778_);
  and (_31073_, _31072_, _31056_);
  nor (_31074_, _31073_, _31070_);
  nor (_31075_, _31074_, _03622_);
  nor (_31076_, _12207_, _11154_);
  nor (_31078_, _31076_, _07777_);
  and (_31079_, _31078_, _31056_);
  nor (_31080_, _31079_, _31075_);
  nor (_31081_, _31080_, _03790_);
  nor (_31082_, _31023_, _05618_);
  nor (_31083_, _31082_, _06828_);
  and (_31084_, _31083_, _31030_);
  nor (_31085_, _31084_, _31081_);
  or (_31086_, _31085_, _18499_);
  and (_31087_, _31064_, _05617_);
  nor (_31089_, _31087_, _07795_);
  and (_31090_, _31089_, _31056_);
  not (_31091_, _31090_);
  nand (_31092_, _31029_, _05617_);
  nor (_31093_, _31028_, _07793_);
  and (_31094_, _31093_, _31092_);
  nor (_31095_, _31094_, _03815_);
  and (_31096_, _31095_, _31091_);
  and (_31097_, _31096_, _31086_);
  nor (_31098_, _31038_, _04246_);
  nor (_31100_, _31098_, _31097_);
  and (_31101_, _31100_, _03514_);
  nor (_31102_, _31037_, _31023_);
  nor (_31103_, _31102_, _03514_);
  or (_31104_, _31103_, _31101_);
  or (_31105_, _31104_, _43004_);
  or (_31106_, _43000_, \oc8051_golden_model_1.TL1 [1]);
  and (_31107_, _31106_, _41806_);
  and (_43650_, _31107_, _31105_);
  not (_31108_, \oc8051_golden_model_1.TL1 [2]);
  nor (_31109_, _05271_, _31108_);
  nor (_31110_, _12538_, _11154_);
  nor (_31111_, _31110_, _31109_);
  nor (_31112_, _31111_, _07793_);
  and (_31113_, _12539_, _05271_);
  nor (_31114_, _31113_, _31109_);
  nor (_31115_, _31114_, _07778_);
  and (_31116_, _05271_, \oc8051_golden_model_1.ACC [2]);
  nor (_31117_, _31116_, _31109_);
  nor (_31118_, _31117_, _03737_);
  nor (_31121_, _31117_, _09029_);
  nor (_31122_, _04409_, _31108_);
  or (_31123_, _31122_, _31121_);
  and (_31124_, _31123_, _04081_);
  nor (_31125_, _12416_, _11154_);
  nor (_31126_, _31125_, _31109_);
  nor (_31127_, _31126_, _04081_);
  or (_31128_, _31127_, _31124_);
  and (_31129_, _31128_, _03996_);
  nor (_31130_, _11154_, _04875_);
  nor (_31132_, _31130_, _31109_);
  nor (_31133_, _31132_, _03996_);
  nor (_31134_, _31133_, _31129_);
  nor (_31135_, _31134_, _03729_);
  or (_31136_, _31135_, _07390_);
  nor (_31137_, _31136_, _31118_);
  and (_31138_, _31132_, _07390_);
  nor (_31139_, _31138_, _31137_);
  nor (_31140_, _31139_, _04481_);
  and (_31141_, _06637_, _05271_);
  nor (_31143_, _31109_, _07400_);
  not (_31144_, _31143_);
  nor (_31145_, _31144_, _31141_);
  nor (_31146_, _31145_, _03222_);
  not (_31147_, _31146_);
  nor (_31148_, _31147_, _31140_);
  nor (_31149_, _12519_, _11154_);
  nor (_31150_, _31149_, _31109_);
  nor (_31151_, _31150_, _03589_);
  or (_31152_, _31151_, _08828_);
  or (_31154_, _31152_, _31148_);
  and (_31155_, _12533_, _05271_);
  or (_31156_, _31109_, _07766_);
  or (_31157_, _31156_, _31155_);
  and (_31158_, _05271_, _06332_);
  nor (_31159_, _31158_, _31109_);
  and (_31160_, _31159_, _03601_);
  nor (_31161_, _31160_, _03780_);
  and (_31162_, _31161_, _31157_);
  and (_31163_, _31162_, _31154_);
  nor (_31165_, _31163_, _31115_);
  nor (_31166_, _31165_, _03622_);
  nor (_31167_, _31109_, _05718_);
  not (_31168_, _31167_);
  nor (_31169_, _31159_, _07777_);
  and (_31170_, _31169_, _31168_);
  nor (_31171_, _31170_, _31166_);
  nor (_31172_, _31171_, _03790_);
  nor (_31173_, _31117_, _06828_);
  and (_31174_, _31173_, _31168_);
  nor (_31176_, _31174_, _03624_);
  not (_31177_, _31176_);
  nor (_31178_, _31177_, _31172_);
  nor (_31179_, _12532_, _11154_);
  or (_31180_, _31109_, _07795_);
  nor (_31181_, _31180_, _31179_);
  or (_31182_, _31181_, _03785_);
  nor (_31183_, _31182_, _31178_);
  nor (_31184_, _31183_, _31112_);
  nor (_31185_, _31184_, _03815_);
  nor (_31187_, _31126_, _04246_);
  or (_31188_, _31187_, _03447_);
  nor (_31189_, _31188_, _31185_);
  and (_31190_, _12592_, _05271_);
  or (_31191_, _31109_, _03514_);
  nor (_31192_, _31191_, _31190_);
  nor (_31193_, _31192_, _31189_);
  or (_31194_, _31193_, _43004_);
  or (_31195_, _43000_, \oc8051_golden_model_1.TL1 [2]);
  and (_31196_, _31195_, _41806_);
  and (_43651_, _31196_, _31194_);
  not (_31198_, \oc8051_golden_model_1.TL1 [3]);
  nor (_31199_, _05271_, _31198_);
  nor (_31200_, _12738_, _11154_);
  nor (_31201_, _31200_, _31199_);
  nor (_31202_, _31201_, _07793_);
  and (_31203_, _12739_, _05271_);
  nor (_31204_, _31203_, _31199_);
  nor (_31205_, _31204_, _07778_);
  and (_31206_, _06592_, _05271_);
  or (_31208_, _31206_, _31199_);
  and (_31209_, _31208_, _04481_);
  and (_31210_, _05271_, \oc8051_golden_model_1.ACC [3]);
  nor (_31211_, _31210_, _31199_);
  nor (_31212_, _31211_, _03737_);
  nor (_31213_, _31211_, _09029_);
  nor (_31214_, _04409_, _31198_);
  or (_31215_, _31214_, _31213_);
  and (_31216_, _31215_, _04081_);
  nor (_31217_, _12627_, _11154_);
  nor (_31219_, _31217_, _31199_);
  nor (_31220_, _31219_, _04081_);
  or (_31221_, _31220_, _31216_);
  and (_31222_, _31221_, _03996_);
  nor (_31223_, _11154_, _05005_);
  nor (_31224_, _31223_, _31199_);
  nor (_31225_, _31224_, _03996_);
  nor (_31226_, _31225_, _31222_);
  nor (_31227_, _31226_, _03729_);
  or (_31228_, _31227_, _07390_);
  nor (_31230_, _31228_, _31212_);
  and (_31231_, _31224_, _07390_);
  or (_31232_, _31231_, _04481_);
  nor (_31233_, _31232_, _31230_);
  or (_31234_, _31233_, _31209_);
  and (_31235_, _31234_, _03589_);
  nor (_31236_, _12718_, _11154_);
  nor (_31237_, _31236_, _31199_);
  nor (_31238_, _31237_, _03589_);
  or (_31239_, _31238_, _08828_);
  or (_31241_, _31239_, _31235_);
  and (_31242_, _12733_, _05271_);
  or (_31243_, _31199_, _07766_);
  or (_31244_, _31243_, _31242_);
  and (_31245_, _05271_, _06276_);
  nor (_31246_, _31245_, _31199_);
  and (_31247_, _31246_, _03601_);
  nor (_31248_, _31247_, _03780_);
  and (_31249_, _31248_, _31244_);
  and (_31250_, _31249_, _31241_);
  nor (_31252_, _31250_, _31205_);
  nor (_31253_, _31252_, _03622_);
  nor (_31254_, _31199_, _05567_);
  not (_31255_, _31254_);
  nor (_31256_, _31246_, _07777_);
  and (_31257_, _31256_, _31255_);
  nor (_31258_, _31257_, _31253_);
  nor (_31259_, _31258_, _03790_);
  nor (_31260_, _31211_, _06828_);
  and (_31261_, _31260_, _31255_);
  nor (_31263_, _31261_, _03624_);
  not (_31264_, _31263_);
  nor (_31265_, _31264_, _31259_);
  nor (_31266_, _12732_, _11154_);
  or (_31267_, _31199_, _07795_);
  nor (_31268_, _31267_, _31266_);
  or (_31269_, _31268_, _03785_);
  nor (_31270_, _31269_, _31265_);
  nor (_31271_, _31270_, _31202_);
  nor (_31272_, _31271_, _03815_);
  nor (_31274_, _31219_, _04246_);
  or (_31275_, _31274_, _03447_);
  nor (_31276_, _31275_, _31272_);
  and (_31277_, _12794_, _05271_);
  or (_31278_, _31199_, _03514_);
  nor (_31279_, _31278_, _31277_);
  nor (_31280_, _31279_, _31276_);
  or (_31281_, _31280_, _43004_);
  or (_31282_, _43000_, \oc8051_golden_model_1.TL1 [3]);
  and (_31283_, _31282_, _41806_);
  and (_43652_, _31283_, _31281_);
  not (_31285_, \oc8051_golden_model_1.TL1 [4]);
  nor (_31286_, _05271_, _31285_);
  nor (_31287_, _12816_, _11154_);
  nor (_31288_, _31287_, _31286_);
  nor (_31289_, _31288_, _07793_);
  and (_31290_, _12817_, _05271_);
  nor (_31291_, _31290_, _31286_);
  nor (_31292_, _31291_, _07778_);
  and (_31293_, _06298_, _05271_);
  nor (_31295_, _31293_, _31286_);
  and (_31296_, _31295_, _03601_);
  nor (_31297_, _05777_, _11154_);
  nor (_31298_, _31297_, _31286_);
  and (_31299_, _31298_, _07390_);
  and (_31300_, _05271_, \oc8051_golden_model_1.ACC [4]);
  nor (_31301_, _31300_, _31286_);
  nor (_31302_, _31301_, _03737_);
  nor (_31303_, _31301_, _09029_);
  nor (_31304_, _04409_, _31285_);
  or (_31306_, _31304_, _31303_);
  and (_31307_, _31306_, _04081_);
  nor (_31308_, _12841_, _11154_);
  nor (_31309_, _31308_, _31286_);
  nor (_31310_, _31309_, _04081_);
  or (_31311_, _31310_, _31307_);
  and (_31312_, _31311_, _03996_);
  nor (_31313_, _31298_, _03996_);
  nor (_31314_, _31313_, _31312_);
  nor (_31315_, _31314_, _03729_);
  or (_31317_, _31315_, _07390_);
  nor (_31318_, _31317_, _31302_);
  nor (_31319_, _31318_, _31299_);
  nor (_31320_, _31319_, _04481_);
  and (_31321_, _06730_, _05271_);
  nor (_31322_, _31286_, _07400_);
  not (_31323_, _31322_);
  nor (_31324_, _31323_, _31321_);
  or (_31325_, _31324_, _03222_);
  nor (_31326_, _31325_, _31320_);
  nor (_31328_, _12933_, _11154_);
  nor (_31329_, _31328_, _31286_);
  nor (_31330_, _31329_, _03589_);
  or (_31331_, _31330_, _03601_);
  nor (_31332_, _31331_, _31326_);
  nor (_31333_, _31332_, _31296_);
  or (_31334_, _31333_, _03600_);
  and (_31335_, _12821_, _05271_);
  or (_31336_, _31335_, _31286_);
  or (_31337_, _31336_, _07766_);
  and (_31339_, _31337_, _07778_);
  and (_31340_, _31339_, _31334_);
  nor (_31341_, _31340_, _31292_);
  nor (_31342_, _31341_, _03622_);
  nor (_31343_, _31286_, _05825_);
  not (_31344_, _31343_);
  nor (_31345_, _31295_, _07777_);
  and (_31346_, _31345_, _31344_);
  nor (_31347_, _31346_, _31342_);
  nor (_31348_, _31347_, _03790_);
  nor (_31350_, _31301_, _06828_);
  and (_31351_, _31350_, _31344_);
  nor (_31352_, _31351_, _03624_);
  not (_31353_, _31352_);
  nor (_31354_, _31353_, _31348_);
  nor (_31355_, _12819_, _11154_);
  or (_31356_, _31286_, _07795_);
  nor (_31357_, _31356_, _31355_);
  or (_31358_, _31357_, _03785_);
  nor (_31359_, _31358_, _31354_);
  nor (_31361_, _31359_, _31289_);
  nor (_31362_, _31361_, _03815_);
  nor (_31363_, _31309_, _04246_);
  or (_31364_, _31363_, _03447_);
  nor (_31365_, _31364_, _31362_);
  and (_31366_, _13003_, _05271_);
  or (_31367_, _31286_, _03514_);
  nor (_31368_, _31367_, _31366_);
  nor (_31369_, _31368_, _31365_);
  or (_31370_, _31369_, _43004_);
  or (_31372_, _43000_, \oc8051_golden_model_1.TL1 [4]);
  and (_31373_, _31372_, _41806_);
  and (_43653_, _31373_, _31370_);
  not (_31374_, \oc8051_golden_model_1.TL1 [5]);
  nor (_31375_, _05271_, _31374_);
  nor (_31376_, _13146_, _11154_);
  nor (_31377_, _31376_, _31375_);
  nor (_31378_, _31377_, _07793_);
  and (_31379_, _13147_, _05271_);
  nor (_31380_, _31379_, _31375_);
  nor (_31382_, _31380_, _07778_);
  and (_31383_, _06684_, _05271_);
  or (_31384_, _31383_, _31375_);
  and (_31385_, _31384_, _04481_);
  and (_31386_, _05271_, \oc8051_golden_model_1.ACC [5]);
  nor (_31387_, _31386_, _31375_);
  nor (_31388_, _31387_, _03737_);
  nor (_31389_, _31387_, _09029_);
  nor (_31390_, _04409_, _31374_);
  or (_31391_, _31390_, _31389_);
  and (_31393_, _31391_, _04081_);
  nor (_31394_, _13014_, _11154_);
  nor (_31395_, _31394_, _31375_);
  nor (_31396_, _31395_, _04081_);
  or (_31397_, _31396_, _31393_);
  and (_31398_, _31397_, _03996_);
  nor (_31399_, _05469_, _11154_);
  nor (_31400_, _31399_, _31375_);
  nor (_31401_, _31400_, _03996_);
  nor (_31402_, _31401_, _31398_);
  nor (_31404_, _31402_, _03729_);
  or (_31405_, _31404_, _07390_);
  nor (_31406_, _31405_, _31388_);
  and (_31407_, _31400_, _07390_);
  or (_31408_, _31407_, _04481_);
  nor (_31409_, _31408_, _31406_);
  or (_31410_, _31409_, _31385_);
  and (_31411_, _31410_, _03589_);
  nor (_31412_, _13127_, _11154_);
  nor (_31413_, _31412_, _31375_);
  nor (_31415_, _31413_, _03589_);
  or (_31416_, _31415_, _08828_);
  or (_31417_, _31416_, _31411_);
  and (_31418_, _13141_, _05271_);
  or (_31419_, _31375_, _07766_);
  or (_31420_, _31419_, _31418_);
  and (_31421_, _06306_, _05271_);
  nor (_31422_, _31421_, _31375_);
  and (_31423_, _31422_, _03601_);
  nor (_31424_, _31423_, _03780_);
  and (_31426_, _31424_, _31420_);
  and (_31427_, _31426_, _31417_);
  nor (_31428_, _31427_, _31382_);
  nor (_31429_, _31428_, _03622_);
  nor (_31430_, _31375_, _05518_);
  not (_31431_, _31430_);
  nor (_31432_, _31422_, _07777_);
  and (_31433_, _31432_, _31431_);
  nor (_31434_, _31433_, _31429_);
  nor (_31435_, _31434_, _03790_);
  nor (_31437_, _31387_, _06828_);
  and (_31438_, _31437_, _31431_);
  nor (_31439_, _31438_, _03624_);
  not (_31440_, _31439_);
  nor (_31441_, _31440_, _31435_);
  nor (_31442_, _13140_, _11154_);
  or (_31443_, _31375_, _07795_);
  nor (_31444_, _31443_, _31442_);
  or (_31445_, _31444_, _03785_);
  nor (_31446_, _31445_, _31441_);
  nor (_31448_, _31446_, _31378_);
  nor (_31449_, _31448_, _03815_);
  nor (_31450_, _31395_, _04246_);
  or (_31451_, _31450_, _03447_);
  nor (_31452_, _31451_, _31449_);
  and (_31453_, _13199_, _05271_);
  or (_31454_, _31375_, _03514_);
  nor (_31455_, _31454_, _31453_);
  nor (_31456_, _31455_, _31452_);
  or (_31457_, _31456_, _43004_);
  or (_31459_, _43000_, \oc8051_golden_model_1.TL1 [5]);
  and (_31460_, _31459_, _41806_);
  and (_43654_, _31460_, _31457_);
  not (_31461_, \oc8051_golden_model_1.TL1 [6]);
  nor (_31462_, _05271_, _31461_);
  nor (_31463_, _13352_, _11154_);
  nor (_31464_, _31463_, _31462_);
  nor (_31465_, _31464_, _07793_);
  and (_31466_, _13353_, _05271_);
  nor (_31467_, _31466_, _31462_);
  nor (_31469_, _31467_, _07778_);
  and (_31470_, _06455_, _05271_);
  or (_31471_, _31470_, _31462_);
  and (_31472_, _31471_, _04481_);
  and (_31473_, _05271_, \oc8051_golden_model_1.ACC [6]);
  nor (_31474_, _31473_, _31462_);
  nor (_31475_, _31474_, _03737_);
  nor (_31476_, _31474_, _09029_);
  nor (_31477_, _04409_, _31461_);
  or (_31478_, _31477_, _31476_);
  and (_31480_, _31478_, _04081_);
  nor (_31481_, _13242_, _11154_);
  nor (_31482_, _31481_, _31462_);
  nor (_31483_, _31482_, _04081_);
  or (_31484_, _31483_, _31480_);
  and (_31485_, _31484_, _03996_);
  nor (_31486_, _05363_, _11154_);
  nor (_31487_, _31486_, _31462_);
  nor (_31488_, _31487_, _03996_);
  nor (_31489_, _31488_, _31485_);
  nor (_31491_, _31489_, _03729_);
  or (_31492_, _31491_, _07390_);
  nor (_31493_, _31492_, _31475_);
  and (_31494_, _31487_, _07390_);
  or (_31495_, _31494_, _04481_);
  nor (_31496_, _31495_, _31493_);
  or (_31497_, _31496_, _31472_);
  and (_31498_, _31497_, _03589_);
  nor (_31499_, _13332_, _11154_);
  nor (_31500_, _31499_, _31462_);
  nor (_31502_, _31500_, _03589_);
  or (_31503_, _31502_, _08828_);
  or (_31504_, _31503_, _31498_);
  and (_31505_, _13347_, _05271_);
  or (_31506_, _31462_, _07766_);
  or (_31507_, _31506_, _31505_);
  and (_31508_, _13339_, _05271_);
  nor (_31509_, _31508_, _31462_);
  and (_31510_, _31509_, _03601_);
  nor (_31511_, _31510_, _03780_);
  and (_31513_, _31511_, _31507_);
  and (_31514_, _31513_, _31504_);
  nor (_31515_, _31514_, _31469_);
  nor (_31516_, _31515_, _03622_);
  nor (_31517_, _31462_, _05412_);
  not (_31518_, _31517_);
  nor (_31519_, _31509_, _07777_);
  and (_31520_, _31519_, _31518_);
  nor (_31521_, _31520_, _31516_);
  nor (_31522_, _31521_, _03790_);
  nor (_31524_, _31474_, _06828_);
  and (_31525_, _31524_, _31518_);
  or (_31526_, _31525_, _31522_);
  and (_31527_, _31526_, _07795_);
  nor (_31528_, _13346_, _11154_);
  nor (_31529_, _31528_, _31462_);
  nor (_31530_, _31529_, _07795_);
  or (_31531_, _31530_, _31527_);
  and (_31532_, _31531_, _07793_);
  nor (_31533_, _31532_, _31465_);
  nor (_31535_, _31533_, _03815_);
  nor (_31536_, _31482_, _04246_);
  or (_31537_, _31536_, _03447_);
  nor (_31538_, _31537_, _31535_);
  and (_31539_, _13402_, _05271_);
  or (_31540_, _31462_, _03514_);
  nor (_31541_, _31540_, _31539_);
  nor (_31542_, _31541_, _31538_);
  or (_31543_, _31542_, _43004_);
  or (_31544_, _43000_, \oc8051_golden_model_1.TL1 [6]);
  and (_31546_, _31544_, _41806_);
  and (_43655_, _31546_, _31543_);
  not (_31547_, \oc8051_golden_model_1.TMOD [0]);
  nor (_31548_, _05286_, _31547_);
  nor (_31549_, _05666_, _11236_);
  nor (_31550_, _31549_, _31548_);
  and (_31551_, _31550_, _17166_);
  and (_31552_, _05286_, \oc8051_golden_model_1.ACC [0]);
  nor (_31553_, _31552_, _31548_);
  nor (_31554_, _31553_, _03737_);
  nor (_31555_, _31553_, _09029_);
  nor (_31556_, _04409_, _31547_);
  or (_31557_, _31556_, _31555_);
  and (_31558_, _31557_, _04081_);
  nor (_31559_, _31550_, _04081_);
  or (_31560_, _31559_, _31558_);
  and (_31561_, _31560_, _03996_);
  and (_31562_, _05286_, _04620_);
  nor (_31563_, _31562_, _31548_);
  nor (_31564_, _31563_, _03996_);
  nor (_31566_, _31564_, _31561_);
  nor (_31567_, _31566_, _03729_);
  or (_31568_, _31567_, _07390_);
  nor (_31569_, _31568_, _31554_);
  and (_31570_, _31563_, _07390_);
  nor (_31571_, _31570_, _31569_);
  nor (_31572_, _31571_, _04481_);
  and (_31573_, _06546_, _05286_);
  nor (_31574_, _31548_, _07400_);
  not (_31575_, _31574_);
  nor (_31577_, _31575_, _31573_);
  nor (_31578_, _31577_, _31572_);
  nor (_31579_, _31578_, _03222_);
  nor (_31580_, _12109_, _11236_);
  or (_31581_, _31548_, _03589_);
  nor (_31582_, _31581_, _31580_);
  or (_31583_, _31582_, _03601_);
  nor (_31584_, _31583_, _31579_);
  and (_31585_, _05286_, _06274_);
  nor (_31586_, _31585_, _31548_);
  nor (_31588_, _31586_, _05886_);
  or (_31589_, _31588_, _31584_);
  and (_31590_, _31589_, _07766_);
  and (_31591_, _12124_, _05286_);
  nor (_31592_, _31591_, _31548_);
  nor (_31593_, _31592_, _07766_);
  or (_31594_, _31593_, _31590_);
  nor (_31595_, _31594_, _03780_);
  and (_31596_, _12128_, _05286_);
  or (_31597_, _31548_, _07778_);
  nor (_31599_, _31597_, _31596_);
  or (_31600_, _31599_, _03622_);
  nor (_31601_, _31600_, _31595_);
  or (_31602_, _31586_, _07777_);
  nor (_31603_, _31602_, _31549_);
  nor (_31604_, _31603_, _31601_);
  nor (_31605_, _31604_, _03790_);
  and (_31606_, _12005_, _05286_);
  or (_31607_, _31606_, _31548_);
  and (_31608_, _31607_, _03790_);
  or (_31610_, _31608_, _31605_);
  and (_31611_, _31610_, _07795_);
  nor (_31612_, _12122_, _11236_);
  nor (_31613_, _31612_, _31548_);
  nor (_31614_, _31613_, _07795_);
  or (_31615_, _31614_, _31611_);
  and (_31616_, _31615_, _07793_);
  nor (_31617_, _12003_, _11236_);
  nor (_31618_, _31617_, _31548_);
  nor (_31619_, _31618_, _07793_);
  nor (_31621_, _31619_, _17166_);
  not (_31622_, _31621_);
  nor (_31623_, _31622_, _31616_);
  nor (_31624_, _31623_, _31551_);
  or (_31625_, _31624_, _43004_);
  or (_31626_, _43000_, \oc8051_golden_model_1.TMOD [0]);
  and (_31627_, _31626_, _41806_);
  and (_43658_, _31627_, _31625_);
  and (_31628_, _06501_, _05286_);
  not (_31629_, \oc8051_golden_model_1.TMOD [1]);
  nor (_31631_, _05286_, _31629_);
  nor (_31632_, _31631_, _07400_);
  not (_31633_, _31632_);
  nor (_31634_, _31633_, _31628_);
  not (_31635_, _31634_);
  and (_31636_, _05286_, _06764_);
  nor (_31637_, _31636_, _31631_);
  and (_31638_, _31637_, _07390_);
  nor (_31639_, _05286_, \oc8051_golden_model_1.TMOD [1]);
  and (_31640_, _05286_, _03274_);
  nor (_31642_, _31640_, _31639_);
  and (_31643_, _31642_, _03729_);
  and (_31644_, _31642_, _04409_);
  nor (_31645_, _04409_, _31629_);
  or (_31646_, _31645_, _31644_);
  and (_31647_, _31646_, _04081_);
  and (_31648_, _12213_, _05286_);
  nor (_31649_, _31648_, _31639_);
  and (_31650_, _31649_, _03610_);
  or (_31651_, _31650_, _31647_);
  and (_31653_, _31651_, _03996_);
  nor (_31654_, _31637_, _03996_);
  nor (_31655_, _31654_, _31653_);
  nor (_31656_, _31655_, _03729_);
  or (_31657_, _31656_, _07390_);
  nor (_31658_, _31657_, _31643_);
  nor (_31659_, _31658_, _31638_);
  nor (_31660_, _31659_, _04481_);
  nor (_31661_, _31660_, _03222_);
  and (_31662_, _31661_, _31635_);
  not (_31664_, _31639_);
  and (_31665_, _12313_, _05286_);
  nor (_31666_, _31665_, _03589_);
  and (_31667_, _31666_, _31664_);
  nor (_31668_, _31667_, _31662_);
  nor (_31669_, _31668_, _08828_);
  nor (_31670_, _12327_, _11236_);
  nor (_31671_, _31670_, _07766_);
  and (_31672_, _05286_, _04303_);
  nor (_31673_, _31672_, _05886_);
  nor (_31675_, _31673_, _31671_);
  nor (_31676_, _31675_, _31639_);
  nor (_31677_, _31676_, _31669_);
  nor (_31678_, _31677_, _03780_);
  nor (_31679_, _12333_, _11236_);
  nor (_31680_, _31679_, _07778_);
  and (_31681_, _31680_, _31664_);
  nor (_31682_, _31681_, _31678_);
  nor (_31683_, _31682_, _03622_);
  nor (_31684_, _12207_, _11236_);
  nor (_31685_, _31684_, _07777_);
  and (_31686_, _31685_, _31664_);
  nor (_31687_, _31686_, _31683_);
  nor (_31688_, _31687_, _03790_);
  nor (_31689_, _31631_, _05618_);
  nor (_31690_, _31689_, _06828_);
  and (_31691_, _31690_, _31642_);
  nor (_31692_, _31691_, _31688_);
  or (_31693_, _31692_, _18499_);
  and (_31694_, _31672_, _05617_);
  nor (_31697_, _31694_, _07795_);
  and (_31698_, _31697_, _31664_);
  nand (_31699_, _31640_, _05617_);
  nor (_31700_, _31639_, _07793_);
  and (_31701_, _31700_, _31699_);
  or (_31702_, _31701_, _03815_);
  nor (_31703_, _31702_, _31698_);
  and (_31704_, _31703_, _31693_);
  nor (_31705_, _31649_, _04246_);
  nor (_31706_, _31705_, _31704_);
  and (_31708_, _31706_, _03514_);
  nor (_31709_, _31648_, _31631_);
  nor (_31710_, _31709_, _03514_);
  or (_31711_, _31710_, _31708_);
  or (_31712_, _31711_, _43004_);
  or (_31713_, _43000_, \oc8051_golden_model_1.TMOD [1]);
  and (_31714_, _31713_, _41806_);
  and (_43659_, _31714_, _31712_);
  not (_31715_, \oc8051_golden_model_1.TMOD [2]);
  nor (_31716_, _05286_, _31715_);
  nor (_31718_, _12538_, _11236_);
  nor (_31719_, _31718_, _31716_);
  nor (_31720_, _31719_, _07793_);
  and (_31721_, _12539_, _05286_);
  nor (_31722_, _31721_, _31716_);
  nor (_31723_, _31722_, _07778_);
  and (_31724_, _05286_, \oc8051_golden_model_1.ACC [2]);
  nor (_31725_, _31724_, _31716_);
  nor (_31726_, _31725_, _03737_);
  nor (_31727_, _31725_, _09029_);
  nor (_31729_, _04409_, _31715_);
  or (_31730_, _31729_, _31727_);
  and (_31731_, _31730_, _04081_);
  nor (_31732_, _12416_, _11236_);
  nor (_31733_, _31732_, _31716_);
  nor (_31734_, _31733_, _04081_);
  or (_31735_, _31734_, _31731_);
  and (_31736_, _31735_, _03996_);
  nor (_31737_, _11236_, _04875_);
  nor (_31738_, _31737_, _31716_);
  nor (_31740_, _31738_, _03996_);
  nor (_31741_, _31740_, _31736_);
  nor (_31742_, _31741_, _03729_);
  or (_31743_, _31742_, _07390_);
  nor (_31744_, _31743_, _31726_);
  and (_31745_, _31738_, _07390_);
  nor (_31746_, _31745_, _31744_);
  nor (_31747_, _31746_, _04481_);
  and (_31748_, _06637_, _05286_);
  nor (_31749_, _31716_, _07400_);
  not (_31751_, _31749_);
  nor (_31752_, _31751_, _31748_);
  nor (_31753_, _31752_, _03222_);
  not (_31754_, _31753_);
  nor (_31755_, _31754_, _31747_);
  nor (_31756_, _12519_, _11236_);
  nor (_31757_, _31756_, _31716_);
  nor (_31758_, _31757_, _03589_);
  or (_31759_, _31758_, _08828_);
  or (_31760_, _31759_, _31755_);
  and (_31762_, _12533_, _05286_);
  or (_31763_, _31716_, _07766_);
  or (_31764_, _31763_, _31762_);
  and (_31765_, _05286_, _06332_);
  nor (_31766_, _31765_, _31716_);
  and (_31767_, _31766_, _03601_);
  nor (_31768_, _31767_, _03780_);
  and (_31769_, _31768_, _31764_);
  and (_31770_, _31769_, _31760_);
  nor (_31771_, _31770_, _31723_);
  nor (_31773_, _31771_, _03622_);
  nor (_31774_, _31716_, _05718_);
  not (_31775_, _31774_);
  nor (_31776_, _31766_, _07777_);
  and (_31777_, _31776_, _31775_);
  nor (_31778_, _31777_, _31773_);
  nor (_31779_, _31778_, _03790_);
  nor (_31780_, _31725_, _06828_);
  and (_31781_, _31780_, _31775_);
  nor (_31782_, _31781_, _03624_);
  not (_31784_, _31782_);
  nor (_31785_, _31784_, _31779_);
  nor (_31786_, _12532_, _11236_);
  or (_31787_, _31716_, _07795_);
  nor (_31788_, _31787_, _31786_);
  or (_31789_, _31788_, _03785_);
  nor (_31790_, _31789_, _31785_);
  nor (_31791_, _31790_, _31720_);
  nor (_31792_, _31791_, _03815_);
  nor (_31793_, _31733_, _04246_);
  or (_31795_, _31793_, _03447_);
  nor (_31796_, _31795_, _31792_);
  and (_31797_, _12592_, _05286_);
  or (_31798_, _31716_, _03514_);
  nor (_31799_, _31798_, _31797_);
  nor (_31800_, _31799_, _31796_);
  or (_31801_, _31800_, _43004_);
  or (_31802_, _43000_, \oc8051_golden_model_1.TMOD [2]);
  and (_31803_, _31802_, _41806_);
  and (_43660_, _31803_, _31801_);
  not (_31805_, \oc8051_golden_model_1.TMOD [3]);
  nor (_31806_, _05286_, _31805_);
  nor (_31807_, _12738_, _11236_);
  nor (_31808_, _31807_, _31806_);
  nor (_31809_, _31808_, _07793_);
  and (_31810_, _12739_, _05286_);
  nor (_31811_, _31810_, _31806_);
  nor (_31812_, _31811_, _07778_);
  and (_31813_, _06592_, _05286_);
  or (_31814_, _31813_, _31806_);
  and (_31816_, _31814_, _04481_);
  and (_31817_, _05286_, \oc8051_golden_model_1.ACC [3]);
  nor (_31818_, _31817_, _31806_);
  nor (_31819_, _31818_, _03737_);
  nor (_31820_, _31818_, _09029_);
  nor (_31821_, _04409_, _31805_);
  or (_31822_, _31821_, _31820_);
  and (_31823_, _31822_, _04081_);
  nor (_31824_, _12627_, _11236_);
  nor (_31825_, _31824_, _31806_);
  nor (_31827_, _31825_, _04081_);
  or (_31828_, _31827_, _31823_);
  and (_31829_, _31828_, _03996_);
  nor (_31830_, _11236_, _05005_);
  nor (_31831_, _31830_, _31806_);
  nor (_31832_, _31831_, _03996_);
  nor (_31833_, _31832_, _31829_);
  nor (_31834_, _31833_, _03729_);
  or (_31835_, _31834_, _07390_);
  nor (_31836_, _31835_, _31819_);
  and (_31838_, _31831_, _07390_);
  or (_31839_, _31838_, _04481_);
  nor (_31840_, _31839_, _31836_);
  or (_31841_, _31840_, _31816_);
  and (_31842_, _31841_, _03589_);
  nor (_31843_, _12718_, _11236_);
  nor (_31844_, _31843_, _31806_);
  nor (_31845_, _31844_, _03589_);
  or (_31846_, _31845_, _08828_);
  or (_31847_, _31846_, _31842_);
  and (_31849_, _12733_, _05286_);
  or (_31850_, _31806_, _07766_);
  or (_31851_, _31850_, _31849_);
  and (_31852_, _05286_, _06276_);
  nor (_31853_, _31852_, _31806_);
  and (_31854_, _31853_, _03601_);
  nor (_31855_, _31854_, _03780_);
  and (_31856_, _31855_, _31851_);
  and (_31857_, _31856_, _31847_);
  nor (_31858_, _31857_, _31812_);
  nor (_31860_, _31858_, _03622_);
  nor (_31861_, _31806_, _05567_);
  not (_31862_, _31861_);
  nor (_31863_, _31853_, _07777_);
  and (_31864_, _31863_, _31862_);
  nor (_31865_, _31864_, _31860_);
  nor (_31866_, _31865_, _03790_);
  nor (_31867_, _31818_, _06828_);
  and (_31868_, _31867_, _31862_);
  or (_31869_, _31868_, _31866_);
  and (_31871_, _31869_, _07795_);
  nor (_31872_, _12732_, _11236_);
  nor (_31873_, _31872_, _31806_);
  nor (_31874_, _31873_, _07795_);
  or (_31875_, _31874_, _31871_);
  and (_31876_, _31875_, _07793_);
  nor (_31877_, _31876_, _31809_);
  nor (_31878_, _31877_, _03815_);
  nor (_31879_, _31825_, _04246_);
  or (_31880_, _31879_, _03447_);
  nor (_31882_, _31880_, _31878_);
  and (_31883_, _12794_, _05286_);
  or (_31884_, _31806_, _03514_);
  nor (_31885_, _31884_, _31883_);
  nor (_31886_, _31885_, _31882_);
  or (_31887_, _31886_, _43004_);
  or (_31888_, _43000_, \oc8051_golden_model_1.TMOD [3]);
  and (_31889_, _31888_, _41806_);
  and (_43663_, _31889_, _31887_);
  not (_31890_, \oc8051_golden_model_1.TMOD [4]);
  nor (_31892_, _05286_, _31890_);
  nor (_31893_, _12816_, _11236_);
  nor (_31894_, _31893_, _31892_);
  nor (_31895_, _31894_, _07793_);
  and (_31896_, _12817_, _05286_);
  nor (_31897_, _31896_, _31892_);
  nor (_31898_, _31897_, _07778_);
  and (_31899_, _06298_, _05286_);
  nor (_31900_, _31899_, _31892_);
  and (_31901_, _31900_, _03601_);
  and (_31903_, _05286_, \oc8051_golden_model_1.ACC [4]);
  nor (_31904_, _31903_, _31892_);
  nor (_31905_, _31904_, _03737_);
  nor (_31906_, _31904_, _09029_);
  nor (_31907_, _04409_, _31890_);
  or (_31908_, _31907_, _31906_);
  and (_31909_, _31908_, _04081_);
  nor (_31910_, _12841_, _11236_);
  nor (_31911_, _31910_, _31892_);
  nor (_31912_, _31911_, _04081_);
  or (_31914_, _31912_, _31909_);
  and (_31915_, _31914_, _03996_);
  nor (_31916_, _05777_, _11236_);
  nor (_31917_, _31916_, _31892_);
  nor (_31918_, _31917_, _03996_);
  nor (_31919_, _31918_, _31915_);
  nor (_31920_, _31919_, _03729_);
  or (_31921_, _31920_, _07390_);
  nor (_31922_, _31921_, _31905_);
  and (_31923_, _31917_, _07390_);
  nor (_31925_, _31923_, _31922_);
  nor (_31926_, _31925_, _04481_);
  and (_31927_, _06730_, _05286_);
  nor (_31928_, _31892_, _07400_);
  not (_31929_, _31928_);
  nor (_31930_, _31929_, _31927_);
  or (_31931_, _31930_, _03222_);
  nor (_31932_, _31931_, _31926_);
  nor (_31933_, _12933_, _11236_);
  nor (_31934_, _31933_, _31892_);
  nor (_31936_, _31934_, _03589_);
  or (_31937_, _31936_, _03601_);
  nor (_31938_, _31937_, _31932_);
  nor (_31939_, _31938_, _31901_);
  or (_31940_, _31939_, _03600_);
  and (_31941_, _12821_, _05286_);
  or (_31942_, _31941_, _31892_);
  or (_31943_, _31942_, _07766_);
  and (_31944_, _31943_, _07778_);
  and (_31945_, _31944_, _31940_);
  nor (_31947_, _31945_, _31898_);
  nor (_31948_, _31947_, _03622_);
  nor (_31949_, _31892_, _05825_);
  not (_31950_, _31949_);
  nor (_31951_, _31900_, _07777_);
  and (_31952_, _31951_, _31950_);
  nor (_31953_, _31952_, _31948_);
  nor (_31954_, _31953_, _03790_);
  nor (_31955_, _31904_, _06828_);
  and (_31956_, _31955_, _31950_);
  nor (_31958_, _31956_, _03624_);
  not (_31959_, _31958_);
  nor (_31960_, _31959_, _31954_);
  nor (_31961_, _12819_, _11236_);
  or (_31962_, _31892_, _07795_);
  nor (_31963_, _31962_, _31961_);
  or (_31964_, _31963_, _03785_);
  nor (_31965_, _31964_, _31960_);
  nor (_31966_, _31965_, _31895_);
  nor (_31967_, _31966_, _03815_);
  nor (_31969_, _31911_, _04246_);
  or (_31970_, _31969_, _03447_);
  nor (_31971_, _31970_, _31967_);
  and (_31972_, _13003_, _05286_);
  or (_31973_, _31892_, _03514_);
  nor (_31974_, _31973_, _31972_);
  nor (_31975_, _31974_, _31971_);
  or (_31976_, _31975_, _43004_);
  or (_31977_, _43000_, \oc8051_golden_model_1.TMOD [4]);
  and (_31978_, _31977_, _41806_);
  and (_43664_, _31978_, _31976_);
  not (_31980_, \oc8051_golden_model_1.TMOD [5]);
  nor (_31981_, _05286_, _31980_);
  nor (_31982_, _13146_, _11236_);
  nor (_31983_, _31982_, _31981_);
  nor (_31984_, _31983_, _07793_);
  and (_31985_, _13147_, _05286_);
  nor (_31986_, _31985_, _31981_);
  nor (_31987_, _31986_, _07778_);
  and (_31988_, _06684_, _05286_);
  or (_31990_, _31988_, _31981_);
  and (_31991_, _31990_, _04481_);
  and (_31992_, _05286_, \oc8051_golden_model_1.ACC [5]);
  nor (_31993_, _31992_, _31981_);
  nor (_31994_, _31993_, _03737_);
  nor (_31995_, _31993_, _09029_);
  nor (_31996_, _04409_, _31980_);
  or (_31997_, _31996_, _31995_);
  and (_31998_, _31997_, _04081_);
  nor (_31999_, _13014_, _11236_);
  nor (_32001_, _31999_, _31981_);
  nor (_32002_, _32001_, _04081_);
  or (_32003_, _32002_, _31998_);
  and (_32004_, _32003_, _03996_);
  nor (_32005_, _05469_, _11236_);
  nor (_32006_, _32005_, _31981_);
  nor (_32007_, _32006_, _03996_);
  nor (_32008_, _32007_, _32004_);
  nor (_32009_, _32008_, _03729_);
  or (_32010_, _32009_, _07390_);
  nor (_32012_, _32010_, _31994_);
  and (_32013_, _32006_, _07390_);
  or (_32014_, _32013_, _04481_);
  nor (_32015_, _32014_, _32012_);
  or (_32016_, _32015_, _31991_);
  and (_32017_, _32016_, _03589_);
  nor (_32018_, _13127_, _11236_);
  nor (_32019_, _32018_, _31981_);
  nor (_32020_, _32019_, _03589_);
  or (_32021_, _32020_, _08828_);
  or (_32023_, _32021_, _32017_);
  and (_32024_, _13141_, _05286_);
  or (_32025_, _31981_, _07766_);
  or (_32026_, _32025_, _32024_);
  and (_32027_, _06306_, _05286_);
  nor (_32028_, _32027_, _31981_);
  and (_32029_, _32028_, _03601_);
  nor (_32030_, _32029_, _03780_);
  and (_32031_, _32030_, _32026_);
  and (_32032_, _32031_, _32023_);
  nor (_32034_, _32032_, _31987_);
  nor (_32035_, _32034_, _03622_);
  nor (_32036_, _31981_, _05518_);
  not (_32037_, _32036_);
  nor (_32038_, _32028_, _07777_);
  and (_32039_, _32038_, _32037_);
  nor (_32040_, _32039_, _32035_);
  nor (_32041_, _32040_, _03790_);
  nor (_32042_, _31993_, _06828_);
  and (_32043_, _32042_, _32037_);
  or (_32045_, _32043_, _32041_);
  and (_32046_, _32045_, _07795_);
  nor (_32047_, _13140_, _11236_);
  nor (_32048_, _32047_, _31981_);
  nor (_32049_, _32048_, _07795_);
  or (_32050_, _32049_, _32046_);
  and (_32051_, _32050_, _07793_);
  nor (_32052_, _32051_, _31984_);
  nor (_32053_, _32052_, _03815_);
  nor (_32054_, _32001_, _04246_);
  or (_32056_, _32054_, _03447_);
  nor (_32057_, _32056_, _32053_);
  and (_32058_, _13199_, _05286_);
  or (_32059_, _31981_, _03514_);
  nor (_32060_, _32059_, _32058_);
  nor (_32061_, _32060_, _32057_);
  or (_32062_, _32061_, _43004_);
  or (_32063_, _43000_, \oc8051_golden_model_1.TMOD [5]);
  and (_32064_, _32063_, _41806_);
  and (_43665_, _32064_, _32062_);
  not (_32066_, \oc8051_golden_model_1.TMOD [6]);
  nor (_32067_, _05286_, _32066_);
  nor (_32068_, _13352_, _11236_);
  nor (_32069_, _32068_, _32067_);
  nor (_32070_, _32069_, _07793_);
  and (_32071_, _13353_, _05286_);
  nor (_32072_, _32071_, _32067_);
  nor (_32073_, _32072_, _07778_);
  and (_32074_, _06455_, _05286_);
  or (_32075_, _32074_, _32067_);
  and (_32077_, _32075_, _04481_);
  and (_32078_, _05286_, \oc8051_golden_model_1.ACC [6]);
  nor (_32079_, _32078_, _32067_);
  nor (_32080_, _32079_, _03737_);
  nor (_32081_, _32079_, _09029_);
  nor (_32082_, _04409_, _32066_);
  or (_32083_, _32082_, _32081_);
  and (_32084_, _32083_, _04081_);
  nor (_32085_, _13242_, _11236_);
  nor (_32086_, _32085_, _32067_);
  nor (_32088_, _32086_, _04081_);
  or (_32089_, _32088_, _32084_);
  and (_32090_, _32089_, _03996_);
  nor (_32091_, _05363_, _11236_);
  nor (_32092_, _32091_, _32067_);
  nor (_32093_, _32092_, _03996_);
  nor (_32094_, _32093_, _32090_);
  nor (_32095_, _32094_, _03729_);
  or (_32096_, _32095_, _07390_);
  nor (_32097_, _32096_, _32080_);
  and (_32099_, _32092_, _07390_);
  or (_32100_, _32099_, _04481_);
  nor (_32101_, _32100_, _32097_);
  or (_32102_, _32101_, _32077_);
  and (_32103_, _32102_, _03589_);
  nor (_32104_, _13332_, _11236_);
  nor (_32105_, _32104_, _32067_);
  nor (_32106_, _32105_, _03589_);
  or (_32107_, _32106_, _08828_);
  or (_32108_, _32107_, _32103_);
  and (_32110_, _13347_, _05286_);
  or (_32111_, _32067_, _07766_);
  or (_32112_, _32111_, _32110_);
  and (_32113_, _13339_, _05286_);
  nor (_32114_, _32113_, _32067_);
  and (_32115_, _32114_, _03601_);
  nor (_32116_, _32115_, _03780_);
  and (_32117_, _32116_, _32112_);
  and (_32118_, _32117_, _32108_);
  nor (_32119_, _32118_, _32073_);
  nor (_32121_, _32119_, _03622_);
  nor (_32122_, _32067_, _05412_);
  not (_32123_, _32122_);
  nor (_32124_, _32114_, _07777_);
  and (_32125_, _32124_, _32123_);
  nor (_32126_, _32125_, _32121_);
  nor (_32127_, _32126_, _03790_);
  nor (_32128_, _32079_, _06828_);
  and (_32129_, _32128_, _32123_);
  or (_32130_, _32129_, _32127_);
  and (_32132_, _32130_, _07795_);
  nor (_32133_, _13346_, _11236_);
  nor (_32134_, _32133_, _32067_);
  nor (_32135_, _32134_, _07795_);
  or (_32136_, _32135_, _32132_);
  and (_32137_, _32136_, _07793_);
  nor (_32138_, _32137_, _32070_);
  nor (_32139_, _32138_, _03815_);
  nor (_32140_, _32086_, _04246_);
  or (_32141_, _32140_, _03447_);
  nor (_32143_, _32141_, _32139_);
  and (_32144_, _13402_, _05286_);
  or (_32145_, _32067_, _03514_);
  nor (_32146_, _32145_, _32144_);
  nor (_32147_, _32146_, _32143_);
  or (_32148_, _32147_, _43004_);
  or (_32149_, _43000_, \oc8051_golden_model_1.TMOD [6]);
  and (_32150_, _32149_, _41806_);
  and (_43666_, _32150_, _32148_);
  and (_32151_, _11975_, _02905_);
  nor (_32153_, _03631_, _03196_);
  not (_32154_, _32153_);
  and (_32155_, _32154_, _04163_);
  and (_32156_, _09854_, \oc8051_golden_model_1.PC [0]);
  and (_32157_, _04163_, \oc8051_golden_model_1.PC [0]);
  nor (_32158_, _32157_, _11444_);
  nor (_32159_, _32158_, _09854_);
  nor (_32160_, _32159_, _32156_);
  and (_32161_, _32160_, _03453_);
  and (_32162_, _11933_, _11940_);
  nor (_32164_, _32162_, _02905_);
  not (_32165_, _03203_);
  and (_32166_, _11328_, _08733_);
  nor (_32167_, _32166_, _02905_);
  not (_32168_, _03201_);
  and (_32169_, _11335_, _07795_);
  nor (_32170_, _32169_, _02905_);
  not (_32171_, _03192_);
  and (_32172_, _11851_, _07777_);
  nor (_32173_, _32172_, _02905_);
  not (_32175_, _03182_);
  and (_32176_, _11345_, _07766_);
  nor (_32177_, _32176_, _02905_);
  and (_32178_, _03601_, _02905_);
  nor (_32179_, _03625_, _03222_);
  and (_32180_, _32179_, _11756_);
  nor (_32181_, _32180_, _02905_);
  nor (_32182_, _04163_, _03227_);
  nor (_32183_, _04163_, _03233_);
  and (_32184_, _04163_, _03980_);
  nor (_32186_, _11630_, _02905_);
  nor (_32187_, _11642_, _02905_);
  and (_32188_, _11642_, _02905_);
  nor (_32189_, _32188_, _32187_);
  and (_32190_, _11630_, _04763_);
  not (_32191_, _32190_);
  nor (_32192_, _32191_, _32189_);
  nor (_32193_, _32192_, _32186_);
  not (_32194_, _32193_);
  nor (_32195_, _32194_, _32184_);
  nor (_32197_, _32195_, _06073_);
  and (_32198_, _11504_, \oc8051_golden_model_1.PC [0]);
  and (_32199_, _04048_, _02905_);
  nor (_32200_, _32199_, _11571_);
  and (_32201_, _32200_, _11624_);
  or (_32202_, _32201_, _32198_);
  nor (_32203_, _32202_, _06072_);
  nor (_32204_, _32203_, _32197_);
  nor (_32205_, _32204_, _04422_);
  and (_32206_, _04422_, \oc8051_golden_model_1.PC [0]);
  nor (_32208_, _32206_, _03610_);
  not (_32209_, _32208_);
  nor (_32210_, _32209_, _32205_);
  not (_32211_, _32210_);
  not (_32212_, _32158_);
  and (_32213_, _32212_, _11367_);
  and (_32214_, _05666_, _05566_);
  and (_32215_, _32214_, _11366_);
  nand (_32216_, _32215_, _12413_);
  nor (_32217_, _32216_, _02905_);
  or (_32219_, _32217_, _04081_);
  or (_32220_, _32219_, _32213_);
  and (_32221_, _32220_, _11362_);
  and (_32222_, _32221_, _32211_);
  nor (_32223_, _11362_, _02905_);
  nor (_32224_, _32223_, _04768_);
  not (_32225_, _32224_);
  nor (_32226_, _32225_, _32222_);
  nor (_32227_, _04163_, _03230_);
  and (_32228_, _11666_, _11659_);
  not (_32230_, _32228_);
  nor (_32231_, _32230_, _32227_);
  not (_32232_, _32231_);
  nor (_32233_, _32232_, _32226_);
  nor (_32234_, _32228_, _02905_);
  nor (_32235_, _32234_, _11670_);
  not (_32236_, _32235_);
  nor (_32237_, _32236_, _32233_);
  or (_32238_, _32237_, _09917_);
  nor (_32239_, _32238_, _32183_);
  and (_32241_, _09969_, _02905_);
  not (_32242_, _32241_);
  nor (_32243_, _32212_, _09969_);
  nor (_32244_, _32243_, _09921_);
  and (_32245_, _32244_, _32242_);
  or (_32246_, _32245_, _03615_);
  or (_32247_, _32246_, _32239_);
  and (_32248_, _32247_, _09920_);
  and (_32249_, _11685_, _02905_);
  and (_32250_, _32158_, _10018_);
  or (_32252_, _32250_, _32249_);
  nor (_32253_, _32252_, _09920_);
  nor (_32254_, _32253_, _32248_);
  and (_32255_, _09876_, _02905_);
  nor (_32256_, _32212_, _09876_);
  nor (_32257_, _32256_, _32255_);
  nor (_32258_, _32257_, _04107_);
  nor (_32259_, _32258_, _32254_);
  nor (_32260_, _32259_, _03604_);
  and (_32261_, _10061_, _02905_);
  nor (_32263_, _32212_, _10061_);
  or (_32264_, _32263_, _32261_);
  and (_32265_, _32264_, _03604_);
  or (_32266_, _32265_, _32260_);
  and (_32267_, _32266_, _11358_);
  and (_32268_, _10025_, _02905_);
  or (_32269_, _32268_, _32267_);
  and (_32270_, _32269_, _03227_);
  or (_32271_, _32270_, _11356_);
  nor (_32272_, _32271_, _32182_);
  nor (_32274_, _11355_, _02905_);
  nor (_32275_, _32274_, _11727_);
  not (_32276_, _32275_);
  nor (_32277_, _32276_, _32272_);
  nor (_32278_, _04163_, _03238_);
  and (_32279_, _11350_, _03248_);
  not (_32280_, _32279_);
  nor (_32281_, _32280_, _32278_);
  not (_32282_, _32281_);
  nor (_32283_, _32282_, _32277_);
  nor (_32284_, _32279_, _02905_);
  nor (_32285_, _32284_, _03224_);
  not (_32286_, _32285_);
  nor (_32287_, _32286_, _32283_);
  nor (_32288_, _04163_, _05897_);
  not (_32289_, _32180_);
  nor (_32290_, _32289_, _32288_);
  not (_32291_, _32290_);
  nor (_32292_, _32291_, _32287_);
  or (_32293_, _32292_, _03169_);
  nor (_32295_, _32293_, _32181_);
  nor (_32296_, _04163_, _03170_);
  or (_32297_, _32296_, _11764_);
  or (_32298_, _32297_, _32295_);
  or (_32299_, _32200_, _11765_);
  and (_32300_, _32299_, _32298_);
  and (_32301_, _32300_, _05886_);
  or (_32302_, _32301_, _32178_);
  and (_32303_, _32302_, _11348_);
  and (_32304_, _11347_, _03329_);
  or (_32306_, _32304_, _32303_);
  and (_32307_, _32306_, _10736_);
  nor (_32308_, _04163_, _10736_);
  or (_32309_, _32308_, _32307_);
  and (_32310_, _32309_, _11820_);
  not (_32311_, _32176_);
  and (_32312_, _08786_, \oc8051_golden_model_1.PC [0]);
  and (_32313_, _32200_, _11826_);
  or (_32314_, _32313_, _32312_);
  and (_32315_, _32314_, _11819_);
  nor (_32316_, _32315_, _32311_);
  not (_32317_, _32316_);
  nor (_32318_, _32317_, _32310_);
  nor (_32319_, _32318_, _32177_);
  and (_32320_, _32319_, _32175_);
  nor (_32321_, _04163_, _32175_);
  or (_32322_, _32321_, _32320_);
  and (_32323_, _32322_, _11842_);
  not (_32324_, _32172_);
  nor (_32325_, _32200_, _11826_);
  nor (_32328_, _08786_, \oc8051_golden_model_1.PC [0]);
  nor (_32329_, _32328_, _11842_);
  not (_32330_, _32329_);
  nor (_32331_, _32330_, _32325_);
  nor (_32332_, _32331_, _32324_);
  not (_32333_, _32332_);
  nor (_32334_, _32333_, _32323_);
  nor (_32335_, _32334_, _32173_);
  and (_32336_, _32335_, _32171_);
  nor (_32337_, _04163_, _32171_);
  or (_32339_, _32337_, _32336_);
  and (_32340_, _32339_, _11338_);
  not (_32341_, _32169_);
  and (_32342_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [0]);
  and (_32343_, _32200_, _07871_);
  or (_32344_, _32343_, _32342_);
  and (_32345_, _32344_, _11337_);
  nor (_32346_, _32345_, _32341_);
  not (_32347_, _32346_);
  nor (_32348_, _32347_, _32340_);
  nor (_32350_, _32348_, _32170_);
  and (_32351_, _32350_, _32168_);
  nor (_32352_, _04163_, _32168_);
  or (_32353_, _32352_, _32351_);
  and (_32354_, _32353_, _11881_);
  nor (_32355_, _07955_, _02905_);
  and (_32356_, _07955_, _02905_);
  nor (_32357_, _32356_, _32355_);
  nor (_32358_, _32357_, _11881_);
  and (_32359_, _11330_, _08588_);
  not (_32361_, _32359_);
  nor (_32362_, _32361_, _32358_);
  not (_32363_, _32362_);
  nor (_32364_, _32363_, _32354_);
  nor (_32365_, _32359_, _02905_);
  or (_32366_, _32365_, _03798_);
  nor (_32367_, _32366_, _32364_);
  and (_32368_, _06546_, _03798_);
  or (_32369_, _32368_, _32367_);
  and (_32370_, _32369_, _06399_);
  nor (_32372_, _04163_, _06399_);
  or (_32373_, _32372_, _32370_);
  and (_32374_, _32373_, _11903_);
  and (_32375_, _32212_, _09854_);
  nor (_32376_, _09854_, _02905_);
  or (_32377_, _32376_, _11903_);
  or (_32378_, _32377_, _32375_);
  and (_32379_, _32378_, _32166_);
  not (_32380_, _32379_);
  nor (_32381_, _32380_, _32374_);
  nor (_32383_, _32381_, _32167_);
  and (_32384_, _32383_, _03516_);
  and (_32385_, _06546_, _03515_);
  or (_32386_, _32385_, _32384_);
  and (_32387_, _32386_, _32165_);
  nor (_32388_, _04163_, _32165_);
  nor (_32389_, _32388_, _32387_);
  nor (_32390_, _32389_, _03628_);
  not (_32391_, _32162_);
  and (_32392_, _32160_, _03628_);
  nor (_32394_, _32392_, _32391_);
  not (_32395_, _32394_);
  nor (_32396_, _32395_, _32390_);
  nor (_32397_, _32396_, _32164_);
  nor (_32398_, _32397_, _05103_);
  and (_32399_, _05103_, _04163_);
  nor (_32400_, _32399_, _03453_);
  not (_32401_, _32400_);
  nor (_32402_, _32401_, _32398_);
  nor (_32403_, _32402_, _32161_);
  and (_32405_, _11957_, _11964_);
  not (_32406_, _32405_);
  nor (_32407_, _32406_, _32403_);
  nor (_32408_, _32405_, \oc8051_golden_model_1.PC [0]);
  nor (_32409_, _32408_, _32154_);
  not (_32410_, _32409_);
  nor (_32411_, _32410_, _32407_);
  or (_32412_, _32411_, _11975_);
  nor (_32413_, _32412_, _32155_);
  or (_32414_, _32413_, _32151_);
  or (_32416_, _32414_, _43004_);
  or (_32417_, _43000_, \oc8051_golden_model_1.PC [0]);
  and (_32418_, _32417_, _41806_);
  and (_43667_, _32418_, _32416_);
  and (_32419_, _11975_, _11442_);
  and (_32420_, _03447_, _02878_);
  and (_32421_, _09854_, _11442_);
  nor (_32422_, _11446_, _11444_);
  nor (_32423_, _32422_, _11447_);
  nor (_32424_, _32423_, _09854_);
  nor (_32426_, _32424_, _32421_);
  and (_32427_, _32426_, _03453_);
  nor (_32428_, _11940_, _11442_);
  nor (_32429_, _05848_, _11442_);
  nor (_32430_, _11328_, _11442_);
  nor (_32431_, _11330_, _11442_);
  and (_32432_, _15120_, _03275_);
  nor (_32433_, _11851_, _11442_);
  nor (_32434_, _11345_, _11442_);
  not (_32435_, _04066_);
  nand (_32437_, _08070_, _32435_);
  and (_32438_, _32437_, _03223_);
  and (_32439_, _08055_, _03275_);
  and (_32440_, _10025_, _03275_);
  nor (_32441_, _03617_, _03606_);
  nand (_32442_, _09969_, _03275_);
  not (_32443_, _32423_);
  or (_32444_, _32443_, _09969_);
  and (_32445_, _32444_, _32442_);
  and (_32446_, _32445_, _09917_);
  nor (_32448_, _11666_, _11442_);
  or (_32449_, _32216_, _11442_);
  or (_32450_, _32443_, _11369_);
  and (_32451_, _32450_, _03610_);
  and (_32452_, _32451_, _32449_);
  or (_32453_, _11624_, \oc8051_golden_model_1.PC [1]);
  nor (_32454_, _11573_, _11571_);
  nor (_32455_, _32454_, _11574_);
  nand (_32456_, _32455_, _11624_);
  and (_32457_, _32456_, _06073_);
  and (_32459_, _32457_, _32453_);
  nor (_32460_, _11630_, _11442_);
  or (_32461_, _04303_, _04763_);
  and (_32462_, _04064_, _03275_);
  and (_32463_, _04729_, \oc8051_golden_model_1.PC [0]);
  nor (_32464_, _32463_, _04409_);
  nand (_32465_, _32464_, \oc8051_golden_model_1.PC [1]);
  or (_32466_, _32464_, \oc8051_golden_model_1.PC [1]);
  nand (_32467_, _32466_, _32465_);
  nor (_32468_, _32467_, _04064_);
  or (_32470_, _32468_, _32462_);
  or (_32471_, _32470_, _03980_);
  and (_32472_, _32471_, _11630_);
  and (_32473_, _32472_, _32461_);
  or (_32474_, _32473_, _32460_);
  and (_32475_, _32474_, _06072_);
  or (_32476_, _32475_, _04422_);
  or (_32477_, _32476_, _32459_);
  nand (_32478_, _04422_, _11442_);
  and (_32479_, _32478_, _04081_);
  and (_32481_, _32479_, _32477_);
  or (_32482_, _32481_, _32452_);
  and (_32483_, _32482_, _11362_);
  nor (_32484_, _11362_, _11442_);
  or (_32485_, _32484_, _03715_);
  or (_32486_, _32485_, _32483_);
  nand (_32487_, _03715_, _02878_);
  and (_32488_, _32487_, _03230_);
  and (_32489_, _32488_, _32486_);
  and (_32490_, _04303_, _04768_);
  or (_32492_, _32490_, _03723_);
  or (_32493_, _32492_, _32489_);
  nand (_32494_, _03723_, _02878_);
  and (_32495_, _32494_, _11659_);
  and (_32496_, _32495_, _32493_);
  nor (_32497_, _11659_, _11442_);
  or (_32498_, _32497_, _03729_);
  or (_32499_, _32498_, _32496_);
  nand (_32500_, _03729_, _02878_);
  and (_32501_, _32500_, _11666_);
  and (_32503_, _32501_, _32499_);
  or (_32504_, _32503_, _32448_);
  and (_32505_, _32504_, _03736_);
  and (_32506_, _03714_, \oc8051_golden_model_1.PC [1]);
  or (_32507_, _32506_, _11670_);
  or (_32508_, _32507_, _32505_);
  or (_32509_, _04303_, _03233_);
  and (_32510_, _32509_, _32508_);
  or (_32511_, _32510_, _03508_);
  nand (_32512_, _03508_, _02878_);
  and (_32514_, _32512_, _09921_);
  and (_32515_, _32514_, _32511_);
  or (_32516_, _32515_, _32446_);
  and (_32517_, _32516_, _32441_);
  or (_32518_, _10018_, _11442_);
  not (_32519_, _32441_);
  or (_32520_, _32443_, _11685_);
  and (_32521_, _32520_, _32519_);
  and (_32522_, _32521_, _32518_);
  or (_32523_, _32522_, _03615_);
  or (_32525_, _32523_, _32517_);
  or (_32526_, _32443_, _09876_);
  nand (_32527_, _09876_, _03275_);
  and (_32528_, _32527_, _32526_);
  or (_32529_, _32528_, _04107_);
  and (_32530_, _32529_, _32525_);
  or (_32531_, _32530_, _03604_);
  and (_32532_, _10061_, _11442_);
  nor (_32533_, _32423_, _10061_);
  or (_32534_, _32533_, _09856_);
  or (_32536_, _32534_, _32532_);
  and (_32537_, _32536_, _11358_);
  and (_32538_, _32537_, _32531_);
  or (_32539_, _32538_, _32440_);
  and (_32540_, _32539_, _06840_);
  and (_32541_, _03719_, \oc8051_golden_model_1.PC [1]);
  or (_32542_, _32541_, _04766_);
  or (_32543_, _32542_, _32540_);
  or (_32544_, _04303_, _03227_);
  and (_32545_, _23519_, _11706_);
  and (_32547_, _32545_, _23262_);
  and (_32548_, _32547_, _32544_);
  and (_32549_, _32548_, _32543_);
  nor (_32550_, _32547_, _02878_);
  or (_32551_, _32550_, _32549_);
  and (_32552_, _32551_, _11355_);
  nor (_32553_, _11355_, _11442_);
  or (_32554_, _32553_, _03753_);
  or (_32555_, _32554_, _32552_);
  nand (_32556_, _03753_, _02878_);
  and (_32558_, _32556_, _03238_);
  and (_32559_, _32558_, _32555_);
  and (_32560_, _04303_, _11727_);
  or (_32561_, _32560_, _03752_);
  or (_32562_, _32561_, _32559_);
  and (_32563_, _03752_, _02878_);
  nor (_32564_, _32563_, _08055_);
  and (_32565_, _32564_, _32562_);
  nor (_32566_, _32565_, _32439_);
  nor (_32567_, _32566_, _32438_);
  and (_32569_, _32438_, _03275_);
  nor (_32570_, _04727_, _03247_);
  or (_32571_, _32570_, _32569_);
  or (_32572_, _32571_, _32567_);
  nand (_32573_, _32570_, _11442_);
  and (_32574_, _32573_, _08186_);
  and (_32575_, _32574_, _32572_);
  nor (_32576_, _08186_, _02878_);
  or (_32577_, _32576_, _07912_);
  or (_32578_, _32577_, _32575_);
  or (_32580_, _03275_, _03248_);
  and (_32581_, _32580_, _03710_);
  and (_32582_, _32581_, _32578_);
  and (_32583_, _03505_, \oc8051_golden_model_1.PC [1]);
  or (_32584_, _32583_, _32582_);
  and (_32585_, _32584_, _05897_);
  and (_32586_, _04303_, _03224_);
  or (_32587_, _32586_, _03625_);
  or (_32588_, _32587_, _32585_);
  nand (_32589_, _03625_, _03275_);
  and (_32591_, _32589_, _11749_);
  and (_32592_, _32591_, _32588_);
  nor (_32593_, _11749_, _02878_);
  or (_32594_, _32593_, _03222_);
  or (_32595_, _32594_, _32592_);
  nand (_32596_, _03275_, _03222_);
  and (_32597_, _32596_, _11756_);
  and (_32598_, _32597_, _32595_);
  nor (_32599_, _11756_, _11442_);
  or (_32600_, _32599_, _03585_);
  or (_32602_, _32600_, _32598_);
  nand (_32603_, _03585_, _02878_);
  and (_32604_, _32603_, _03170_);
  and (_32605_, _32604_, _32602_);
  and (_32606_, _04303_, _03169_);
  or (_32607_, _32606_, _11764_);
  or (_32608_, _32607_, _32605_);
  nand (_32609_, _32455_, _11764_);
  and (_32610_, _32609_, _05894_);
  and (_32611_, _32610_, _32608_);
  nor (_32613_, _03601_, \oc8051_golden_model_1.PC [1]);
  nor (_32614_, _32613_, _05895_);
  or (_32615_, _32614_, _32611_);
  nand (_32616_, _03601_, _03275_);
  and (_32617_, _32616_, _08364_);
  and (_32618_, _32617_, _32615_);
  and (_32619_, _08363_, \oc8051_golden_model_1.PC [1]);
  or (_32620_, _32619_, _32618_);
  nand (_32621_, _32620_, _11348_);
  nor (_32622_, _11348_, _03345_);
  nor (_32623_, _32622_, _03584_);
  nand (_32624_, _32623_, _32621_);
  and (_32625_, _03584_, _02878_);
  nor (_32626_, _32625_, _03178_);
  nand (_32627_, _32626_, _32624_);
  and (_32628_, _04303_, _03178_);
  nor (_32629_, _32628_, _11819_);
  nand (_32630_, _32629_, _32627_);
  nor (_32631_, _32455_, _08786_);
  and (_32632_, _08786_, \oc8051_golden_model_1.PC [1]);
  nor (_32635_, _32632_, _11820_);
  not (_32636_, _32635_);
  nor (_32637_, _32636_, _32631_);
  nor (_32638_, _32637_, _11824_);
  and (_32639_, _32638_, _32630_);
  or (_32640_, _32639_, _32434_);
  nand (_32641_, _32640_, _11341_);
  nor (_32642_, _11341_, _02878_);
  nor (_32643_, _32642_, _03600_);
  nand (_32644_, _32643_, _32641_);
  and (_32646_, _03600_, _03275_);
  nor (_32647_, _32646_, _03780_);
  and (_32648_, _32647_, _32644_);
  and (_32649_, _03780_, \oc8051_golden_model_1.PC [1]);
  or (_32650_, _32649_, _32648_);
  nand (_32651_, _32650_, _32175_);
  and (_32652_, _04303_, _03182_);
  nor (_32653_, _32652_, _11841_);
  nand (_32654_, _32653_, _32651_);
  nor (_32655_, _32455_, _11826_);
  nor (_32657_, _08786_, _02878_);
  nor (_32658_, _32657_, _11842_);
  not (_32659_, _32658_);
  nor (_32660_, _32659_, _32655_);
  nor (_32661_, _32660_, _11853_);
  and (_32662_, _32661_, _32654_);
  or (_32663_, _32662_, _32433_);
  nand (_32664_, _32663_, _08430_);
  nor (_32665_, _08430_, _02878_);
  nor (_32666_, _32665_, _03622_);
  nand (_32668_, _32666_, _32664_);
  and (_32669_, _03622_, _03275_);
  nor (_32670_, _32669_, _03790_);
  and (_32671_, _32670_, _32668_);
  and (_32672_, _03790_, \oc8051_golden_model_1.PC [1]);
  or (_32673_, _32672_, _32671_);
  nand (_32674_, _32673_, _32171_);
  and (_32675_, _04303_, _03192_);
  nor (_32676_, _32675_, _11337_);
  nand (_32677_, _32676_, _32674_);
  and (_32679_, \oc8051_golden_model_1.PSW [7], _02878_);
  and (_32680_, _32455_, _07871_);
  or (_32681_, _32680_, _32679_);
  and (_32682_, _32681_, _11337_);
  nor (_32683_, _32682_, _15120_);
  and (_32684_, _32683_, _32677_);
  or (_32685_, _32684_, _32432_);
  nand (_32686_, _08450_, _12559_);
  nor (_32687_, _15123_, _15127_);
  and (_32688_, _32687_, _32686_);
  nand (_32690_, _32688_, _32685_);
  and (_32691_, _03605_, _03200_);
  nor (_32692_, _32688_, _11442_);
  nor (_32693_, _32692_, _32691_);
  nand (_32694_, _32693_, _32690_);
  and (_32695_, _32691_, _11442_);
  nor (_32696_, _32695_, _08460_);
  nand (_32697_, _32696_, _32694_);
  nor (_32698_, _08459_, _02878_);
  nor (_32699_, _32698_, _03624_);
  nand (_32701_, _32699_, _32697_);
  and (_32702_, _03624_, _03275_);
  nor (_32703_, _32702_, _03785_);
  and (_32704_, _32703_, _32701_);
  and (_32705_, _03785_, \oc8051_golden_model_1.PC [1]);
  or (_32706_, _32705_, _32704_);
  nand (_32707_, _32706_, _32168_);
  and (_32708_, _04303_, _03201_);
  nor (_32709_, _32708_, _11880_);
  nand (_32710_, _32709_, _32707_);
  nor (_32712_, _32455_, _07871_);
  and (_32713_, _07871_, \oc8051_golden_model_1.PC [1]);
  nor (_32714_, _32713_, _11881_);
  not (_32715_, _32714_);
  nor (_32716_, _32715_, _32712_);
  nor (_32717_, _32716_, _11885_);
  and (_32718_, _32717_, _32710_);
  or (_32719_, _32718_, _32431_);
  nand (_32720_, _32719_, _08507_);
  nor (_32721_, _08507_, _02878_);
  nor (_32723_, _32721_, _08587_);
  nand (_32724_, _32723_, _32720_);
  and (_32725_, _08587_, _11442_);
  nor (_32726_, _32725_, _03798_);
  and (_32727_, _32726_, _32724_);
  nor (_32728_, _06501_, _10652_);
  or (_32729_, _32728_, _32727_);
  nand (_32730_, _32729_, _06399_);
  and (_32731_, _04303_, _03188_);
  nor (_32732_, _32731_, _03621_);
  nand (_32734_, _32732_, _32730_);
  nor (_32735_, _09854_, _03275_);
  and (_32736_, _32443_, _09854_);
  or (_32737_, _32736_, _11903_);
  nor (_32738_, _32737_, _32735_);
  nor (_32739_, _32738_, _11907_);
  and (_32740_, _32739_, _32734_);
  or (_32741_, _32740_, _32430_);
  nand (_32742_, _32741_, _08702_);
  nor (_32743_, _08702_, _02878_);
  nor (_32745_, _32743_, _08732_);
  nand (_32746_, _32745_, _32742_);
  and (_32747_, _08732_, _11442_);
  nor (_32748_, _32747_, _03515_);
  and (_32749_, _32748_, _32746_);
  nor (_32750_, _06501_, _03516_);
  or (_32751_, _32750_, _32749_);
  nand (_32752_, _32751_, _32165_);
  and (_32753_, _04303_, _03203_);
  nor (_32754_, _32753_, _03628_);
  nand (_32756_, _32754_, _32752_);
  and (_32757_, _32426_, _03628_);
  nor (_32758_, _32757_, _12561_);
  and (_32759_, _32758_, _32756_);
  or (_32760_, _32759_, _32429_);
  nand (_32761_, _32760_, _06409_);
  and (_32762_, _04533_, _03275_);
  nor (_32763_, _32762_, _03815_);
  nand (_32764_, _32763_, _32761_);
  not (_32765_, _11940_);
  and (_32767_, _03815_, _02878_);
  nor (_32768_, _32767_, _32765_);
  and (_32769_, _32768_, _32764_);
  or (_32770_, _32769_, _32428_);
  nand (_32771_, _32770_, _04540_);
  and (_32772_, _05103_, _04303_);
  nor (_32773_, _32772_, _03453_);
  and (_32774_, _32773_, _32771_);
  or (_32775_, _32774_, _32427_);
  nand (_32776_, _32775_, _11955_);
  nor (_32778_, _11955_, _03275_);
  nor (_32779_, _32778_, _04552_);
  nand (_32780_, _32779_, _32776_);
  and (_32781_, _04552_, _03275_);
  nor (_32782_, _32781_, _03447_);
  and (_32783_, _32782_, _32780_);
  or (_32784_, _32783_, _32420_);
  nand (_32785_, _32784_, _11964_);
  nor (_32786_, _11964_, _03275_);
  nor (_32787_, _32786_, _32154_);
  nand (_32789_, _32787_, _32785_);
  and (_32790_, _32154_, _04303_);
  nor (_32791_, _32790_, _11975_);
  and (_32792_, _32791_, _32789_);
  or (_32793_, _32792_, _32419_);
  or (_32794_, _32793_, _43004_);
  or (_32795_, _43000_, \oc8051_golden_model_1.PC [1]);
  and (_32796_, _32795_, _41806_);
  and (_43670_, _32796_, _32794_);
  and (_32797_, _03447_, _03210_);
  nor (_32799_, _11328_, _03266_);
  nor (_32800_, _11330_, _03266_);
  nor (_32801_, _11335_, _03266_);
  nor (_32802_, _11851_, _03266_);
  nor (_32803_, _11345_, _03266_);
  and (_32804_, _03505_, _03245_);
  nor (_32805_, _32547_, _03210_);
  not (_32806_, _03266_);
  and (_32807_, _10025_, _32806_);
  and (_32808_, _03980_, _03946_);
  nor (_32810_, _11643_, _03266_);
  and (_32811_, _03979_, _03245_);
  or (_32812_, _04409_, \oc8051_golden_model_1.PC [2]);
  nor (_32813_, _32812_, _04729_);
  or (_32814_, _32813_, _32811_);
  not (_32815_, _11632_);
  and (_32816_, _32190_, _32815_);
  and (_32817_, _32816_, _32814_);
  or (_32818_, _32817_, _32810_);
  or (_32819_, _32818_, _32808_);
  and (_32821_, _32819_, _06072_);
  and (_32822_, _11578_, _11575_);
  nor (_32823_, _32822_, _11579_);
  nand (_32824_, _32823_, _11624_);
  or (_32825_, _11624_, _03245_);
  and (_32826_, _32825_, _06073_);
  and (_32827_, _32826_, _32824_);
  or (_32828_, _32827_, _32821_);
  and (_32829_, _32828_, _05966_);
  and (_32830_, _04422_, _32806_);
  or (_32832_, _32830_, _03610_);
  or (_32833_, _32832_, _32829_);
  and (_32834_, _11451_, _11448_);
  nor (_32835_, _32834_, _11452_);
  not (_32836_, _32835_);
  and (_32837_, _32836_, _11367_);
  and (_32838_, _11440_, _11369_);
  or (_32839_, _32838_, _04081_);
  or (_32840_, _32839_, _32837_);
  and (_32841_, _32840_, _11362_);
  and (_32843_, _32841_, _32833_);
  nor (_32844_, _11362_, _03266_);
  or (_32845_, _32844_, _03715_);
  or (_32846_, _32845_, _32843_);
  nand (_32847_, _03715_, _03210_);
  and (_32848_, _32847_, _03230_);
  and (_32849_, _32848_, _32846_);
  and (_32850_, _03946_, _04768_);
  or (_32851_, _32850_, _03723_);
  or (_32852_, _32851_, _32849_);
  nand (_32854_, _03723_, _03210_);
  and (_32855_, _32854_, _11659_);
  and (_32856_, _32855_, _32852_);
  nor (_32857_, _11659_, _03266_);
  or (_32858_, _32857_, _03729_);
  or (_32859_, _32858_, _32856_);
  nand (_32860_, _03729_, _03210_);
  and (_32861_, _32860_, _11666_);
  and (_32862_, _32861_, _32859_);
  nor (_32863_, _11666_, _03266_);
  or (_32865_, _32863_, _03714_);
  or (_32866_, _32865_, _32862_);
  nand (_32867_, _03714_, _03210_);
  and (_32868_, _32867_, _03233_);
  and (_32869_, _32868_, _32866_);
  and (_32870_, _03946_, _11670_);
  or (_32871_, _32870_, _03508_);
  or (_32872_, _32871_, _32869_);
  nand (_32873_, _03508_, _03210_);
  and (_32874_, _32873_, _09921_);
  and (_32876_, _32874_, _32872_);
  or (_32877_, _32836_, _09969_);
  nand (_32878_, _11439_, _09969_);
  and (_32879_, _32878_, _09917_);
  nand (_32880_, _32879_, _32877_);
  nand (_32881_, _32880_, _23483_);
  or (_32882_, _32881_, _32876_);
  or (_32883_, _32836_, _09876_);
  nand (_32884_, _11439_, _09876_);
  and (_32885_, _32884_, _32883_);
  or (_32887_, _32885_, _04107_);
  or (_32888_, _32836_, _11685_);
  or (_32889_, _11440_, _10018_);
  and (_32890_, _32889_, _32888_);
  or (_32891_, _32890_, _09920_);
  and (_32892_, _32891_, _32887_);
  and (_32893_, _32892_, _32882_);
  or (_32894_, _32893_, _03604_);
  and (_32895_, _11440_, _10061_);
  nor (_32896_, _32835_, _10061_);
  or (_32898_, _32896_, _09856_);
  or (_32899_, _32898_, _32895_);
  and (_32900_, _32899_, _11358_);
  and (_32901_, _32900_, _32894_);
  or (_32902_, _32901_, _32807_);
  and (_32903_, _32902_, _06840_);
  and (_32904_, _03719_, _03245_);
  or (_32905_, _32904_, _04766_);
  or (_32906_, _32905_, _32903_);
  or (_32907_, _03946_, _03227_);
  and (_32909_, _32907_, _32547_);
  and (_32910_, _32909_, _32906_);
  or (_32911_, _32910_, _32805_);
  and (_32912_, _32911_, _11355_);
  nor (_32913_, _11355_, _03266_);
  or (_32914_, _32913_, _03753_);
  or (_32915_, _32914_, _32912_);
  nand (_32916_, _03753_, _03210_);
  and (_32917_, _32916_, _03238_);
  and (_32918_, _32917_, _32915_);
  and (_32920_, _03946_, _11727_);
  or (_32921_, _32920_, _03752_);
  or (_32922_, _32921_, _32918_);
  nand (_32923_, _03752_, _03210_);
  and (_32924_, _32923_, _11350_);
  and (_32925_, _32924_, _32922_);
  nor (_32926_, _11350_, _03266_);
  or (_32927_, _32926_, _32925_);
  and (_32928_, _32927_, _08186_);
  nor (_32929_, _08186_, _03210_);
  or (_32931_, _32929_, _07912_);
  or (_32932_, _32931_, _32928_);
  or (_32933_, _32806_, _03248_);
  and (_32934_, _32933_, _03710_);
  and (_32935_, _32934_, _32932_);
  or (_32936_, _32935_, _32804_);
  and (_32937_, _32936_, _05897_);
  and (_32938_, _03946_, _03224_);
  or (_32939_, _32938_, _03625_);
  or (_32940_, _32939_, _32937_);
  and (_32942_, _11439_, _03625_);
  nor (_32943_, _32942_, _04475_);
  and (_32944_, _32943_, _32940_);
  and (_32945_, _04475_, _03245_);
  or (_32946_, _06835_, _03969_);
  or (_32947_, _32946_, _32945_);
  or (_32948_, _32947_, _32944_);
  nand (_32949_, _32946_, _03210_);
  and (_32950_, _32949_, _11748_);
  and (_32951_, _32950_, _32948_);
  nor (_32953_, _11748_, _03210_);
  or (_32954_, _32953_, _03222_);
  or (_32955_, _32954_, _32951_);
  nand (_32956_, _11439_, _03222_);
  and (_32957_, _32956_, _11756_);
  and (_32958_, _32957_, _32955_);
  nor (_32959_, _11756_, _03266_);
  or (_32960_, _32959_, _03585_);
  or (_32961_, _32960_, _32958_);
  nand (_32962_, _03585_, _03210_);
  and (_32964_, _32962_, _03170_);
  and (_32965_, _32964_, _32961_);
  and (_32966_, _03946_, _03169_);
  or (_32967_, _32966_, _32965_);
  and (_32968_, _32967_, _11765_);
  nor (_32969_, _32823_, _11765_);
  or (_32970_, _32969_, _06168_);
  or (_32971_, _32970_, _32968_);
  or (_32972_, _05894_, _03245_);
  and (_32973_, _32972_, _05886_);
  and (_32974_, _32973_, _32971_);
  and (_32975_, _11440_, _03601_);
  or (_32976_, _32975_, _08363_);
  or (_32977_, _32976_, _32974_);
  and (_32978_, _08363_, _03210_);
  nor (_32979_, _32978_, _11347_);
  and (_32980_, _32979_, _32977_);
  and (_32981_, _11347_, _03262_);
  or (_32982_, _32981_, _03584_);
  or (_32983_, _32982_, _32980_);
  nand (_32986_, _03584_, _03210_);
  and (_32987_, _32986_, _10736_);
  and (_32988_, _32987_, _32983_);
  and (_32989_, _03946_, _03178_);
  or (_32990_, _32989_, _11819_);
  or (_32991_, _32990_, _32988_);
  nor (_32992_, _32823_, _08786_);
  nand (_32993_, _08786_, _03245_);
  nand (_32994_, _32993_, _11819_);
  or (_32995_, _32994_, _32992_);
  and (_32997_, _32995_, _11345_);
  and (_32998_, _32997_, _32991_);
  or (_32999_, _32998_, _32803_);
  and (_33000_, _32999_, _11341_);
  nor (_33001_, _11341_, _03210_);
  or (_33002_, _33001_, _03600_);
  or (_33003_, _33002_, _33000_);
  nand (_33004_, _11439_, _03600_);
  and (_33005_, _33004_, _07778_);
  and (_33006_, _33005_, _33003_);
  and (_33008_, _03780_, _03245_);
  or (_33009_, _33008_, _33006_);
  and (_33010_, _33009_, _32175_);
  and (_33011_, _03946_, _03182_);
  or (_33012_, _33011_, _11841_);
  or (_33013_, _33012_, _33010_);
  or (_33014_, _32823_, _11826_);
  or (_33015_, _08786_, _03210_);
  and (_33016_, _33015_, _11841_);
  and (_33017_, _33016_, _33014_);
  nor (_33019_, _33017_, _11853_);
  and (_33020_, _33019_, _33013_);
  or (_33021_, _33020_, _32802_);
  and (_33022_, _33021_, _08430_);
  nor (_33023_, _08430_, _03210_);
  or (_33024_, _33023_, _03622_);
  or (_33025_, _33024_, _33022_);
  nand (_33026_, _11439_, _03622_);
  and (_33027_, _33026_, _06828_);
  and (_33028_, _33027_, _33025_);
  and (_33029_, _03790_, _03245_);
  or (_33030_, _33029_, _33028_);
  and (_33031_, _33030_, _32171_);
  and (_33032_, _03946_, _03192_);
  or (_33033_, _33032_, _11337_);
  or (_33034_, _33033_, _33031_);
  nor (_33035_, _32823_, \oc8051_golden_model_1.PSW [7]);
  or (_33036_, _03210_, _07871_);
  nand (_33037_, _33036_, _11337_);
  or (_33038_, _33037_, _33035_);
  and (_33040_, _33038_, _11335_);
  and (_33041_, _33040_, _33034_);
  or (_33042_, _33041_, _32801_);
  and (_33043_, _33042_, _08459_);
  nor (_33044_, _08459_, _03210_);
  or (_33045_, _33044_, _03624_);
  or (_33046_, _33045_, _33043_);
  nand (_33047_, _11439_, _03624_);
  and (_33048_, _33047_, _07793_);
  and (_33049_, _33048_, _33046_);
  and (_33051_, _03785_, _03245_);
  or (_33052_, _33051_, _33049_);
  and (_33053_, _33052_, _32168_);
  and (_33054_, _03946_, _03201_);
  or (_33055_, _33054_, _11880_);
  or (_33056_, _33055_, _33053_);
  nor (_33057_, _32823_, _07871_);
  or (_33058_, _03210_, \oc8051_golden_model_1.PSW [7]);
  nand (_33059_, _33058_, _11880_);
  or (_33060_, _33059_, _33057_);
  and (_33062_, _33060_, _11330_);
  and (_33063_, _33062_, _33056_);
  or (_33064_, _33063_, _32800_);
  and (_33065_, _33064_, _08507_);
  nor (_33066_, _08507_, _03210_);
  or (_33067_, _33066_, _08587_);
  or (_33068_, _33067_, _33065_);
  nand (_33069_, _08587_, _03266_);
  and (_33070_, _33069_, _10652_);
  and (_33071_, _33070_, _33068_);
  nor (_33073_, _06637_, _10652_);
  or (_33074_, _33073_, _33071_);
  and (_33075_, _33074_, _06399_);
  and (_33076_, _03946_, _03188_);
  or (_33077_, _33076_, _03621_);
  or (_33078_, _33077_, _33075_);
  and (_33079_, _32836_, _09854_);
  nor (_33080_, _11439_, _09854_);
  or (_33081_, _33080_, _11903_);
  or (_33082_, _33081_, _33079_);
  and (_33084_, _33082_, _11328_);
  and (_33085_, _33084_, _33078_);
  or (_33086_, _33085_, _32799_);
  and (_33087_, _33086_, _08702_);
  nor (_33088_, _08702_, _03210_);
  or (_33089_, _33088_, _08732_);
  or (_33090_, _33089_, _33087_);
  nand (_33091_, _08732_, _03266_);
  and (_33092_, _33091_, _03516_);
  and (_33093_, _33092_, _33090_);
  nor (_33095_, _06637_, _03516_);
  or (_33096_, _33095_, _33093_);
  and (_33097_, _33096_, _32165_);
  and (_33098_, _03946_, _03203_);
  or (_33099_, _33098_, _03628_);
  or (_33100_, _33099_, _33097_);
  nor (_33101_, _32835_, _09854_);
  and (_33102_, _11440_, _09854_);
  nor (_33103_, _33102_, _33101_);
  nand (_33104_, _33103_, _03628_);
  and (_33106_, _33104_, _11933_);
  and (_33107_, _33106_, _33100_);
  nor (_33108_, _11933_, _03266_);
  or (_33109_, _33108_, _03815_);
  or (_33110_, _33109_, _33107_);
  and (_33111_, _03815_, _03210_);
  nor (_33112_, _33111_, _32765_);
  and (_33113_, _33112_, _33110_);
  nor (_33114_, _11940_, _03266_);
  or (_33115_, _33114_, _33113_);
  and (_33117_, _33115_, _04540_);
  and (_33118_, _05103_, _03946_);
  nor (_33119_, _33118_, _03453_);
  not (_33120_, _33119_);
  or (_33121_, _33120_, _33117_);
  and (_33122_, _33103_, _03453_);
  nor (_33123_, _33122_, _11958_);
  nand (_33124_, _33123_, _33121_);
  nor (_33125_, _11957_, _03266_);
  nor (_33126_, _33125_, _03447_);
  and (_33128_, _33126_, _33124_);
  or (_33129_, _33128_, _32797_);
  nand (_33130_, _33129_, _11964_);
  nor (_33131_, _11964_, _32806_);
  nor (_33132_, _33131_, _32154_);
  nand (_33133_, _33132_, _33130_);
  and (_33134_, _32154_, _03946_);
  nor (_33135_, _33134_, _11975_);
  and (_33136_, _33135_, _33133_);
  and (_33137_, _11975_, _03266_);
  or (_33139_, _33137_, _33136_);
  or (_33140_, _33139_, _43004_);
  or (_33141_, _43000_, \oc8051_golden_model_1.PC [2]);
  and (_33142_, _33141_, _41806_);
  and (_43671_, _33142_, _33140_);
  and (_33143_, _03447_, _03297_);
  and (_33144_, _03815_, _03297_);
  nor (_33145_, _11328_, _03650_);
  nor (_33146_, _11330_, _03650_);
  nor (_33147_, _11335_, _03650_);
  nor (_33149_, _11851_, _03650_);
  nor (_33150_, _11345_, _03650_);
  and (_33151_, _08363_, _03648_);
  and (_33152_, _03505_, _03648_);
  nor (_33153_, _11350_, _03650_);
  nor (_33154_, _32547_, _03297_);
  and (_33155_, _10025_, _03311_);
  and (_33156_, _11504_, _03648_);
  or (_33157_, _11568_, _11567_);
  and (_33158_, _33157_, _11580_);
  nor (_33160_, _33157_, _11580_);
  nor (_33161_, _33160_, _33158_);
  not (_33162_, _33161_);
  and (_33163_, _33162_, _11624_);
  or (_33164_, _33163_, _06072_);
  or (_33165_, _33164_, _33156_);
  and (_33166_, _03980_, _03708_);
  nor (_33167_, _11642_, _03650_);
  and (_33168_, _03979_, _03648_);
  not (_33169_, _04729_);
  nor (_33171_, _04409_, \oc8051_golden_model_1.PC [3]);
  and (_33172_, _33171_, _33169_);
  nor (_33173_, _33172_, _33168_);
  nor (_33174_, _33173_, _11632_);
  nor (_33175_, _33174_, _33167_);
  nor (_33176_, _33175_, _32191_);
  nor (_33177_, _11630_, _03650_);
  or (_33178_, _33177_, _06073_);
  or (_33179_, _33178_, _33176_);
  or (_33180_, _33179_, _33166_);
  and (_33182_, _33180_, _33165_);
  nand (_33183_, _33182_, _05966_);
  and (_33184_, _04422_, _03311_);
  nor (_33185_, _33184_, _03610_);
  and (_33186_, _33185_, _33183_);
  or (_33187_, _11435_, _11367_);
  or (_33188_, _11437_, _11436_);
  and (_33189_, _33188_, _11453_);
  nor (_33190_, _33188_, _11453_);
  nor (_33191_, _33190_, _33189_);
  not (_33193_, _33191_);
  or (_33194_, _33193_, _11369_);
  nand (_33195_, _33194_, _33187_);
  and (_33196_, _33195_, _03610_);
  nor (_33197_, _33196_, _33186_);
  nand (_33198_, _33197_, _11362_);
  nor (_33199_, _11362_, _03650_);
  nor (_33200_, _33199_, _03715_);
  nand (_33201_, _33200_, _33198_);
  and (_33202_, _03715_, _03297_);
  nor (_33204_, _33202_, _04768_);
  nand (_33205_, _33204_, _33201_);
  and (_33206_, _03708_, _04768_);
  nor (_33207_, _33206_, _03723_);
  nand (_33208_, _33207_, _33205_);
  and (_33209_, _03723_, _03297_);
  nor (_33210_, _33209_, _11660_);
  nand (_33211_, _33210_, _33208_);
  nor (_33212_, _11659_, _03650_);
  nor (_33213_, _33212_, _03729_);
  nand (_33215_, _33213_, _33211_);
  and (_33216_, _03729_, _03297_);
  nor (_33217_, _33216_, _11668_);
  nand (_33218_, _33217_, _33215_);
  nor (_33219_, _11666_, _03650_);
  nor (_33220_, _33219_, _03714_);
  nand (_33221_, _33220_, _33218_);
  and (_33222_, _03714_, _03297_);
  nor (_33223_, _33222_, _11670_);
  nand (_33224_, _33223_, _33221_);
  and (_33226_, _03708_, _11670_);
  nor (_33227_, _33226_, _03508_);
  nand (_33228_, _33227_, _33224_);
  and (_33229_, _03508_, _03297_);
  nor (_33230_, _33229_, _09917_);
  nand (_33231_, _33230_, _33228_);
  not (_33232_, _23483_);
  and (_33233_, _11434_, _09969_);
  nor (_33234_, _33193_, _09969_);
  or (_33235_, _33234_, _09921_);
  nor (_33237_, _33235_, _33233_);
  nor (_33238_, _33237_, _33232_);
  nand (_33239_, _33238_, _33231_);
  and (_33240_, _11434_, _09876_);
  nor (_33241_, _33193_, _09876_);
  nor (_33242_, _33241_, _33240_);
  nor (_33243_, _33242_, _04107_);
  or (_33244_, _11435_, _10018_);
  or (_33245_, _33193_, _11685_);
  nand (_33246_, _33245_, _33244_);
  and (_33248_, _33246_, _09919_);
  nor (_33249_, _33248_, _33243_);
  nand (_33250_, _33249_, _33239_);
  nand (_33251_, _33250_, _09856_);
  nor (_33252_, _33191_, _10061_);
  and (_33253_, _11435_, _10061_);
  or (_33254_, _33253_, _09856_);
  nor (_33255_, _33254_, _33252_);
  nor (_33256_, _33255_, _10025_);
  and (_33257_, _33256_, _33251_);
  or (_33259_, _33257_, _33155_);
  nand (_33260_, _33259_, _06840_);
  and (_33261_, _03719_, _03648_);
  nor (_33262_, _33261_, _04766_);
  nand (_33263_, _33262_, _33260_);
  not (_33264_, _32547_);
  nor (_33265_, _03708_, _03227_);
  nor (_33266_, _33265_, _33264_);
  and (_33267_, _33266_, _33263_);
  or (_33268_, _33267_, _33154_);
  nand (_33270_, _33268_, _11355_);
  nor (_33271_, _11355_, _03650_);
  nor (_33272_, _33271_, _03753_);
  nand (_33273_, _33272_, _33270_);
  and (_33274_, _03753_, _03297_);
  nor (_33275_, _33274_, _11727_);
  nand (_33276_, _33275_, _33273_);
  and (_33277_, _03708_, _11727_);
  nor (_33278_, _33277_, _03752_);
  nand (_33279_, _33278_, _33276_);
  and (_33281_, _03752_, _03297_);
  not (_33282_, _33281_);
  and (_33283_, _33282_, _11350_);
  and (_33284_, _33283_, _33279_);
  or (_33285_, _33284_, _33153_);
  nand (_33286_, _33285_, _08186_);
  nor (_33287_, _08186_, _03297_);
  nor (_33288_, _33287_, _07912_);
  nand (_33289_, _33288_, _33286_);
  nor (_33290_, _03248_, _03311_);
  nor (_33292_, _33290_, _03505_);
  and (_33293_, _33292_, _33289_);
  or (_33294_, _33293_, _33152_);
  nand (_33295_, _33294_, _05897_);
  and (_33296_, _03708_, _03224_);
  nor (_33297_, _33296_, _03625_);
  nand (_33298_, _33297_, _33295_);
  not (_33299_, _11749_);
  and (_33300_, _11434_, _03625_);
  nor (_33301_, _33300_, _33299_);
  nand (_33303_, _33301_, _33298_);
  nor (_33304_, _11749_, _03297_);
  nor (_33305_, _33304_, _03222_);
  nand (_33306_, _33305_, _33303_);
  and (_33307_, _11434_, _03222_);
  nor (_33308_, _33307_, _11758_);
  nand (_33309_, _33308_, _33306_);
  nor (_33310_, _11756_, _03650_);
  nor (_33311_, _33310_, _03585_);
  and (_33312_, _33311_, _33309_);
  and (_33314_, _03585_, _03297_);
  or (_33315_, _33314_, _03169_);
  or (_33316_, _33315_, _33312_);
  and (_33317_, _03708_, _03169_);
  nor (_33318_, _33317_, _11764_);
  nand (_33319_, _33318_, _33316_);
  and (_33320_, _33161_, _11764_);
  nor (_33321_, _33320_, _06168_);
  nand (_33322_, _33321_, _33319_);
  nor (_33323_, _05894_, _03297_);
  nor (_33325_, _33323_, _03601_);
  nand (_33326_, _33325_, _33322_);
  and (_33327_, _11434_, _03601_);
  nor (_33328_, _33327_, _08363_);
  and (_33329_, _33328_, _33326_);
  or (_33330_, _33329_, _33151_);
  nand (_33331_, _33330_, _11348_);
  nor (_33332_, _11348_, _03307_);
  nor (_33333_, _33332_, _03584_);
  nand (_33334_, _33333_, _33331_);
  and (_33336_, _03584_, _03297_);
  nor (_33337_, _33336_, _03178_);
  nand (_33338_, _33337_, _33334_);
  and (_33339_, _03708_, _03178_);
  nor (_33340_, _33339_, _11819_);
  nand (_33341_, _33340_, _33338_);
  and (_33342_, _08786_, _03297_);
  and (_33343_, _33161_, _11826_);
  or (_33344_, _33343_, _33342_);
  and (_33345_, _33344_, _11819_);
  nor (_33346_, _33345_, _11824_);
  and (_33347_, _33346_, _33341_);
  or (_33348_, _33347_, _33150_);
  nand (_33349_, _33348_, _11341_);
  nor (_33350_, _11341_, _03297_);
  nor (_33351_, _33350_, _03600_);
  and (_33352_, _33351_, _33349_);
  and (_33353_, _11434_, _03600_);
  or (_33354_, _33353_, _03780_);
  nor (_33355_, _33354_, _33352_);
  and (_33358_, _03780_, _03648_);
  or (_33359_, _33358_, _33355_);
  nand (_33360_, _33359_, _32175_);
  and (_33361_, _03708_, _03182_);
  nor (_33362_, _33361_, _11841_);
  nand (_33363_, _33362_, _33360_);
  or (_33364_, _33161_, _11826_);
  or (_33365_, _08786_, _03297_);
  and (_33366_, _33365_, _11841_);
  and (_33367_, _33366_, _33364_);
  nor (_33369_, _33367_, _11853_);
  and (_33370_, _33369_, _33363_);
  or (_33371_, _33370_, _33149_);
  nand (_33372_, _33371_, _08430_);
  nor (_33373_, _08430_, _03297_);
  nor (_33374_, _33373_, _03622_);
  and (_33375_, _33374_, _33372_);
  and (_33376_, _11434_, _03622_);
  or (_33377_, _33376_, _03790_);
  nor (_33378_, _33377_, _33375_);
  and (_33380_, _03790_, _03648_);
  or (_33381_, _33380_, _33378_);
  nand (_33382_, _33381_, _32171_);
  and (_33383_, _03708_, _03192_);
  nor (_33384_, _33383_, _11337_);
  nand (_33385_, _33384_, _33382_);
  and (_33386_, _03297_, \oc8051_golden_model_1.PSW [7]);
  and (_33387_, _33161_, _07871_);
  or (_33388_, _33387_, _33386_);
  and (_33389_, _33388_, _11337_);
  nor (_33391_, _33389_, _11864_);
  and (_33392_, _33391_, _33385_);
  or (_33393_, _33392_, _33147_);
  nand (_33394_, _33393_, _08459_);
  nor (_33395_, _08459_, _03297_);
  nor (_33396_, _33395_, _03624_);
  and (_33397_, _33396_, _33394_);
  and (_33398_, _11434_, _03624_);
  or (_33399_, _33398_, _03785_);
  nor (_33400_, _33399_, _33397_);
  and (_33402_, _03785_, _03648_);
  or (_33403_, _33402_, _33400_);
  nand (_33404_, _33403_, _32168_);
  and (_33405_, _03708_, _03201_);
  nor (_33406_, _33405_, _11880_);
  nand (_33407_, _33406_, _33404_);
  nor (_33408_, _33161_, _07871_);
  nor (_33409_, _03297_, \oc8051_golden_model_1.PSW [7]);
  nor (_33410_, _33409_, _11881_);
  not (_33411_, _33410_);
  nor (_33413_, _33411_, _33408_);
  nor (_33414_, _33413_, _11885_);
  and (_33415_, _33414_, _33407_);
  or (_33416_, _33415_, _33146_);
  nand (_33417_, _33416_, _08507_);
  nor (_33418_, _08507_, _03297_);
  nor (_33419_, _33418_, _08587_);
  and (_33420_, _33419_, _33417_);
  and (_33421_, _08587_, _03650_);
  or (_33422_, _33421_, _03798_);
  nor (_33424_, _33422_, _33420_);
  and (_33425_, _08636_, _03798_);
  or (_33426_, _33425_, _33424_);
  nand (_33427_, _33426_, _06399_);
  and (_33428_, _03708_, _03188_);
  nor (_33429_, _33428_, _03621_);
  nand (_33430_, _33429_, _33427_);
  and (_33431_, _33193_, _09854_);
  nor (_33432_, _11434_, _09854_);
  or (_33433_, _33432_, _11903_);
  or (_33435_, _33433_, _33431_);
  and (_33436_, _33435_, _11328_);
  and (_33437_, _33436_, _33430_);
  or (_33438_, _33437_, _33145_);
  nand (_33439_, _33438_, _08702_);
  nor (_33440_, _08702_, _03297_);
  nor (_33441_, _33440_, _08732_);
  and (_33442_, _33441_, _33439_);
  and (_33443_, _08732_, _03650_);
  or (_33444_, _33443_, _03515_);
  nor (_33446_, _33444_, _33442_);
  and (_33447_, _08636_, _03515_);
  or (_33448_, _33447_, _33446_);
  nand (_33449_, _33448_, _32165_);
  and (_33450_, _03708_, _03203_);
  nor (_33451_, _33450_, _03628_);
  nand (_33452_, _33451_, _33449_);
  nor (_33453_, _33191_, _09854_);
  and (_33454_, _11435_, _09854_);
  nor (_33455_, _33454_, _33453_);
  and (_33457_, _33455_, _03628_);
  nor (_33458_, _33457_, _11934_);
  nand (_33459_, _33458_, _33452_);
  nor (_33460_, _11933_, _03650_);
  nor (_33461_, _33460_, _03815_);
  and (_33462_, _33461_, _33459_);
  or (_33463_, _33462_, _33144_);
  nand (_33464_, _33463_, _11940_);
  nor (_33465_, _11940_, _03311_);
  nor (_33466_, _33465_, _05103_);
  nand (_33468_, _33466_, _33464_);
  and (_33469_, _05103_, _03708_);
  nor (_33470_, _33469_, _03453_);
  nand (_33471_, _33470_, _33468_);
  and (_33472_, _33455_, _03453_);
  nor (_33473_, _33472_, _11958_);
  nand (_33474_, _33473_, _33471_);
  nor (_33475_, _11957_, _03650_);
  nor (_33476_, _33475_, _03447_);
  and (_33477_, _33476_, _33474_);
  or (_33479_, _33477_, _33143_);
  nand (_33480_, _33479_, _11964_);
  nor (_33481_, _11964_, _03311_);
  nor (_33482_, _33481_, _32154_);
  nand (_33483_, _33482_, _33480_);
  and (_33484_, _32154_, _03708_);
  nor (_33485_, _33484_, _11975_);
  and (_33486_, _33485_, _33483_);
  and (_33487_, _11975_, _03650_);
  or (_33488_, _33487_, _33486_);
  or (_33490_, _33488_, _43004_);
  or (_33491_, _43000_, \oc8051_golden_model_1.PC [3]);
  and (_33492_, _33491_, _41806_);
  and (_43672_, _33492_, _33490_);
  and (_33493_, _06236_, _05103_);
  and (_33494_, _11565_, _03780_);
  and (_33495_, _11564_, _08786_);
  and (_33496_, _11585_, _11582_);
  nor (_33497_, _33496_, _11586_);
  and (_33498_, _33497_, _11826_);
  or (_33500_, _33498_, _33495_);
  and (_33501_, _33500_, _11819_);
  nor (_33502_, _32547_, _11564_);
  not (_33503_, \oc8051_golden_model_1.PC [4]);
  nor (_33504_, _02892_, _33503_);
  and (_33505_, _02892_, _33503_);
  nor (_33506_, _33505_, _33504_);
  not (_33507_, _33506_);
  and (_33508_, _33507_, _10025_);
  and (_33509_, _11565_, _03714_);
  nor (_33511_, _33506_, _11659_);
  and (_33512_, _11458_, _11455_);
  nor (_33513_, _33512_, _11459_);
  or (_33514_, _33513_, _11369_);
  and (_33515_, _33514_, _03610_);
  or (_33516_, _11430_, _11367_);
  and (_33517_, _33516_, _33515_);
  nand (_33518_, _33497_, _11624_);
  or (_33519_, _11624_, _11565_);
  and (_33520_, _33519_, _06073_);
  nand (_33522_, _33520_, _33518_);
  not (_33523_, _11647_);
  and (_33524_, _06236_, _03980_);
  nor (_33525_, _33506_, _11642_);
  and (_33526_, _11565_, _03979_);
  nor (_33527_, _04409_, \oc8051_golden_model_1.PC [4]);
  and (_33528_, _33527_, _33169_);
  nor (_33529_, _33528_, _33526_);
  nor (_33530_, _33529_, _11632_);
  nor (_33531_, _33530_, _33525_);
  nor (_33533_, _33531_, _03980_);
  nor (_33534_, _33533_, _11631_);
  not (_33535_, _33534_);
  nor (_33536_, _33535_, _33524_);
  nor (_33537_, _33507_, _11630_);
  nor (_33538_, _33537_, _06073_);
  not (_33539_, _33538_);
  nor (_33540_, _33539_, _33536_);
  nor (_33541_, _33540_, _33523_);
  and (_33542_, _33541_, _33522_);
  or (_33544_, _33542_, _33517_);
  and (_33545_, _33544_, _11362_);
  nor (_33546_, _33507_, _11653_);
  or (_33547_, _33546_, _03715_);
  or (_33548_, _33547_, _33545_);
  and (_33549_, _11565_, _03715_);
  nor (_33550_, _33549_, _04768_);
  and (_33551_, _33550_, _33548_);
  nor (_33552_, _06236_, _03230_);
  or (_33553_, _33552_, _03723_);
  nor (_33555_, _33553_, _33551_);
  and (_33556_, _11565_, _03723_);
  or (_33557_, _33556_, _33555_);
  and (_33558_, _33557_, _11659_);
  or (_33559_, _33558_, _33511_);
  nand (_33560_, _33559_, _03737_);
  and (_33561_, _11565_, _03729_);
  nor (_33562_, _33561_, _11668_);
  nand (_33563_, _33562_, _33560_);
  nor (_33564_, _33507_, _11666_);
  nor (_33566_, _33564_, _03714_);
  and (_33567_, _33566_, _33563_);
  or (_33568_, _33567_, _33509_);
  nand (_33569_, _33568_, _03233_);
  and (_33570_, _06236_, _11670_);
  nor (_33571_, _33570_, _03508_);
  nand (_33572_, _33571_, _33569_);
  and (_33573_, _11564_, _03508_);
  nor (_33574_, _33573_, _09917_);
  nand (_33575_, _33574_, _33572_);
  and (_33577_, _11430_, _09969_);
  not (_33578_, _33513_);
  nor (_33579_, _33578_, _09969_);
  or (_33580_, _33579_, _09921_);
  nor (_33581_, _33580_, _33577_);
  nor (_33582_, _33581_, _33232_);
  nand (_33583_, _33582_, _33575_);
  and (_33584_, _11430_, _09876_);
  nor (_33585_, _33578_, _09876_);
  nor (_33586_, _33585_, _33584_);
  nor (_33588_, _33586_, _04107_);
  and (_33589_, _33578_, _10018_);
  or (_33590_, _11430_, _10018_);
  nand (_33591_, _33590_, _09919_);
  nor (_33592_, _33591_, _33589_);
  nor (_33593_, _33592_, _33588_);
  nand (_33594_, _33593_, _33583_);
  nand (_33595_, _33594_, _09856_);
  and (_33596_, _11430_, _10061_);
  not (_33597_, _10061_);
  and (_33599_, _33513_, _33597_);
  or (_33600_, _33599_, _33596_);
  and (_33601_, _33600_, _03604_);
  nor (_33602_, _33601_, _10025_);
  and (_33603_, _33602_, _33595_);
  or (_33604_, _33603_, _33508_);
  nand (_33605_, _33604_, _06840_);
  and (_33606_, _11565_, _03719_);
  nor (_33607_, _33606_, _04766_);
  nand (_33608_, _33607_, _33605_);
  nor (_33610_, _06236_, _03227_);
  nor (_33611_, _33610_, _33264_);
  and (_33612_, _33611_, _33608_);
  or (_33613_, _33612_, _33502_);
  nand (_33614_, _33613_, _11355_);
  nor (_33615_, _33506_, _11355_);
  nor (_33616_, _33615_, _03753_);
  and (_33617_, _33616_, _33614_);
  and (_33618_, _11564_, _03753_);
  or (_33619_, _33618_, _33617_);
  and (_33621_, _33619_, _03238_);
  nor (_33622_, _06236_, _03238_);
  or (_33623_, _33622_, _03752_);
  or (_33624_, _33623_, _33621_);
  and (_33625_, _11565_, _03752_);
  not (_33626_, _33625_);
  and (_33627_, _33626_, _11350_);
  nand (_33628_, _33627_, _33624_);
  nor (_33629_, _33507_, _11350_);
  nor (_33630_, _33629_, _08187_);
  nand (_33632_, _33630_, _33628_);
  nor (_33633_, _11564_, _08186_);
  nor (_33634_, _33633_, _07912_);
  and (_33635_, _33634_, _33632_);
  nor (_33636_, _33507_, _03248_);
  or (_33637_, _33636_, _03505_);
  nor (_33638_, _33637_, _33635_);
  and (_33639_, _11565_, _03505_);
  or (_33640_, _33639_, _33638_);
  nand (_33641_, _33640_, _05897_);
  and (_33643_, _06236_, _03224_);
  nor (_33644_, _33643_, _03625_);
  nand (_33645_, _33644_, _33641_);
  and (_33646_, _11430_, _03625_);
  nor (_33647_, _33646_, _33299_);
  nand (_33648_, _33647_, _33645_);
  nor (_33649_, _11749_, _11564_);
  nor (_33650_, _33649_, _03222_);
  and (_33651_, _33650_, _33648_);
  and (_33652_, _11430_, _03222_);
  nor (_33654_, _33652_, _33651_);
  nand (_33655_, _33654_, _11756_);
  nor (_33656_, _33506_, _11756_);
  nor (_33657_, _33656_, _03585_);
  and (_33658_, _33657_, _33655_);
  and (_33659_, _11564_, _03585_);
  or (_33660_, _33659_, _03169_);
  or (_33661_, _33660_, _33658_);
  and (_33662_, _06236_, _03169_);
  nor (_33663_, _33662_, _11764_);
  nand (_33665_, _33663_, _33661_);
  and (_33666_, _33497_, _11764_);
  nor (_33667_, _33666_, _06168_);
  nand (_33668_, _33667_, _33665_);
  nor (_33669_, _11564_, _05894_);
  nor (_33670_, _33669_, _03601_);
  nand (_33671_, _33670_, _33668_);
  and (_33672_, _11430_, _03601_);
  nor (_33673_, _33672_, _08363_);
  nand (_33674_, _33673_, _33671_);
  and (_33676_, _11565_, _08363_);
  nor (_33677_, _33676_, _11347_);
  nand (_33678_, _33677_, _33674_);
  and (_33679_, _11795_, _11792_);
  nor (_33680_, _33679_, _11796_);
  and (_33681_, _33680_, _11347_);
  nor (_33682_, _33681_, _03584_);
  and (_33683_, _33682_, _33678_);
  and (_33684_, _11565_, _03584_);
  or (_33685_, _33684_, _33683_);
  nand (_33687_, _33685_, _10736_);
  and (_33688_, _06236_, _03178_);
  nor (_33689_, _33688_, _11819_);
  and (_33690_, _33689_, _33687_);
  or (_33691_, _33690_, _33501_);
  nand (_33692_, _33691_, _11345_);
  nor (_33693_, _33507_, _11345_);
  nor (_33694_, _33693_, _11342_);
  nand (_33695_, _33694_, _33692_);
  nor (_33696_, _11564_, _11341_);
  nor (_33698_, _33696_, _03600_);
  nand (_33699_, _33698_, _33695_);
  and (_33700_, _11430_, _03600_);
  nor (_33701_, _33700_, _03780_);
  and (_33702_, _33701_, _33699_);
  or (_33703_, _33702_, _33494_);
  nand (_33704_, _33703_, _32175_);
  and (_33705_, _06236_, _03182_);
  nor (_33706_, _33705_, _11841_);
  nand (_33707_, _33706_, _33704_);
  or (_33709_, _11565_, _08786_);
  nand (_33710_, _33497_, _08786_);
  and (_33711_, _33710_, _33709_);
  or (_33712_, _33711_, _11842_);
  nand (_33713_, _33712_, _33707_);
  nand (_33714_, _33713_, _11851_);
  nor (_33715_, _33507_, _11851_);
  nor (_33716_, _33715_, _08431_);
  nand (_33717_, _33716_, _33714_);
  nor (_33718_, _11564_, _08430_);
  nor (_33720_, _33718_, _03622_);
  nand (_33721_, _33720_, _33717_);
  and (_33722_, _11430_, _03622_);
  nor (_33723_, _33722_, _03790_);
  and (_33724_, _33723_, _33721_);
  and (_33725_, _11565_, _03790_);
  or (_33726_, _33725_, _33724_);
  nand (_33727_, _33726_, _32171_);
  and (_33728_, _06236_, _03192_);
  nor (_33729_, _33728_, _11337_);
  and (_33731_, _33729_, _33727_);
  and (_33732_, _11564_, \oc8051_golden_model_1.PSW [7]);
  and (_33733_, _33497_, _07871_);
  or (_33734_, _33733_, _33732_);
  and (_33735_, _33734_, _11337_);
  or (_33736_, _33735_, _33731_);
  nand (_33737_, _33736_, _11335_);
  nor (_33738_, _33507_, _11335_);
  nor (_33739_, _33738_, _08460_);
  nand (_33740_, _33739_, _33737_);
  nor (_33742_, _11564_, _08459_);
  nor (_33743_, _33742_, _03624_);
  nand (_33744_, _33743_, _33740_);
  and (_33745_, _11430_, _03624_);
  nor (_33746_, _33745_, _03785_);
  and (_33747_, _33746_, _33744_);
  and (_33748_, _11565_, _03785_);
  or (_33749_, _33748_, _33747_);
  nand (_33750_, _33749_, _32168_);
  and (_33751_, _06236_, _03201_);
  nor (_33753_, _33751_, _11880_);
  nand (_33754_, _33753_, _33750_);
  nand (_33755_, _11564_, _07871_);
  nand (_33756_, _33497_, \oc8051_golden_model_1.PSW [7]);
  and (_33757_, _33756_, _33755_);
  or (_33758_, _33757_, _11881_);
  nand (_33759_, _33758_, _33754_);
  nand (_33760_, _33759_, _11330_);
  nor (_33761_, _33507_, _11330_);
  nor (_33762_, _33761_, _08508_);
  nand (_33764_, _33762_, _33760_);
  nor (_33765_, _11564_, _08507_);
  nor (_33766_, _33765_, _08587_);
  nand (_33767_, _33766_, _33764_);
  and (_33768_, _33506_, _08587_);
  nor (_33769_, _33768_, _03798_);
  and (_33770_, _33769_, _33767_);
  nor (_33771_, _06730_, _10652_);
  or (_33772_, _33771_, _33770_);
  nand (_33773_, _33772_, _06399_);
  and (_33775_, _06236_, _03188_);
  nor (_33776_, _33775_, _03621_);
  and (_33777_, _33776_, _33773_);
  nor (_33778_, _11431_, _09854_);
  and (_33779_, _33513_, _09854_);
  nor (_33780_, _33779_, _33778_);
  nor (_33781_, _33780_, _11903_);
  or (_33782_, _33781_, _33777_);
  nand (_33783_, _33782_, _11328_);
  nor (_33784_, _33507_, _11328_);
  nor (_33785_, _33784_, _08703_);
  nand (_33786_, _33785_, _33783_);
  nor (_33787_, _11564_, _08702_);
  nor (_33788_, _33787_, _08732_);
  nand (_33789_, _33788_, _33786_);
  and (_33790_, _33506_, _08732_);
  nor (_33791_, _33790_, _03515_);
  nand (_33792_, _33791_, _33789_);
  nor (_33793_, _06730_, _03516_);
  nor (_33794_, _33793_, _03203_);
  nand (_33796_, _33794_, _33792_);
  nor (_33797_, _06236_, _32165_);
  nor (_33798_, _33797_, _03628_);
  nand (_33799_, _33798_, _33796_);
  and (_33800_, _11431_, _09854_);
  nor (_33801_, _33513_, _09854_);
  nor (_33802_, _33801_, _33800_);
  nor (_33803_, _33802_, _03816_);
  nor (_33804_, _33803_, _11934_);
  nand (_33805_, _33804_, _33799_);
  nor (_33807_, _33507_, _11933_);
  nor (_33808_, _33807_, _03815_);
  nand (_33809_, _33808_, _33805_);
  and (_33810_, _11565_, _03815_);
  nor (_33811_, _33810_, _32765_);
  nand (_33812_, _33811_, _33809_);
  nor (_33813_, _33507_, _11940_);
  nor (_33814_, _33813_, _05103_);
  and (_33815_, _33814_, _33812_);
  or (_33816_, _33815_, _33493_);
  nand (_33818_, _33816_, _03823_);
  nor (_33819_, _33802_, _03823_);
  nor (_33820_, _33819_, _11958_);
  nand (_33821_, _33820_, _33818_);
  nor (_33822_, _33507_, _11957_);
  nor (_33823_, _33822_, _03447_);
  nand (_33824_, _33823_, _33821_);
  not (_33825_, _11964_);
  and (_33826_, _11565_, _03447_);
  nor (_33827_, _33826_, _33825_);
  nand (_33829_, _33827_, _33824_);
  nor (_33830_, _33507_, _11964_);
  nor (_33831_, _33830_, _32154_);
  nand (_33832_, _33831_, _33829_);
  and (_33833_, _32154_, _06236_);
  nor (_33834_, _33833_, _11975_);
  and (_33835_, _33834_, _33832_);
  and (_33836_, _33506_, _11975_);
  or (_33837_, _33836_, _33835_);
  or (_33838_, _33837_, _43004_);
  or (_33840_, _43000_, \oc8051_golden_model_1.PC [4]);
  and (_33841_, _33840_, _41806_);
  and (_43673_, _33841_, _33838_);
  nor (_33842_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_33843_, _11559_, _02905_);
  nor (_33844_, _33843_, _33842_);
  and (_33845_, _33844_, _11975_);
  and (_33846_, _11559_, _03447_);
  nor (_33847_, _33844_, _11328_);
  nor (_33848_, _33844_, _11330_);
  nor (_33850_, _33844_, _11335_);
  nor (_33851_, _33844_, _11851_);
  nor (_33852_, _33844_, _11345_);
  and (_33853_, _11560_, _03584_);
  and (_33854_, _11560_, _03505_);
  nor (_33855_, _32547_, _11559_);
  and (_33856_, _11504_, _11560_);
  or (_33857_, _11562_, _11561_);
  and (_33858_, _33857_, _11587_);
  nor (_33859_, _33857_, _11587_);
  or (_33861_, _33859_, _33858_);
  and (_33862_, _33861_, _11624_);
  or (_33863_, _33862_, _06072_);
  or (_33864_, _33863_, _33856_);
  and (_33865_, _06267_, _03980_);
  nor (_33866_, _33844_, _11643_);
  and (_33867_, _11560_, _03979_);
  or (_33868_, _04409_, \oc8051_golden_model_1.PC [5]);
  nor (_33869_, _33868_, _04729_);
  or (_33870_, _33869_, _33867_);
  and (_33871_, _33870_, _32816_);
  or (_33872_, _33871_, _06073_);
  or (_33873_, _33872_, _33866_);
  or (_33874_, _33873_, _33865_);
  and (_33875_, _33874_, _33864_);
  nand (_33876_, _33875_, _05966_);
  not (_33877_, _33844_);
  and (_33878_, _33877_, _04422_);
  nor (_33879_, _33878_, _03610_);
  and (_33880_, _33879_, _33876_);
  or (_33883_, _11426_, _11367_);
  or (_33884_, _11428_, _11427_);
  and (_33885_, _33884_, _11460_);
  nor (_33886_, _33884_, _11460_);
  or (_33887_, _33886_, _33885_);
  or (_33888_, _33887_, _11369_);
  nand (_33889_, _33888_, _33883_);
  and (_33890_, _33889_, _03610_);
  nor (_33891_, _33890_, _33880_);
  nand (_33892_, _33891_, _11362_);
  nor (_33894_, _33844_, _11362_);
  nor (_33895_, _33894_, _03715_);
  nand (_33896_, _33895_, _33892_);
  and (_33897_, _11559_, _03715_);
  nor (_33898_, _33897_, _04768_);
  nand (_33899_, _33898_, _33896_);
  and (_33900_, _06267_, _04768_);
  nor (_33901_, _33900_, _03723_);
  nand (_33902_, _33901_, _33899_);
  and (_33903_, _11559_, _03723_);
  nor (_33905_, _33903_, _11660_);
  nand (_33906_, _33905_, _33902_);
  nor (_33907_, _33844_, _11659_);
  nor (_33908_, _33907_, _03729_);
  nand (_33909_, _33908_, _33906_);
  and (_33910_, _11559_, _03729_);
  nor (_33911_, _33910_, _11668_);
  nand (_33912_, _33911_, _33909_);
  nor (_33913_, _33844_, _11666_);
  nor (_33914_, _33913_, _03714_);
  nand (_33916_, _33914_, _33912_);
  and (_33917_, _11559_, _03714_);
  nor (_33918_, _33917_, _11670_);
  nand (_33919_, _33918_, _33916_);
  and (_33920_, _06267_, _11670_);
  nor (_33921_, _33920_, _03508_);
  nand (_33922_, _33921_, _33919_);
  and (_33923_, _11559_, _03508_);
  nor (_33924_, _33923_, _09917_);
  nand (_33925_, _33924_, _33922_);
  and (_33927_, _11425_, _09969_);
  not (_33928_, _33927_);
  nor (_33929_, _33887_, _09969_);
  nor (_33930_, _33929_, _09921_);
  and (_33931_, _33930_, _33928_);
  nor (_33932_, _33931_, _33232_);
  nand (_33933_, _33932_, _33925_);
  and (_33934_, _11425_, _09876_);
  nor (_33935_, _33887_, _09876_);
  nor (_33936_, _33935_, _33934_);
  nor (_33938_, _33936_, _04107_);
  or (_33939_, _11426_, _10018_);
  or (_33940_, _33887_, _11685_);
  nand (_33941_, _33940_, _33939_);
  and (_33942_, _33941_, _09919_);
  nor (_33943_, _33942_, _33938_);
  nand (_33944_, _33943_, _33933_);
  nand (_33945_, _33944_, _09856_);
  nand (_33946_, _11425_, _10061_);
  or (_33947_, _33887_, _10061_);
  and (_33949_, _33947_, _33946_);
  or (_33950_, _33949_, _09856_);
  and (_33951_, _33950_, _33945_);
  or (_33952_, _33951_, _10025_);
  nand (_33953_, _33844_, _10025_);
  and (_33954_, _33953_, _33952_);
  nand (_33955_, _33954_, _06840_);
  and (_33956_, _11560_, _03719_);
  nor (_33957_, _33956_, _04766_);
  nand (_33958_, _33957_, _33955_);
  nor (_33960_, _06267_, _03227_);
  nor (_33961_, _33960_, _33264_);
  and (_33962_, _33961_, _33958_);
  or (_33963_, _33962_, _33855_);
  nand (_33964_, _33963_, _11355_);
  nor (_33965_, _33844_, _11355_);
  nor (_33966_, _33965_, _03753_);
  nand (_33967_, _33966_, _33964_);
  and (_33968_, _11559_, _03753_);
  nor (_33969_, _33968_, _11727_);
  nand (_33971_, _33969_, _33967_);
  and (_33972_, _06267_, _11727_);
  nor (_33973_, _33972_, _03752_);
  nand (_33974_, _33973_, _33971_);
  and (_33975_, _11559_, _03752_);
  not (_33976_, _33975_);
  and (_33977_, _33976_, _11350_);
  and (_33978_, _33977_, _33974_);
  nor (_33979_, _33844_, _11350_);
  or (_33980_, _33979_, _33978_);
  nand (_33982_, _33980_, _08186_);
  nor (_33983_, _11559_, _08186_);
  nor (_33984_, _33983_, _07912_);
  nand (_33985_, _33984_, _33982_);
  nor (_33986_, _33877_, _03248_);
  nor (_33987_, _33986_, _03505_);
  and (_33988_, _33987_, _33985_);
  or (_33989_, _33988_, _33854_);
  nand (_33990_, _33989_, _05897_);
  and (_33991_, _06267_, _03224_);
  nor (_33993_, _33991_, _03625_);
  nand (_33994_, _33993_, _33990_);
  and (_33995_, _11425_, _03625_);
  nor (_33996_, _33995_, _33299_);
  nand (_33997_, _33996_, _33994_);
  nor (_33998_, _11749_, _11559_);
  nor (_33999_, _33998_, _03222_);
  nand (_34000_, _33999_, _33997_);
  and (_34001_, _11425_, _03222_);
  nor (_34002_, _34001_, _11758_);
  nand (_34004_, _34002_, _34000_);
  nor (_34005_, _33844_, _11756_);
  nor (_34006_, _34005_, _03585_);
  nand (_34007_, _34006_, _34004_);
  nor (_34008_, _11559_, _03169_);
  or (_34009_, _34008_, _11760_);
  nand (_34010_, _34009_, _34007_);
  and (_34011_, _06267_, _03169_);
  nor (_34012_, _34011_, _11764_);
  nand (_34013_, _34012_, _34010_);
  nor (_34015_, _33861_, _11765_);
  nor (_34016_, _34015_, _06168_);
  nand (_34017_, _34016_, _34013_);
  nor (_34018_, _11559_, _05894_);
  nor (_34019_, _34018_, _03601_);
  nand (_34020_, _34019_, _34017_);
  and (_34021_, _11425_, _03601_);
  nor (_34022_, _34021_, _08363_);
  nand (_34023_, _34022_, _34020_);
  and (_34024_, _11560_, _08363_);
  nor (_34026_, _34024_, _11347_);
  nand (_34027_, _34026_, _34023_);
  and (_34028_, _11797_, _11790_);
  not (_34029_, _34028_);
  nor (_34030_, _11798_, _11348_);
  and (_34031_, _34030_, _34029_);
  nor (_34032_, _34031_, _03584_);
  and (_34033_, _34032_, _34027_);
  or (_34034_, _34033_, _33853_);
  nand (_34035_, _34034_, _10736_);
  and (_34037_, _06267_, _03178_);
  nor (_34038_, _34037_, _11819_);
  nand (_34039_, _34038_, _34035_);
  and (_34040_, _11559_, _08786_);
  nor (_34041_, _33861_, _08786_);
  or (_34042_, _34041_, _34040_);
  and (_34043_, _34042_, _11819_);
  nor (_34044_, _34043_, _11824_);
  and (_34045_, _34044_, _34039_);
  or (_34046_, _34045_, _33852_);
  nand (_34048_, _34046_, _11341_);
  nor (_34049_, _11559_, _11341_);
  nor (_34050_, _34049_, _03600_);
  and (_34051_, _34050_, _34048_);
  and (_34052_, _11425_, _03600_);
  or (_34053_, _34052_, _03780_);
  nor (_34054_, _34053_, _34051_);
  and (_34055_, _11560_, _03780_);
  or (_34056_, _34055_, _34054_);
  nand (_34057_, _34056_, _32175_);
  and (_34059_, _06267_, _03182_);
  nor (_34060_, _34059_, _11841_);
  nand (_34061_, _34060_, _34057_);
  nand (_34062_, _33861_, _08786_);
  or (_34063_, _11559_, _08786_);
  and (_34064_, _34063_, _11841_);
  and (_34065_, _34064_, _34062_);
  nor (_34066_, _34065_, _11853_);
  and (_34067_, _34066_, _34061_);
  or (_34068_, _34067_, _33851_);
  nand (_34070_, _34068_, _08430_);
  nor (_34071_, _11559_, _08430_);
  nor (_34072_, _34071_, _03622_);
  and (_34073_, _34072_, _34070_);
  and (_34074_, _11425_, _03622_);
  or (_34075_, _34074_, _03790_);
  nor (_34076_, _34075_, _34073_);
  and (_34077_, _11560_, _03790_);
  or (_34078_, _34077_, _34076_);
  nand (_34079_, _34078_, _32171_);
  and (_34081_, _06267_, _03192_);
  nor (_34082_, _34081_, _11337_);
  nand (_34083_, _34082_, _34079_);
  and (_34084_, _33861_, _07871_);
  nor (_34085_, _11559_, _07871_);
  nor (_34086_, _34085_, _11338_);
  not (_34087_, _34086_);
  nor (_34088_, _34087_, _34084_);
  nor (_34089_, _34088_, _11864_);
  and (_34090_, _34089_, _34083_);
  or (_34092_, _34090_, _33850_);
  nand (_34093_, _34092_, _08459_);
  nor (_34094_, _11559_, _08459_);
  nor (_34095_, _34094_, _03624_);
  and (_34096_, _34095_, _34093_);
  and (_34097_, _11425_, _03624_);
  or (_34098_, _34097_, _03785_);
  nor (_34099_, _34098_, _34096_);
  and (_34100_, _11560_, _03785_);
  or (_34101_, _34100_, _34099_);
  nand (_34103_, _34101_, _32168_);
  and (_34104_, _06267_, _03201_);
  nor (_34105_, _34104_, _11880_);
  nand (_34106_, _34105_, _34103_);
  and (_34107_, _33861_, \oc8051_golden_model_1.PSW [7]);
  nor (_34108_, _11559_, \oc8051_golden_model_1.PSW [7]);
  nor (_34109_, _34108_, _11881_);
  not (_34110_, _34109_);
  nor (_34111_, _34110_, _34107_);
  nor (_34112_, _34111_, _11885_);
  and (_34114_, _34112_, _34106_);
  or (_34115_, _34114_, _33848_);
  nand (_34116_, _34115_, _08507_);
  nor (_34117_, _11559_, _08507_);
  nor (_34118_, _34117_, _08587_);
  nand (_34119_, _34118_, _34116_);
  and (_34120_, _33844_, _08587_);
  nor (_34121_, _34120_, _03798_);
  and (_34122_, _34121_, _34119_);
  nor (_34123_, _06684_, _10652_);
  or (_34125_, _34123_, _34122_);
  nand (_34126_, _34125_, _06399_);
  and (_34127_, _06267_, _03188_);
  nor (_34128_, _34127_, _03621_);
  nand (_34129_, _34128_, _34126_);
  and (_34130_, _33887_, _09854_);
  nor (_34131_, _11425_, _09854_);
  or (_34132_, _34131_, _11903_);
  or (_34133_, _34132_, _34130_);
  and (_34134_, _34133_, _11328_);
  and (_34136_, _34134_, _34129_);
  or (_34137_, _34136_, _33847_);
  nand (_34138_, _34137_, _08702_);
  nor (_34139_, _11559_, _08702_);
  nor (_34140_, _34139_, _08732_);
  nand (_34141_, _34140_, _34138_);
  and (_34142_, _33844_, _08732_);
  nor (_34143_, _34142_, _03515_);
  and (_34144_, _34143_, _34141_);
  nor (_34145_, _06684_, _03516_);
  or (_34146_, _34145_, _34144_);
  nand (_34147_, _34146_, _32165_);
  and (_34148_, _06267_, _03203_);
  nor (_34149_, _34148_, _03628_);
  nand (_34150_, _34149_, _34147_);
  and (_34151_, _11425_, _09854_);
  nor (_34152_, _33887_, _09854_);
  or (_34153_, _34152_, _34151_);
  and (_34154_, _34153_, _03628_);
  nor (_34155_, _34154_, _11934_);
  nand (_34158_, _34155_, _34150_);
  nor (_34159_, _33844_, _11933_);
  nor (_34160_, _34159_, _03815_);
  nand (_34161_, _34160_, _34158_);
  and (_34162_, _11559_, _03815_);
  nor (_34163_, _34162_, _32765_);
  and (_34164_, _34163_, _34161_);
  nor (_34165_, _33844_, _11940_);
  or (_34166_, _34165_, _34164_);
  nand (_34167_, _34166_, _04540_);
  and (_34169_, _06267_, _05103_);
  nor (_34170_, _34169_, _03453_);
  nand (_34171_, _34170_, _34167_);
  and (_34172_, _34153_, _03453_);
  nor (_34173_, _34172_, _11958_);
  nand (_34174_, _34173_, _34171_);
  nor (_34175_, _33844_, _11957_);
  nor (_34176_, _34175_, _03447_);
  and (_34177_, _34176_, _34174_);
  or (_34178_, _34177_, _33846_);
  nand (_34180_, _34178_, _11964_);
  nor (_34181_, _33877_, _11964_);
  nor (_34182_, _34181_, _32154_);
  nand (_34183_, _34182_, _34180_);
  and (_34184_, _32154_, _06267_);
  nor (_34185_, _34184_, _11975_);
  and (_34186_, _34185_, _34183_);
  or (_34187_, _34186_, _33845_);
  or (_34188_, _34187_, _43004_);
  or (_34189_, _43000_, \oc8051_golden_model_1.PC [5]);
  and (_34191_, _34189_, _41806_);
  and (_43674_, _34191_, _34188_);
  and (_34192_, _06204_, _05103_);
  and (_34193_, _06077_, _11315_);
  nor (_34194_, _34193_, \oc8051_golden_model_1.PC [6]);
  nor (_34195_, _34194_, _11316_);
  not (_34196_, _34195_);
  and (_34197_, _34196_, _08732_);
  and (_34198_, _11418_, _03624_);
  and (_34199_, _11418_, _03622_);
  and (_34201_, _11418_, _03600_);
  nor (_34202_, _34196_, _11350_);
  and (_34203_, _11552_, _03714_);
  nor (_34204_, _34195_, _11653_);
  and (_34205_, _06204_, _03980_);
  nor (_34206_, _04729_, \oc8051_golden_model_1.PC [6]);
  or (_34207_, _34206_, _04409_);
  and (_34208_, _11551_, _04409_);
  nor (_34209_, _34208_, _11632_);
  and (_34210_, _34209_, _34207_);
  or (_34212_, _34195_, _11642_);
  nand (_34213_, _34212_, _11630_);
  or (_34214_, _34213_, _34210_);
  and (_34215_, _34214_, _04763_);
  nor (_34216_, _34215_, _34205_);
  nor (_34217_, _34196_, _11630_);
  nor (_34218_, _34217_, _06073_);
  not (_34219_, _34218_);
  nor (_34220_, _34219_, _34216_);
  and (_34221_, _11589_, _11556_);
  nor (_34223_, _34221_, _11590_);
  nand (_34224_, _34223_, _11624_);
  or (_34225_, _11624_, _11552_);
  and (_34226_, _34225_, _06073_);
  and (_34227_, _34226_, _34224_);
  or (_34228_, _34227_, _34220_);
  nand (_34229_, _34228_, _11647_);
  or (_34230_, _11418_, _11367_);
  and (_34231_, _11462_, _11422_);
  nor (_34232_, _34231_, _11463_);
  not (_34234_, _34232_);
  or (_34235_, _34234_, _11369_);
  and (_34236_, _34235_, _03610_);
  nand (_34237_, _34236_, _34230_);
  nand (_34238_, _34237_, _34229_);
  and (_34239_, _34238_, _11362_);
  or (_34240_, _34239_, _34204_);
  nand (_34241_, _34240_, _04055_);
  and (_34242_, _11552_, _03715_);
  nor (_34243_, _34242_, _04768_);
  and (_34245_, _34243_, _34241_);
  nor (_34246_, _06204_, _03230_);
  or (_34247_, _34246_, _03723_);
  nor (_34248_, _34247_, _34245_);
  and (_34249_, _11552_, _03723_);
  or (_34250_, _34249_, _34248_);
  and (_34251_, _34250_, _11659_);
  nor (_34252_, _34195_, _11659_);
  or (_34253_, _34252_, _34251_);
  nand (_34254_, _34253_, _03737_);
  and (_34256_, _11552_, _03729_);
  nor (_34257_, _34256_, _11668_);
  nand (_34258_, _34257_, _34254_);
  nor (_34259_, _34196_, _11666_);
  nor (_34260_, _34259_, _03714_);
  and (_34261_, _34260_, _34258_);
  or (_34262_, _34261_, _34203_);
  nand (_34263_, _34262_, _03233_);
  and (_34264_, _06204_, _11670_);
  nor (_34265_, _34264_, _03508_);
  nand (_34267_, _34265_, _34263_);
  and (_34268_, _11551_, _03508_);
  nor (_34269_, _34268_, _09917_);
  nand (_34270_, _34269_, _34267_);
  and (_34271_, _11417_, _09969_);
  nor (_34272_, _34234_, _09969_);
  or (_34273_, _34272_, _09921_);
  nor (_34274_, _34273_, _34271_);
  nor (_34275_, _34274_, _33232_);
  and (_34276_, _34275_, _34270_);
  and (_34278_, _34234_, _10018_);
  and (_34279_, _11418_, _11685_);
  nor (_34280_, _34279_, _34278_);
  and (_34281_, _34280_, _32519_);
  nor (_34282_, _34281_, _34276_);
  and (_34283_, _11418_, _09876_);
  nor (_34284_, _34232_, _09876_);
  or (_34285_, _34284_, _04107_);
  or (_34286_, _34285_, _34283_);
  nand (_34287_, _34286_, _34282_);
  nand (_34289_, _34287_, _09856_);
  nand (_34290_, _11417_, _10061_);
  nand (_34291_, _34232_, _33597_);
  and (_34292_, _34291_, _34290_);
  or (_34293_, _34292_, _09856_);
  and (_34294_, _34293_, _34289_);
  or (_34295_, _34294_, _10025_);
  nand (_34296_, _34195_, _10025_);
  and (_34297_, _34296_, _34295_);
  nand (_34298_, _34297_, _06840_);
  and (_34300_, _11552_, _03719_);
  nor (_34301_, _34300_, _04766_);
  nand (_34302_, _34301_, _34298_);
  nor (_34303_, _06204_, _03227_);
  nor (_34304_, _34303_, _33264_);
  and (_34305_, _34304_, _34302_);
  nor (_34306_, _32547_, _11551_);
  or (_34307_, _34306_, _34305_);
  nand (_34308_, _34307_, _11355_);
  nor (_34309_, _34195_, _11355_);
  nor (_34311_, _34309_, _03753_);
  and (_34312_, _34311_, _34308_);
  and (_34313_, _11551_, _03753_);
  or (_34314_, _34313_, _34312_);
  and (_34315_, _34314_, _03238_);
  nor (_34316_, _06204_, _03238_);
  or (_34317_, _34316_, _03752_);
  or (_34318_, _34317_, _34315_);
  and (_34319_, _11552_, _03752_);
  not (_34320_, _34319_);
  and (_34322_, _34320_, _11350_);
  and (_34323_, _34322_, _34318_);
  or (_34324_, _34323_, _34202_);
  and (_34325_, _34324_, _08186_);
  nor (_34326_, _11552_, _08186_);
  or (_34327_, _34326_, _34325_);
  and (_34328_, _34327_, _03248_);
  nor (_34329_, _34196_, _03248_);
  or (_34330_, _34329_, _03505_);
  or (_34331_, _34330_, _34328_);
  and (_34333_, _11552_, _03505_);
  nor (_34334_, _34333_, _03224_);
  nand (_34335_, _34334_, _34331_);
  nor (_34336_, _06204_, _05897_);
  nor (_34337_, _34336_, _03625_);
  nand (_34338_, _34337_, _34335_);
  and (_34339_, _11418_, _03625_);
  nor (_34340_, _34339_, _33299_);
  nand (_34341_, _34340_, _34338_);
  nor (_34342_, _11749_, _11552_);
  nor (_34344_, _34342_, _03222_);
  nand (_34345_, _34344_, _34341_);
  and (_34346_, _11418_, _03222_);
  nor (_34347_, _34346_, _11758_);
  nand (_34348_, _34347_, _34345_);
  nor (_34349_, _34196_, _11756_);
  nor (_34350_, _34349_, _03585_);
  nand (_34351_, _34350_, _34348_);
  and (_34352_, _11552_, _03585_);
  nor (_34353_, _34352_, _03169_);
  and (_34355_, _34353_, _34351_);
  nor (_34356_, _06204_, _03170_);
  or (_34357_, _34356_, _34355_);
  and (_34358_, _34357_, _11765_);
  and (_34359_, _34223_, _11764_);
  or (_34360_, _34359_, _34358_);
  nand (_34361_, _34360_, _05894_);
  nor (_34362_, _11552_, _05894_);
  nor (_34363_, _34362_, _03601_);
  nand (_34364_, _34363_, _34361_);
  and (_34366_, _11418_, _03601_);
  nor (_34367_, _34366_, _08363_);
  nand (_34368_, _34367_, _34364_);
  and (_34369_, _11551_, _08363_);
  nor (_34370_, _34369_, _11347_);
  nand (_34371_, _34370_, _34368_);
  and (_34372_, _11799_, _11786_);
  nor (_34373_, _34372_, _11800_);
  nor (_34374_, _34373_, _11348_);
  nor (_34375_, _34374_, _03584_);
  nand (_34377_, _34375_, _34371_);
  and (_34378_, _11551_, _03584_);
  nor (_34379_, _34378_, _03178_);
  nand (_34380_, _34379_, _34377_);
  and (_34381_, _06204_, _03178_);
  nor (_34382_, _34381_, _11819_);
  nand (_34383_, _34382_, _34380_);
  and (_34384_, _11551_, _08786_);
  and (_34385_, _34223_, _11826_);
  or (_34386_, _34385_, _34384_);
  and (_34388_, _34386_, _11819_);
  nor (_34389_, _34388_, _11824_);
  nand (_34390_, _34389_, _34383_);
  nor (_34391_, _34195_, _11345_);
  nor (_34392_, _34391_, _11342_);
  nand (_34393_, _34392_, _34390_);
  nor (_34394_, _11552_, _11341_);
  nor (_34395_, _34394_, _03600_);
  and (_34396_, _34395_, _34393_);
  or (_34397_, _34396_, _34201_);
  nand (_34399_, _34397_, _07778_);
  and (_34400_, _11552_, _03780_);
  nor (_34401_, _34400_, _03182_);
  and (_34402_, _34401_, _34399_);
  nor (_34403_, _06204_, _32175_);
  or (_34404_, _34403_, _34402_);
  nand (_34405_, _34404_, _11842_);
  or (_34406_, _34223_, _11826_);
  or (_34407_, _11551_, _08786_);
  and (_34408_, _34407_, _11841_);
  and (_34410_, _34408_, _34406_);
  nor (_34411_, _34410_, _11853_);
  nand (_34412_, _34411_, _34405_);
  nor (_34413_, _34195_, _11851_);
  nor (_34414_, _34413_, _08431_);
  nand (_34415_, _34414_, _34412_);
  nor (_34416_, _11552_, _08430_);
  nor (_34417_, _34416_, _03622_);
  and (_34418_, _34417_, _34415_);
  or (_34419_, _34418_, _34199_);
  nand (_34421_, _34419_, _06828_);
  and (_34422_, _11552_, _03790_);
  nor (_34423_, _34422_, _03192_);
  and (_34424_, _34423_, _34421_);
  nor (_34425_, _06204_, _32171_);
  or (_34426_, _34425_, _34424_);
  nand (_34427_, _34426_, _11338_);
  and (_34428_, _11551_, \oc8051_golden_model_1.PSW [7]);
  and (_34429_, _34223_, _07871_);
  or (_34430_, _34429_, _34428_);
  and (_34432_, _34430_, _11337_);
  nor (_34433_, _34432_, _11864_);
  nand (_34434_, _34433_, _34427_);
  nor (_34435_, _34195_, _11335_);
  nor (_34436_, _34435_, _08460_);
  nand (_34437_, _34436_, _34434_);
  nor (_34438_, _11552_, _08459_);
  nor (_34439_, _34438_, _03624_);
  and (_34440_, _34439_, _34437_);
  or (_34441_, _34440_, _34198_);
  nand (_34443_, _34441_, _07793_);
  and (_34444_, _11552_, _03785_);
  nor (_34445_, _34444_, _03201_);
  and (_34446_, _34445_, _34443_);
  nor (_34447_, _06204_, _32168_);
  or (_34448_, _34447_, _34446_);
  nand (_34449_, _34448_, _11881_);
  nor (_34450_, _34223_, _07871_);
  nor (_34451_, _11551_, \oc8051_golden_model_1.PSW [7]);
  nor (_34452_, _34451_, _11881_);
  not (_34454_, _34452_);
  nor (_34455_, _34454_, _34450_);
  nor (_34456_, _34455_, _11885_);
  nand (_34457_, _34456_, _34449_);
  nor (_34458_, _34195_, _11330_);
  nor (_34459_, _34458_, _08508_);
  nand (_34460_, _34459_, _34457_);
  nor (_34461_, _11552_, _08507_);
  nor (_34462_, _34461_, _08587_);
  nand (_34463_, _34462_, _34460_);
  and (_34465_, _34196_, _08587_);
  nor (_34466_, _34465_, _03798_);
  nand (_34467_, _34466_, _34463_);
  and (_34468_, _06455_, _03798_);
  nor (_34469_, _34468_, _03188_);
  nand (_34470_, _34469_, _34467_);
  and (_34471_, _06204_, _03188_);
  nor (_34472_, _34471_, _03621_);
  nand (_34473_, _34472_, _34470_);
  nor (_34474_, _11417_, _09854_);
  and (_34476_, _34234_, _09854_);
  or (_34477_, _34476_, _11903_);
  nor (_34478_, _34477_, _34474_);
  nor (_34479_, _34478_, _11907_);
  nand (_34480_, _34479_, _34473_);
  nor (_34481_, _34195_, _11328_);
  nor (_34482_, _34481_, _08703_);
  nand (_34483_, _34482_, _34480_);
  nor (_34484_, _11552_, _08702_);
  nor (_34485_, _34484_, _08732_);
  and (_34487_, _34485_, _34483_);
  or (_34488_, _34487_, _34197_);
  nand (_34489_, _34488_, _03516_);
  nor (_34490_, _06455_, _03516_);
  nor (_34491_, _34490_, _03203_);
  nand (_34492_, _34491_, _34489_);
  nor (_34493_, _06204_, _32165_);
  nor (_34494_, _34493_, _03628_);
  and (_34495_, _34494_, _34492_);
  nor (_34496_, _34232_, _09854_);
  and (_34498_, _11418_, _09854_);
  nor (_34499_, _34498_, _34496_);
  nor (_34500_, _34499_, _03816_);
  or (_34501_, _34500_, _34495_);
  and (_34502_, _34501_, _11933_);
  nor (_34503_, _34195_, _11933_);
  or (_34504_, _34503_, _34502_);
  nand (_34505_, _34504_, _04246_);
  and (_34506_, _11552_, _03815_);
  nor (_34507_, _34506_, _32765_);
  nand (_34509_, _34507_, _34505_);
  nor (_34510_, _34196_, _11940_);
  nor (_34511_, _34510_, _05103_);
  and (_34512_, _34511_, _34509_);
  or (_34513_, _34512_, _34192_);
  nand (_34514_, _34513_, _03823_);
  nor (_34515_, _34499_, _03823_);
  nor (_34516_, _34515_, _11958_);
  nand (_34517_, _34516_, _34514_);
  nor (_34518_, _34196_, _11957_);
  nor (_34520_, _34518_, _03447_);
  nand (_34521_, _34520_, _34517_);
  and (_34522_, _11552_, _03447_);
  nor (_34523_, _34522_, _33825_);
  nand (_34524_, _34523_, _34521_);
  nor (_34525_, _34196_, _11964_);
  nor (_34526_, _34525_, _32154_);
  nand (_34527_, _34526_, _34524_);
  and (_34528_, _32154_, _06204_);
  nor (_34529_, _34528_, _11975_);
  and (_34531_, _34529_, _34527_);
  and (_34532_, _34195_, _11975_);
  or (_34533_, _34532_, _34531_);
  or (_34534_, _34533_, _43004_);
  or (_34535_, _43000_, \oc8051_golden_model_1.PC [6]);
  and (_34536_, _34535_, _41806_);
  and (_43675_, _34536_, _34534_);
  and (_34537_, _06082_, _03447_);
  and (_34538_, _06082_, _03815_);
  nor (_34539_, _11316_, \oc8051_golden_model_1.PC [7]);
  nor (_34541_, _34539_, _11317_);
  nor (_34542_, _34541_, _11328_);
  nor (_34543_, _34541_, _11330_);
  nor (_34544_, _34541_, _11335_);
  nor (_34545_, _34541_, _11851_);
  nor (_34546_, _34541_, _11345_);
  and (_34547_, _06143_, _03505_);
  nor (_34548_, _34541_, _11350_);
  nor (_34549_, _32547_, _06082_);
  not (_34550_, _34541_);
  and (_34552_, _34550_, _10025_);
  and (_34553_, _11504_, _06143_);
  or (_34554_, _11547_, _11548_);
  and (_34555_, _34554_, _11591_);
  nor (_34556_, _34554_, _11591_);
  nor (_34557_, _34556_, _34555_);
  not (_34558_, _34557_);
  and (_34559_, _34558_, _11624_);
  or (_34560_, _34559_, _06072_);
  or (_34561_, _34560_, _34553_);
  and (_34563_, _05881_, _03980_);
  nor (_34564_, _34541_, _11642_);
  and (_34565_, _06143_, _03979_);
  nor (_34566_, _04409_, \oc8051_golden_model_1.PC [7]);
  and (_34567_, _34566_, _33169_);
  nor (_34568_, _34567_, _34565_);
  nor (_34569_, _34568_, _11632_);
  nor (_34570_, _34569_, _34564_);
  nor (_34571_, _34570_, _32191_);
  nor (_34572_, _34541_, _11630_);
  or (_34574_, _34572_, _06073_);
  or (_34575_, _34574_, _34571_);
  or (_34576_, _34575_, _34563_);
  and (_34577_, _34576_, _34561_);
  nand (_34578_, _34577_, _05966_);
  and (_34579_, _34550_, _04422_);
  nor (_34580_, _34579_, _03610_);
  and (_34581_, _34580_, _34578_);
  or (_34582_, _11367_, _06749_);
  or (_34583_, _11413_, _11414_);
  and (_34585_, _34583_, _11464_);
  nor (_34586_, _34583_, _11464_);
  nor (_34587_, _34586_, _34585_);
  not (_34588_, _34587_);
  or (_34589_, _34588_, _11369_);
  nand (_34590_, _34589_, _34582_);
  and (_34591_, _34590_, _03610_);
  nor (_34592_, _34591_, _34581_);
  nand (_34593_, _34592_, _11362_);
  nor (_34594_, _34541_, _11362_);
  nor (_34596_, _34594_, _03715_);
  nand (_34597_, _34596_, _34593_);
  and (_34598_, _06082_, _03715_);
  nor (_34599_, _34598_, _04768_);
  nand (_34600_, _34599_, _34597_);
  and (_34601_, _05881_, _04768_);
  nor (_34602_, _34601_, _03723_);
  nand (_34603_, _34602_, _34600_);
  and (_34604_, _06082_, _03723_);
  nor (_34605_, _34604_, _11660_);
  nand (_34607_, _34605_, _34603_);
  nor (_34608_, _34541_, _11659_);
  nor (_34609_, _34608_, _03729_);
  nand (_34610_, _34609_, _34607_);
  and (_34611_, _06082_, _03729_);
  nor (_34612_, _34611_, _11668_);
  nand (_34613_, _34612_, _34610_);
  nor (_34614_, _34541_, _11666_);
  nor (_34615_, _34614_, _03714_);
  nand (_34616_, _34615_, _34613_);
  and (_34618_, _06082_, _03714_);
  nor (_34619_, _34618_, _11670_);
  nand (_34620_, _34619_, _34616_);
  and (_34621_, _05881_, _11670_);
  nor (_34622_, _34621_, _03508_);
  nand (_34623_, _34622_, _34620_);
  and (_34624_, _06082_, _03508_);
  nor (_34625_, _34624_, _09917_);
  nand (_34626_, _34625_, _34623_);
  and (_34627_, _09969_, _06748_);
  nor (_34629_, _34588_, _09969_);
  or (_34630_, _34629_, _34627_);
  nor (_34631_, _34630_, _09921_);
  nor (_34632_, _34631_, _09919_);
  nand (_34633_, _34632_, _34626_);
  or (_34634_, _10018_, _06749_);
  or (_34635_, _34588_, _11685_);
  nand (_34636_, _34635_, _34634_);
  nand (_34637_, _34636_, _32519_);
  and (_34638_, _34637_, _34633_);
  or (_34640_, _34638_, _03615_);
  and (_34641_, _09876_, _06748_);
  nor (_34642_, _34588_, _09876_);
  nor (_34643_, _34642_, _34641_);
  or (_34644_, _34643_, _04107_);
  and (_34645_, _34644_, _34640_);
  or (_34646_, _34645_, _03604_);
  and (_34647_, _10061_, _06749_);
  nor (_34648_, _34587_, _10061_);
  or (_34649_, _34648_, _09856_);
  or (_34651_, _34649_, _34647_);
  and (_34652_, _34651_, _11358_);
  and (_34653_, _34652_, _34646_);
  or (_34654_, _34653_, _34552_);
  nand (_34655_, _34654_, _06840_);
  and (_34656_, _06143_, _03719_);
  nor (_34657_, _34656_, _04766_);
  nand (_34658_, _34657_, _34655_);
  nor (_34659_, _05881_, _03227_);
  nor (_34660_, _34659_, _33264_);
  and (_34662_, _34660_, _34658_);
  or (_34663_, _34662_, _34549_);
  nand (_34664_, _34663_, _11355_);
  nor (_34665_, _34541_, _11355_);
  nor (_34666_, _34665_, _03753_);
  nand (_34667_, _34666_, _34664_);
  and (_34668_, _06082_, _03753_);
  nor (_34669_, _34668_, _11727_);
  nand (_34670_, _34669_, _34667_);
  and (_34671_, _05881_, _11727_);
  nor (_34673_, _34671_, _03752_);
  nand (_34674_, _34673_, _34670_);
  and (_34675_, _06082_, _03752_);
  not (_34676_, _34675_);
  and (_34677_, _34676_, _11350_);
  and (_34678_, _34677_, _34674_);
  or (_34679_, _34678_, _34548_);
  nand (_34680_, _34679_, _08186_);
  nor (_34681_, _08186_, _06082_);
  nor (_34682_, _34681_, _07912_);
  nand (_34684_, _34682_, _34680_);
  nor (_34685_, _34550_, _03248_);
  nor (_34686_, _34685_, _03505_);
  and (_34687_, _34686_, _34684_);
  or (_34688_, _34687_, _34547_);
  nand (_34689_, _34688_, _05897_);
  and (_34690_, _05881_, _03224_);
  nor (_34691_, _34690_, _03625_);
  nand (_34692_, _34691_, _34689_);
  and (_34693_, _06748_, _03625_);
  nor (_34695_, _34693_, _33299_);
  nand (_34696_, _34695_, _34692_);
  nor (_34697_, _11749_, _06082_);
  nor (_34698_, _34697_, _03222_);
  nand (_34699_, _34698_, _34696_);
  and (_34700_, _06748_, _03222_);
  nor (_34701_, _34700_, _11758_);
  nand (_34702_, _34701_, _34699_);
  nor (_34703_, _34541_, _11756_);
  nor (_34704_, _34703_, _03585_);
  nand (_34706_, _34704_, _34702_);
  nor (_34707_, _06082_, _03169_);
  or (_34708_, _34707_, _11760_);
  nand (_34709_, _34708_, _34706_);
  and (_34710_, _05881_, _03169_);
  nor (_34711_, _34710_, _11764_);
  nand (_34712_, _34711_, _34709_);
  and (_34713_, _34557_, _11764_);
  nor (_34714_, _34713_, _06168_);
  nand (_34715_, _34714_, _34712_);
  nor (_34717_, _06082_, _05894_);
  nor (_34718_, _34717_, _03601_);
  nand (_34719_, _34718_, _34715_);
  and (_34720_, _06748_, _03601_);
  nor (_34721_, _34720_, _08363_);
  nand (_34722_, _34721_, _34719_);
  and (_34723_, _08363_, _06143_);
  nor (_34724_, _34723_, _11347_);
  nand (_34725_, _34724_, _34722_);
  or (_34726_, _11781_, _11782_);
  and (_34728_, _34726_, _11801_);
  nor (_34729_, _34726_, _11801_);
  or (_34730_, _34729_, _34728_);
  nor (_34731_, _34730_, _11348_);
  nor (_34732_, _34731_, _03584_);
  and (_34733_, _34732_, _34725_);
  and (_34734_, _06143_, _03584_);
  or (_34735_, _34734_, _34733_);
  nand (_34736_, _34735_, _10736_);
  and (_34737_, _05881_, _03178_);
  nor (_34739_, _34737_, _11819_);
  nand (_34740_, _34739_, _34736_);
  and (_34741_, _08786_, _06082_);
  and (_34742_, _34557_, _11826_);
  or (_34743_, _34742_, _34741_);
  and (_34744_, _34743_, _11819_);
  nor (_34745_, _34744_, _11824_);
  and (_34746_, _34745_, _34740_);
  or (_34747_, _34746_, _34546_);
  nand (_34748_, _34747_, _11341_);
  nor (_34750_, _11341_, _06082_);
  nor (_34751_, _34750_, _03600_);
  and (_34752_, _34751_, _34748_);
  and (_34753_, _06748_, _03600_);
  or (_34754_, _34753_, _03780_);
  nor (_34755_, _34754_, _34752_);
  and (_34756_, _06143_, _03780_);
  or (_34757_, _34756_, _34755_);
  nand (_34758_, _34757_, _32175_);
  and (_34759_, _05881_, _03182_);
  nor (_34761_, _34759_, _11841_);
  nand (_34762_, _34761_, _34758_);
  or (_34763_, _34557_, _11826_);
  or (_34764_, _08786_, _06082_);
  and (_34765_, _34764_, _11841_);
  and (_34766_, _34765_, _34763_);
  nor (_34767_, _34766_, _11853_);
  and (_34768_, _34767_, _34762_);
  or (_34769_, _34768_, _34545_);
  nand (_34770_, _34769_, _08430_);
  nor (_34771_, _08430_, _06082_);
  nor (_34772_, _34771_, _03622_);
  and (_34773_, _34772_, _34770_);
  and (_34774_, _06748_, _03622_);
  or (_34775_, _34774_, _03790_);
  nor (_34776_, _34775_, _34773_);
  and (_34777_, _06143_, _03790_);
  or (_34778_, _34777_, _34776_);
  nand (_34779_, _34778_, _32171_);
  and (_34780_, _05881_, _03192_);
  nor (_34783_, _34780_, _11337_);
  nand (_34784_, _34783_, _34779_);
  and (_34785_, _06082_, \oc8051_golden_model_1.PSW [7]);
  and (_34786_, _34557_, _07871_);
  or (_34787_, _34786_, _34785_);
  and (_34788_, _34787_, _11337_);
  nor (_34789_, _34788_, _11864_);
  and (_34790_, _34789_, _34784_);
  or (_34791_, _34790_, _34544_);
  nand (_34792_, _34791_, _08459_);
  nor (_34794_, _08459_, _06082_);
  nor (_34795_, _34794_, _03624_);
  and (_34796_, _34795_, _34792_);
  and (_34797_, _06748_, _03624_);
  or (_34798_, _34797_, _03785_);
  nor (_34799_, _34798_, _34796_);
  and (_34800_, _06143_, _03785_);
  or (_34801_, _34800_, _34799_);
  nand (_34802_, _34801_, _32168_);
  and (_34803_, _05881_, _03201_);
  nor (_34805_, _34803_, _11880_);
  nand (_34806_, _34805_, _34802_);
  nor (_34807_, _34557_, _07871_);
  nor (_34808_, _06082_, \oc8051_golden_model_1.PSW [7]);
  nor (_34809_, _34808_, _11881_);
  not (_34810_, _34809_);
  nor (_34811_, _34810_, _34807_);
  nor (_34812_, _34811_, _11885_);
  and (_34813_, _34812_, _34806_);
  or (_34814_, _34813_, _34543_);
  nand (_34816_, _34814_, _08507_);
  nor (_34817_, _08507_, _06082_);
  nor (_34818_, _34817_, _08587_);
  nand (_34819_, _34818_, _34816_);
  and (_34820_, _34541_, _08587_);
  nor (_34821_, _34820_, _03798_);
  and (_34822_, _34821_, _34819_);
  nor (_34823_, _06069_, _10652_);
  or (_34824_, _34823_, _34822_);
  nand (_34825_, _34824_, _06399_);
  and (_34827_, _05881_, _03188_);
  nor (_34828_, _34827_, _03621_);
  nand (_34829_, _34828_, _34825_);
  and (_34830_, _34588_, _09854_);
  nor (_34831_, _09854_, _06748_);
  or (_34832_, _34831_, _11903_);
  or (_34833_, _34832_, _34830_);
  and (_34834_, _34833_, _11328_);
  and (_34835_, _34834_, _34829_);
  or (_34836_, _34835_, _34542_);
  nand (_34838_, _34836_, _08702_);
  nor (_34839_, _08702_, _06082_);
  nor (_34840_, _34839_, _08732_);
  nand (_34841_, _34840_, _34838_);
  and (_34842_, _34541_, _08732_);
  nor (_34843_, _34842_, _03515_);
  and (_34844_, _34843_, _34841_);
  nor (_34845_, _06069_, _03516_);
  or (_34846_, _34845_, _34844_);
  nand (_34847_, _34846_, _32165_);
  and (_34849_, _05881_, _03203_);
  nor (_34850_, _34849_, _03628_);
  nand (_34851_, _34850_, _34847_);
  and (_34852_, _09854_, _06749_);
  nor (_34853_, _34587_, _09854_);
  nor (_34854_, _34853_, _34852_);
  and (_34855_, _34854_, _03628_);
  nor (_34856_, _34855_, _11934_);
  nand (_34857_, _34856_, _34851_);
  nor (_34858_, _34541_, _11933_);
  nor (_34860_, _34858_, _03815_);
  and (_34861_, _34860_, _34857_);
  or (_34862_, _34861_, _34538_);
  nand (_34863_, _34862_, _11940_);
  nor (_34864_, _34550_, _11940_);
  nor (_34865_, _34864_, _05103_);
  nand (_34866_, _34865_, _34863_);
  and (_34867_, _05881_, _05103_);
  nor (_34868_, _34867_, _03453_);
  nand (_34869_, _34868_, _34866_);
  and (_34871_, _34854_, _03453_);
  nor (_34872_, _34871_, _11958_);
  nand (_34873_, _34872_, _34869_);
  nor (_34874_, _34541_, _11957_);
  nor (_34875_, _34874_, _03447_);
  and (_34876_, _34875_, _34873_);
  or (_34877_, _34876_, _34537_);
  nand (_34878_, _34877_, _11964_);
  nor (_34879_, _34550_, _11964_);
  nor (_34880_, _34879_, _32154_);
  nand (_34882_, _34880_, _34878_);
  and (_34883_, _32154_, _05881_);
  nor (_34884_, _34883_, _11975_);
  and (_34885_, _34884_, _34882_);
  and (_34886_, _34541_, _11975_);
  or (_34887_, _34886_, _34885_);
  or (_34888_, _34887_, _43004_);
  or (_34889_, _43000_, \oc8051_golden_model_1.PC [7]);
  and (_34890_, _34889_, _41806_);
  and (_43676_, _34890_, _34888_);
  nor (_34892_, _04048_, _11968_);
  nor (_34893_, _04048_, _11944_);
  and (_34894_, _11469_, _03624_);
  nor (_34895_, _11337_, _03192_);
  nor (_34896_, _11595_, _05894_);
  and (_34897_, _11595_, _03585_);
  or (_34898_, _11468_, _10018_);
  nor (_34899_, _11472_, _11466_);
  nor (_34900_, _34899_, _11473_);
  or (_34901_, _34900_, _11685_);
  nand (_34903_, _34901_, _34898_);
  nand (_34904_, _34903_, _09919_);
  and (_34905_, _11468_, _09969_);
  not (_34906_, _34900_);
  nor (_34907_, _34906_, _09969_);
  or (_34908_, _34907_, _34905_);
  nor (_34909_, _34908_, _09921_);
  and (_34910_, _11595_, _03714_);
  nor (_34911_, _03723_, _04768_);
  and (_34912_, _11595_, _03715_);
  or (_34914_, _11468_, _11367_);
  or (_34915_, _34900_, _11369_);
  and (_34916_, _34915_, _34914_);
  or (_34917_, _34916_, _04081_);
  and (_34918_, _11504_, _11595_);
  nor (_34919_, _11599_, _11593_);
  nor (_34920_, _34919_, _11600_);
  and (_34921_, _34920_, _11624_);
  nor (_34922_, _34921_, _34918_);
  nand (_34923_, _34922_, _06073_);
  nand (_34925_, _11596_, _03979_);
  or (_34926_, _04409_, \oc8051_golden_model_1.PC [8]);
  or (_34927_, _34926_, _04729_);
  and (_34928_, _34927_, _34925_);
  or (_34929_, _34928_, _11632_);
  nor (_34930_, _11317_, \oc8051_golden_model_1.PC [8]);
  nor (_34931_, _34930_, _11318_);
  or (_34932_, _34931_, _11642_);
  and (_34933_, _34932_, _34929_);
  nor (_34934_, _34933_, _32191_);
  nor (_34936_, _34931_, _11630_);
  nor (_34937_, _34936_, _34934_);
  nor (_34938_, _34937_, _06073_);
  nor (_34939_, _34938_, _04422_);
  and (_34940_, _34939_, _34923_);
  and (_34941_, _34931_, _04422_);
  or (_34942_, _34941_, _03610_);
  or (_34943_, _34942_, _34940_);
  nand (_34944_, _34943_, _34917_);
  nand (_34945_, _34944_, _11362_);
  nor (_34947_, _34931_, _11362_);
  nor (_34948_, _34947_, _03715_);
  and (_34949_, _34948_, _34945_);
  or (_34950_, _34949_, _34912_);
  nand (_34951_, _34950_, _34911_);
  and (_34952_, _11595_, _03723_);
  nor (_34953_, _34952_, _11660_);
  nand (_34954_, _34953_, _34951_);
  nor (_34955_, _34931_, _11659_);
  nor (_34956_, _34955_, _03729_);
  nand (_34958_, _34956_, _34954_);
  and (_34959_, _11595_, _03729_);
  nor (_34960_, _34959_, _11668_);
  nand (_34961_, _34960_, _34958_);
  nor (_34962_, _34931_, _11666_);
  nor (_34963_, _34962_, _03714_);
  and (_34964_, _34963_, _34961_);
  or (_34965_, _34964_, _34910_);
  nand (_34966_, _34965_, _11671_);
  and (_34967_, _11595_, _03508_);
  nor (_34969_, _34967_, _09917_);
  and (_34970_, _34969_, _34966_);
  or (_34971_, _34970_, _34909_);
  nand (_34972_, _34971_, _09920_);
  nand (_34973_, _34972_, _34904_);
  or (_34974_, _34973_, _03615_);
  nor (_34975_, _34906_, _09876_);
  and (_34976_, _11468_, _09876_);
  nor (_34977_, _34976_, _34975_);
  or (_34978_, _34977_, _04107_);
  and (_34980_, _34978_, _34974_);
  or (_34981_, _34980_, _03604_);
  and (_34982_, _11468_, _10061_);
  and (_34983_, _34900_, _33597_);
  or (_34984_, _34983_, _34982_);
  and (_34985_, _34984_, _03604_);
  nor (_34986_, _34985_, _10025_);
  nand (_34987_, _34986_, _34981_);
  not (_34988_, _34931_);
  and (_34989_, _34988_, _10025_);
  nor (_34991_, _34989_, _03719_);
  nand (_34992_, _34991_, _34987_);
  and (_34993_, _11595_, _03719_);
  nor (_34994_, _34993_, _04766_);
  nand (_34995_, _34994_, _34992_);
  nand (_34996_, _34995_, _32547_);
  nor (_34997_, _32547_, _11596_);
  nor (_34998_, _34997_, _11356_);
  nand (_34999_, _34998_, _34996_);
  nor (_35000_, _34931_, _11355_);
  nor (_35002_, _35000_, _03753_);
  nand (_35003_, _35002_, _34999_);
  and (_35004_, _11595_, _03753_);
  nor (_35005_, _35004_, _11727_);
  nand (_35006_, _35005_, _35003_);
  nand (_35007_, _35006_, _09668_);
  and (_35008_, _11595_, _03752_);
  not (_35009_, _35008_);
  and (_35010_, _35009_, _11350_);
  nand (_35011_, _35010_, _35007_);
  nor (_35013_, _34931_, _11350_);
  nor (_35014_, _35013_, _08187_);
  and (_35015_, _35014_, _35011_);
  nor (_35016_, _11596_, _08186_);
  or (_35017_, _35016_, _07912_);
  nor (_35018_, _35017_, _35015_);
  nor (_35019_, _34931_, _03248_);
  or (_35020_, _35019_, _35018_);
  nand (_35021_, _35020_, _03710_);
  and (_35022_, _11596_, _03505_);
  nor (_35024_, _35022_, _23690_);
  and (_35025_, _35024_, _35021_);
  and (_35026_, _11468_, _03625_);
  nor (_35027_, _35026_, _35025_);
  nand (_35028_, _35027_, _11749_);
  nor (_35029_, _11749_, _11595_);
  nor (_35030_, _35029_, _03222_);
  nand (_35031_, _35030_, _35028_);
  and (_35032_, _11468_, _03222_);
  nor (_35033_, _35032_, _11758_);
  nand (_35035_, _35033_, _35031_);
  nor (_35036_, _34931_, _11756_);
  nor (_35037_, _35036_, _03585_);
  and (_35038_, _35037_, _35035_);
  or (_35039_, _35038_, _34897_);
  nor (_35040_, _11764_, _03169_);
  nand (_35041_, _35040_, _35039_);
  and (_35042_, _34920_, _11764_);
  nor (_35043_, _35042_, _06168_);
  and (_35044_, _35043_, _35041_);
  or (_35046_, _35044_, _34896_);
  nand (_35047_, _35046_, _05886_);
  and (_35048_, _11469_, _03601_);
  nor (_35049_, _35048_, _08363_);
  nand (_35050_, _35049_, _35047_);
  and (_35051_, _11595_, _08363_);
  nor (_35052_, _35051_, _11347_);
  nand (_35053_, _35052_, _35050_);
  nor (_35054_, _11803_, \oc8051_golden_model_1.DPH [0]);
  nor (_35055_, _35054_, _11804_);
  nor (_35057_, _35055_, _11348_);
  nor (_35058_, _35057_, _03584_);
  nand (_35059_, _35058_, _35053_);
  and (_35060_, _11595_, _03584_);
  nor (_35061_, _35060_, _03178_);
  nand (_35062_, _35061_, _35059_);
  nand (_35063_, _35062_, _11820_);
  and (_35064_, _11595_, _08786_);
  and (_35065_, _34920_, _11826_);
  or (_35066_, _35065_, _35064_);
  and (_35068_, _35066_, _11819_);
  nor (_35069_, _35068_, _11824_);
  nand (_35070_, _35069_, _35063_);
  nor (_35071_, _34931_, _11345_);
  nor (_35072_, _35071_, _11342_);
  nand (_35073_, _35072_, _35070_);
  nor (_35074_, _11596_, _11341_);
  nor (_35075_, _35074_, _03600_);
  nand (_35076_, _35075_, _35073_);
  and (_35077_, _11469_, _03600_);
  nor (_35079_, _35077_, _03780_);
  nand (_35080_, _35079_, _35076_);
  and (_35081_, _11595_, _03780_);
  nor (_35082_, _35081_, _03182_);
  nand (_35083_, _35082_, _35080_);
  nand (_35084_, _35083_, _11842_);
  or (_35085_, _34920_, _11826_);
  or (_35086_, _11595_, _08786_);
  and (_35087_, _35086_, _11841_);
  and (_35088_, _35087_, _35085_);
  nor (_35090_, _35088_, _11853_);
  nand (_35091_, _35090_, _35084_);
  nor (_35092_, _34931_, _11851_);
  nor (_35093_, _35092_, _08431_);
  and (_35094_, _35093_, _35091_);
  nor (_35095_, _11596_, _08430_);
  or (_35096_, _35095_, _03622_);
  or (_35097_, _35096_, _35094_);
  and (_35098_, _11469_, _03622_);
  nor (_35099_, _35098_, _03790_);
  and (_35101_, _35099_, _35097_);
  and (_35102_, _11595_, _03790_);
  or (_35103_, _35102_, _35101_);
  nand (_35104_, _35103_, _34895_);
  and (_35105_, _11595_, \oc8051_golden_model_1.PSW [7]);
  and (_35106_, _34920_, _07871_);
  or (_35107_, _35106_, _35105_);
  and (_35108_, _35107_, _11337_);
  nor (_35109_, _35108_, _11864_);
  nand (_35110_, _35109_, _35104_);
  nor (_35112_, _34931_, _11335_);
  nor (_35113_, _35112_, _08460_);
  nand (_35114_, _35113_, _35110_);
  nor (_35115_, _11596_, _08459_);
  nor (_35116_, _35115_, _03624_);
  and (_35117_, _35116_, _35114_);
  or (_35118_, _35117_, _34894_);
  nand (_35119_, _35118_, _07793_);
  nor (_35120_, _11880_, _03201_);
  and (_35121_, _11596_, _03785_);
  not (_35123_, _35121_);
  and (_35124_, _35123_, _35120_);
  nand (_35125_, _35124_, _35119_);
  nor (_35126_, _34920_, _07871_);
  nor (_35127_, _11595_, \oc8051_golden_model_1.PSW [7]);
  nor (_35128_, _35127_, _11881_);
  not (_35129_, _35128_);
  nor (_35130_, _35129_, _35126_);
  nor (_35131_, _35130_, _11885_);
  nand (_35132_, _35131_, _35125_);
  nor (_35134_, _34931_, _11330_);
  nor (_35135_, _35134_, _08508_);
  and (_35136_, _35135_, _35132_);
  nor (_35137_, _11596_, _08507_);
  or (_35138_, _35137_, _08587_);
  or (_35139_, _35138_, _35136_);
  and (_35140_, _34988_, _08587_);
  nor (_35141_, _35140_, _03798_);
  nand (_35142_, _35141_, _35139_);
  and (_35143_, _04620_, _03798_);
  nor (_35145_, _35143_, _03188_);
  nand (_35146_, _35145_, _35142_);
  nand (_35147_, _35146_, _11903_);
  and (_35148_, _34906_, _09854_);
  nor (_35149_, _11468_, _09854_);
  or (_35150_, _35149_, _11903_);
  or (_35151_, _35150_, _35148_);
  and (_35152_, _35151_, _11328_);
  nand (_35153_, _35152_, _35147_);
  nor (_35154_, _34931_, _11328_);
  nor (_35156_, _35154_, _08703_);
  and (_35157_, _35156_, _35153_);
  nor (_35158_, _11596_, _08702_);
  or (_35159_, _35158_, _08732_);
  or (_35160_, _35159_, _35157_);
  and (_35161_, _34988_, _08732_);
  nor (_35162_, _35161_, _03515_);
  nand (_35163_, _35162_, _35160_);
  and (_35164_, _04620_, _03515_);
  nor (_35165_, _35164_, _03203_);
  nand (_35167_, _35165_, _35163_);
  nand (_35168_, _35167_, _03816_);
  and (_35169_, _11469_, _09854_);
  nor (_35170_, _34900_, _09854_);
  nor (_35171_, _35170_, _35169_);
  and (_35172_, _35171_, _03628_);
  nor (_35173_, _35172_, _11934_);
  nand (_35174_, _35173_, _35168_);
  nor (_35175_, _34931_, _11933_);
  nor (_35176_, _35175_, _03815_);
  nand (_35178_, _35176_, _35174_);
  and (_35179_, _11595_, _03815_);
  nor (_35180_, _35179_, _32765_);
  nand (_35181_, _35180_, _35178_);
  nor (_35182_, _34931_, _11940_);
  nor (_35183_, _35182_, _03629_);
  and (_35184_, _35183_, _35181_);
  or (_35185_, _35184_, _34893_);
  nor (_35186_, _03198_, _03453_);
  nand (_35187_, _35186_, _35185_);
  and (_35189_, _35171_, _03453_);
  nor (_35190_, _35189_, _11958_);
  nand (_35191_, _35190_, _35187_);
  nor (_35192_, _34931_, _11957_);
  nor (_35193_, _35192_, _03447_);
  nand (_35194_, _35193_, _35191_);
  and (_35195_, _11595_, _03447_);
  nor (_35196_, _35195_, _33825_);
  nand (_35197_, _35196_, _35194_);
  nor (_35198_, _34931_, _11964_);
  nor (_35200_, _35198_, _03631_);
  and (_35201_, _35200_, _35197_);
  or (_35202_, _35201_, _34892_);
  and (_35203_, _35202_, _24553_);
  and (_35204_, _34931_, _11975_);
  or (_35205_, _35204_, _35203_);
  or (_35206_, _35205_, _43004_);
  or (_35207_, _43000_, \oc8051_golden_model_1.PC [8]);
  and (_35208_, _35207_, _41806_);
  and (_43677_, _35208_, _35206_);
  nor (_35210_, _03414_, _11968_);
  nor (_35211_, _03414_, _11944_);
  nor (_35212_, _11318_, \oc8051_golden_model_1.PC [9]);
  nor (_35213_, _35212_, _11319_);
  nor (_35214_, _35213_, _11328_);
  nor (_35215_, _35213_, _11330_);
  and (_35216_, _11408_, _03624_);
  nor (_35217_, _35213_, _11335_);
  and (_35218_, _11408_, _03622_);
  nor (_35219_, _35213_, _11851_);
  and (_35221_, _11408_, _03600_);
  nor (_35222_, _35213_, _11345_);
  and (_35223_, _11542_, _03585_);
  nor (_35224_, _35213_, _11350_);
  not (_35225_, _35213_);
  and (_35226_, _35225_, _10025_);
  and (_35227_, _11408_, _09876_);
  nor (_35228_, _11473_, _11470_);
  and (_35229_, _35228_, _11412_);
  nor (_35230_, _35228_, _11412_);
  nor (_35232_, _35230_, _35229_);
  nor (_35233_, _35232_, _09876_);
  nor (_35234_, _35233_, _35227_);
  or (_35235_, _35234_, _04107_);
  and (_35236_, _35213_, _04422_);
  and (_35237_, _11504_, _11542_);
  nor (_35238_, _11600_, _11597_);
  and (_35239_, _35238_, _11546_);
  nor (_35240_, _35238_, _11546_);
  nor (_35241_, _35240_, _35239_);
  nor (_35243_, _35241_, _11504_);
  or (_35244_, _35243_, _35237_);
  nor (_35245_, _35244_, _06072_);
  nand (_35246_, _35213_, _04064_);
  and (_35247_, _11630_, _33169_);
  or (_35248_, _35247_, _35213_);
  and (_35249_, _11543_, _03979_);
  nor (_35250_, _35249_, _11632_);
  or (_35251_, _04409_, \oc8051_golden_model_1.PC [9]);
  or (_35252_, _35251_, _04729_);
  nand (_35254_, _35252_, _35250_);
  nand (_35255_, _35254_, _32190_);
  and (_35256_, _35255_, _35248_);
  nor (_35257_, _35256_, _06073_);
  and (_35258_, _35257_, _35246_);
  or (_35259_, _35258_, _04422_);
  nor (_35260_, _35259_, _35245_);
  or (_35261_, _35260_, _35236_);
  and (_35262_, _35261_, _04081_);
  not (_35263_, _35262_);
  not (_35265_, _11362_);
  and (_35266_, _11408_, _11369_);
  not (_35267_, _35232_);
  and (_35268_, _35267_, _11367_);
  nor (_35269_, _35268_, _35266_);
  nor (_35270_, _35269_, _04081_);
  nor (_35271_, _35270_, _35265_);
  and (_35272_, _35271_, _35263_);
  nor (_35273_, _35213_, _11362_);
  nor (_35274_, _35273_, _03715_);
  not (_35276_, _35274_);
  nor (_35277_, _35276_, _35272_);
  and (_35278_, _11542_, _03715_);
  or (_35279_, _35278_, _04768_);
  nor (_35280_, _35279_, _35277_);
  nor (_35281_, _35280_, _03723_);
  and (_35282_, _11542_, _03723_);
  nor (_35283_, _35282_, _11660_);
  not (_35284_, _35283_);
  nor (_35285_, _35284_, _35281_);
  nor (_35287_, _35213_, _11659_);
  nor (_35288_, _35287_, _03729_);
  not (_35289_, _35288_);
  or (_35290_, _35289_, _35285_);
  and (_35291_, _11542_, _03729_);
  nor (_35292_, _35291_, _11668_);
  nand (_35293_, _35292_, _35290_);
  nor (_35294_, _35213_, _11666_);
  nor (_35295_, _35294_, _03714_);
  nand (_35296_, _35295_, _35293_);
  and (_35298_, _11542_, _03714_);
  nor (_35299_, _35298_, _11670_);
  nand (_35300_, _35299_, _35296_);
  nand (_35301_, _35300_, _03510_);
  and (_35302_, _11542_, _03508_);
  nor (_35303_, _35302_, _09917_);
  and (_35304_, _35303_, _35301_);
  and (_35305_, _11408_, _09969_);
  nor (_35306_, _35232_, _09969_);
  or (_35307_, _35306_, _35305_);
  nor (_35309_, _35307_, _09921_);
  or (_35310_, _35309_, _35304_);
  nand (_35311_, _35310_, _09920_);
  and (_35312_, _35267_, _10018_);
  and (_35313_, _11408_, _11685_);
  or (_35314_, _35313_, _09920_);
  or (_35315_, _35314_, _35312_);
  nand (_35316_, _35315_, _35311_);
  or (_35317_, _35316_, _03615_);
  and (_35318_, _35317_, _35235_);
  or (_35320_, _35318_, _03604_);
  and (_35321_, _11408_, _10061_);
  nor (_35322_, _35232_, _10061_);
  or (_35323_, _35322_, _35321_);
  and (_35324_, _35323_, _03604_);
  nor (_35325_, _35324_, _10025_);
  and (_35326_, _35325_, _35320_);
  or (_35327_, _35326_, _35226_);
  nand (_35328_, _35327_, _06840_);
  and (_35329_, _11543_, _03719_);
  not (_35331_, _35329_);
  not (_35332_, _11715_);
  and (_35333_, _23519_, _35332_);
  and (_35334_, _35333_, _35331_);
  and (_35335_, _35334_, _11712_);
  and (_35336_, _35335_, _11710_);
  nand (_35337_, _35336_, _35328_);
  nor (_35338_, _32547_, _11543_);
  nor (_35339_, _35338_, _11356_);
  nand (_35340_, _35339_, _35337_);
  nor (_35342_, _35213_, _11355_);
  nor (_35343_, _35342_, _03753_);
  and (_35344_, _35343_, _35340_);
  and (_35345_, _11542_, _03753_);
  or (_35346_, _35345_, _35344_);
  nand (_35347_, _35346_, _11728_);
  and (_35348_, _11542_, _03752_);
  not (_35349_, _35348_);
  and (_35350_, _35349_, _11350_);
  and (_35351_, _35350_, _35347_);
  or (_35353_, _35351_, _35224_);
  nand (_35354_, _35353_, _08186_);
  nor (_35355_, _11542_, _08186_);
  nor (_35356_, _35355_, _07912_);
  nand (_35357_, _35356_, _35354_);
  nor (_35358_, _35225_, _03248_);
  nor (_35359_, _35358_, _03505_);
  nand (_35360_, _35359_, _35357_);
  and (_35361_, _11543_, _03505_);
  nor (_35362_, _35361_, _23690_);
  nand (_35364_, _35362_, _35360_);
  and (_35365_, _11408_, _03625_);
  nor (_35366_, _35365_, _33299_);
  nand (_35367_, _35366_, _35364_);
  nor (_35368_, _11749_, _11542_);
  nor (_35369_, _35368_, _03222_);
  nand (_35370_, _35369_, _35367_);
  and (_35371_, _11408_, _03222_);
  nor (_35372_, _35371_, _11758_);
  nand (_35373_, _35372_, _35370_);
  nor (_35375_, _35213_, _11756_);
  nor (_35376_, _35375_, _03585_);
  and (_35377_, _35376_, _35373_);
  or (_35378_, _35377_, _35223_);
  nand (_35379_, _35378_, _35040_);
  nor (_35380_, _35241_, _11765_);
  nor (_35381_, _35380_, _06168_);
  nand (_35382_, _35381_, _35379_);
  nor (_35383_, _11542_, _05894_);
  nor (_35384_, _35383_, _03601_);
  nand (_35386_, _35384_, _35382_);
  and (_35387_, _11408_, _03601_);
  nor (_35388_, _35387_, _08363_);
  nand (_35389_, _35388_, _35386_);
  and (_35390_, _11543_, _08363_);
  nor (_35391_, _35390_, _11347_);
  and (_35392_, _35391_, _35389_);
  nor (_35393_, _11804_, \oc8051_golden_model_1.DPH [1]);
  not (_35394_, _35393_);
  nor (_35395_, _11805_, _11348_);
  and (_35397_, _35395_, _35394_);
  or (_35398_, _35397_, _35392_);
  nand (_35399_, _35398_, _10263_);
  and (_35400_, _11542_, _03584_);
  nor (_35401_, _35400_, _03178_);
  nand (_35402_, _35401_, _35399_);
  nand (_35403_, _35402_, _11820_);
  and (_35404_, _11542_, _08786_);
  nor (_35405_, _35241_, _08786_);
  or (_35406_, _35405_, _35404_);
  and (_35408_, _35406_, _11819_);
  nor (_35409_, _35408_, _11824_);
  and (_35410_, _35409_, _35403_);
  or (_35411_, _35410_, _35222_);
  nand (_35412_, _35411_, _11341_);
  nor (_35413_, _11542_, _11341_);
  nor (_35414_, _35413_, _03600_);
  and (_35415_, _35414_, _35412_);
  or (_35416_, _35415_, _35221_);
  nand (_35417_, _35416_, _07778_);
  and (_35419_, _11542_, _03780_);
  nor (_35420_, _35419_, _03182_);
  nand (_35421_, _35420_, _35417_);
  nand (_35422_, _35421_, _11842_);
  nand (_35423_, _35241_, _08786_);
  or (_35424_, _11542_, _08786_);
  and (_35425_, _35424_, _11841_);
  and (_35426_, _35425_, _35423_);
  nor (_35427_, _35426_, _11853_);
  and (_35428_, _35427_, _35422_);
  or (_35430_, _35428_, _35219_);
  nand (_35431_, _35430_, _08430_);
  nor (_35432_, _11542_, _08430_);
  nor (_35433_, _35432_, _03622_);
  and (_35434_, _35433_, _35431_);
  or (_35435_, _35434_, _35218_);
  nand (_35436_, _35435_, _06828_);
  and (_35437_, _11542_, _03790_);
  nor (_35438_, _35437_, _03192_);
  nand (_35439_, _35438_, _35436_);
  nand (_35441_, _35439_, _11338_);
  and (_35442_, _11542_, \oc8051_golden_model_1.PSW [7]);
  nor (_35443_, _35241_, \oc8051_golden_model_1.PSW [7]);
  or (_35444_, _35443_, _35442_);
  and (_35445_, _35444_, _11337_);
  nor (_35446_, _35445_, _11864_);
  and (_35447_, _35446_, _35441_);
  or (_35448_, _35447_, _35217_);
  nand (_35449_, _35448_, _08459_);
  nor (_35450_, _11542_, _08459_);
  nor (_35452_, _35450_, _03624_);
  and (_35453_, _35452_, _35449_);
  or (_35454_, _35453_, _35216_);
  nand (_35455_, _35454_, _07793_);
  and (_35456_, _11542_, _03785_);
  nor (_35457_, _35456_, _03201_);
  nand (_35458_, _35457_, _35455_);
  nand (_35459_, _35458_, _11881_);
  and (_35460_, _35241_, \oc8051_golden_model_1.PSW [7]);
  nor (_35461_, _11542_, \oc8051_golden_model_1.PSW [7]);
  nor (_35463_, _35461_, _11881_);
  not (_35464_, _35463_);
  nor (_35465_, _35464_, _35460_);
  nor (_35466_, _35465_, _11885_);
  and (_35467_, _35466_, _35459_);
  or (_35468_, _35467_, _35215_);
  nand (_35469_, _35468_, _08507_);
  nor (_35470_, _11542_, _08507_);
  nor (_35471_, _35470_, _08587_);
  nand (_35472_, _35471_, _35469_);
  and (_35474_, _35213_, _08587_);
  nor (_35475_, _35474_, _03798_);
  nand (_35476_, _35475_, _35472_);
  nor (_35477_, _03621_, _03188_);
  not (_35478_, _35477_);
  and (_35479_, _04406_, _03798_);
  nor (_35480_, _35479_, _35478_);
  nand (_35481_, _35480_, _35476_);
  and (_35482_, _35267_, _09854_);
  nor (_35483_, _11409_, _09854_);
  nor (_35485_, _35483_, _35482_);
  nor (_35486_, _35485_, _11903_);
  nor (_35487_, _35486_, _11907_);
  and (_35488_, _35487_, _35481_);
  or (_35489_, _35488_, _35214_);
  nand (_35490_, _35489_, _08702_);
  nor (_35491_, _11542_, _08702_);
  nor (_35492_, _35491_, _08732_);
  nand (_35493_, _35492_, _35490_);
  and (_35494_, _35213_, _08732_);
  nor (_35497_, _35494_, _03515_);
  nand (_35498_, _35497_, _35493_);
  not (_35499_, _23212_);
  and (_35500_, _04406_, _03515_);
  nor (_35501_, _35500_, _35499_);
  nand (_35502_, _35501_, _35498_);
  nor (_35503_, _35267_, _09854_);
  and (_35504_, _11409_, _09854_);
  nor (_35505_, _35504_, _35503_);
  and (_35506_, _35505_, _03628_);
  nor (_35508_, _35506_, _11934_);
  nand (_35509_, _35508_, _35502_);
  nor (_35510_, _35213_, _11933_);
  nor (_35511_, _35510_, _03815_);
  nand (_35512_, _35511_, _35509_);
  and (_35513_, _11542_, _03815_);
  nor (_35514_, _35513_, _32765_);
  nand (_35515_, _35514_, _35512_);
  nor (_35516_, _35213_, _11940_);
  nor (_35517_, _35516_, _03629_);
  and (_35520_, _35517_, _35515_);
  or (_35521_, _35520_, _35211_);
  nand (_35522_, _35521_, _35186_);
  and (_35523_, _35505_, _03453_);
  nor (_35524_, _35523_, _11958_);
  nand (_35525_, _35524_, _35522_);
  nor (_35526_, _35213_, _11957_);
  nor (_35527_, _35526_, _03447_);
  nand (_35528_, _35527_, _35525_);
  and (_35529_, _11542_, _03447_);
  nor (_35531_, _35529_, _33825_);
  nand (_35532_, _35531_, _35528_);
  nor (_35533_, _35213_, _11964_);
  nor (_35534_, _35533_, _03631_);
  and (_35535_, _35534_, _35532_);
  or (_35536_, _35535_, _35210_);
  and (_35537_, _35536_, _24553_);
  and (_35538_, _35213_, _11975_);
  or (_35539_, _35538_, _35537_);
  or (_35540_, _35539_, _43004_);
  or (_35543_, _43000_, \oc8051_golden_model_1.PC [9]);
  and (_35544_, _35543_, _41806_);
  and (_43678_, _35544_, _35540_);
  nor (_35545_, _11319_, \oc8051_golden_model_1.PC [10]);
  nor (_35546_, _35545_, _11320_);
  and (_35547_, _35546_, _11975_);
  or (_35548_, _35546_, _11957_);
  not (_35549_, _35546_);
  nand (_35550_, _35549_, _08732_);
  nand (_35551_, _35549_, _08587_);
  nand (_35553_, _11395_, _03624_);
  nand (_35554_, _11395_, _03622_);
  nor (_35555_, _35549_, _11756_);
  or (_35556_, _11529_, _08186_);
  nor (_35557_, _35549_, _11666_);
  or (_35558_, _35546_, _11659_);
  nor (_35559_, _35549_, _11653_);
  nor (_35560_, _11477_, _11474_);
  not (_35561_, _35560_);
  and (_35562_, _35561_, _11405_);
  nor (_35565_, _35561_, _11405_);
  nor (_35566_, _35565_, _35562_);
  or (_35567_, _35566_, _11369_);
  or (_35568_, _11394_, _11367_);
  and (_35569_, _35568_, _03610_);
  and (_35570_, _35569_, _35567_);
  nor (_35571_, _11604_, _11601_);
  not (_35572_, _35571_);
  and (_35573_, _35572_, _11539_);
  nor (_35574_, _35572_, _11539_);
  nor (_35576_, _35574_, _35573_);
  and (_35577_, _35576_, _11624_);
  and (_35578_, _11504_, _11529_);
  or (_35579_, _35578_, _06072_);
  or (_35580_, _35579_, _35577_);
  or (_35581_, _35546_, _11643_);
  not (_35582_, _03979_);
  or (_35583_, _11529_, _35582_);
  or (_35584_, _04409_, \oc8051_golden_model_1.PC [10]);
  or (_35585_, _35584_, _04729_);
  and (_35587_, _35585_, _35583_);
  nand (_35588_, _11630_, _32815_);
  or (_35589_, _35588_, _35587_);
  and (_35590_, _35589_, _35581_);
  or (_35591_, _06073_, _03980_);
  or (_35592_, _35591_, _35590_);
  and (_35593_, _35592_, _11647_);
  and (_35594_, _35593_, _35580_);
  or (_35595_, _35594_, _35570_);
  and (_35596_, _35595_, _11362_);
  or (_35598_, _35596_, _35559_);
  and (_35599_, _35598_, _03730_);
  and (_35600_, _11529_, _14265_);
  nor (_35601_, _35600_, _04768_);
  nand (_35602_, _35601_, _11659_);
  or (_35603_, _35602_, _35599_);
  and (_35604_, _35603_, _35558_);
  or (_35605_, _35604_, _03729_);
  or (_35606_, _11529_, _03737_);
  and (_35607_, _35606_, _11666_);
  and (_35609_, _35607_, _35605_);
  or (_35610_, _35609_, _35557_);
  and (_35611_, _35610_, _03736_);
  and (_35612_, _11529_, _03714_);
  or (_35613_, _35612_, _11670_);
  or (_35614_, _35613_, _35611_);
  and (_35615_, _35614_, _03510_);
  and (_35616_, _11529_, _03508_);
  or (_35617_, _35616_, _09917_);
  or (_35618_, _35617_, _35615_);
  or (_35620_, _35566_, _09969_);
  nand (_35621_, _11395_, _09969_);
  and (_35622_, _35621_, _35620_);
  or (_35623_, _35622_, _09921_);
  and (_35624_, _35623_, _35618_);
  or (_35625_, _35624_, _32519_);
  and (_35626_, _11394_, _11685_);
  and (_35627_, _35566_, _10018_);
  or (_35628_, _35627_, _35626_);
  or (_35629_, _35628_, _09920_);
  and (_35631_, _35629_, _35625_);
  or (_35632_, _35631_, _03615_);
  and (_35633_, _11394_, _09876_);
  and (_35634_, _35566_, _11693_);
  or (_35635_, _35634_, _04107_);
  or (_35636_, _35635_, _35633_);
  and (_35637_, _35636_, _09856_);
  and (_35638_, _35637_, _35632_);
  or (_35639_, _35566_, _10061_);
  nand (_35640_, _11395_, _10061_);
  and (_35642_, _35640_, _03604_);
  and (_35643_, _35642_, _35639_);
  or (_35644_, _35643_, _10025_);
  or (_35645_, _35644_, _35638_);
  nand (_35646_, _35549_, _10025_);
  and (_35647_, _32547_, _06840_);
  and (_35648_, _35647_, _35646_);
  and (_35649_, _35648_, _35645_);
  not (_35650_, _11529_);
  nor (_35651_, _35647_, _35650_);
  nand (_35653_, _11355_, _03227_);
  or (_35654_, _35653_, _35651_);
  or (_35655_, _35654_, _35649_);
  or (_35656_, _35546_, _11355_);
  and (_35657_, _35656_, _09669_);
  and (_35658_, _35657_, _35655_);
  nand (_35659_, _11529_, _03753_);
  nand (_35660_, _35659_, _11728_);
  or (_35661_, _35660_, _35658_);
  nand (_35662_, _35650_, _03752_);
  and (_35664_, _35662_, _11350_);
  and (_35665_, _35664_, _35661_);
  nor (_35666_, _35549_, _11350_);
  or (_35667_, _35666_, _08187_);
  or (_35668_, _35667_, _35665_);
  and (_35669_, _35668_, _35556_);
  or (_35670_, _35669_, _07912_);
  or (_35671_, _35546_, _03248_);
  and (_35672_, _35671_, _03710_);
  and (_35673_, _35672_, _35670_);
  nand (_35675_, _11529_, _03505_);
  nand (_35676_, _35675_, _23689_);
  or (_35677_, _35676_, _35673_);
  nand (_35678_, _11395_, _03625_);
  and (_35679_, _35678_, _11749_);
  and (_35680_, _35679_, _35677_);
  nor (_35681_, _11749_, _35650_);
  or (_35682_, _35681_, _03222_);
  or (_35683_, _35682_, _35680_);
  nand (_35684_, _11395_, _03222_);
  and (_35686_, _35684_, _11756_);
  and (_35687_, _35686_, _35683_);
  nor (_35688_, _35687_, _35555_);
  nor (_35689_, _35688_, _03585_);
  nand (_35690_, _11529_, _03585_);
  nand (_35691_, _35690_, _35040_);
  or (_35692_, _35691_, _35689_);
  or (_35693_, _35576_, _11765_);
  and (_35694_, _35693_, _05894_);
  and (_35695_, _35694_, _35692_);
  nor (_35697_, _35650_, _05894_);
  or (_35698_, _35697_, _03601_);
  or (_35699_, _35698_, _35695_);
  nand (_35700_, _11395_, _03601_);
  and (_35701_, _35700_, _08364_);
  and (_35702_, _35701_, _35699_);
  and (_35703_, _11529_, _08363_);
  or (_35704_, _35703_, _11347_);
  or (_35705_, _35704_, _35702_);
  nor (_35706_, _11805_, \oc8051_golden_model_1.DPH [2]);
  nor (_35708_, _35706_, _11806_);
  or (_35709_, _35708_, _11348_);
  and (_35710_, _35709_, _10263_);
  and (_35711_, _35710_, _35705_);
  and (_35712_, _11529_, _03584_);
  or (_35713_, _35712_, _35711_);
  nor (_35714_, _11819_, _03178_);
  and (_35715_, _35714_, _35713_);
  or (_35716_, _35576_, _08786_);
  or (_35717_, _11529_, _11826_);
  and (_35719_, _35717_, _11819_);
  and (_35720_, _35719_, _35716_);
  or (_35721_, _35720_, _11824_);
  or (_35722_, _35721_, _35715_);
  or (_35723_, _35546_, _11345_);
  and (_35724_, _35723_, _11341_);
  and (_35725_, _35724_, _35722_);
  and (_35726_, _11529_, _11342_);
  or (_35727_, _35726_, _03600_);
  or (_35728_, _35727_, _35725_);
  nand (_35730_, _11395_, _03600_);
  and (_35731_, _35730_, _35728_);
  or (_35732_, _35731_, _03780_);
  nand (_35733_, _35650_, _03780_);
  and (_35734_, _35733_, _23991_);
  and (_35735_, _35734_, _35732_);
  or (_35736_, _35576_, _11826_);
  or (_35737_, _11529_, _08786_);
  and (_35738_, _35737_, _11841_);
  and (_35739_, _35738_, _35736_);
  or (_35741_, _35739_, _11853_);
  or (_35742_, _35741_, _35735_);
  or (_35743_, _35546_, _11851_);
  and (_35744_, _35743_, _08430_);
  and (_35745_, _35744_, _35742_);
  nor (_35746_, _35650_, _08430_);
  or (_35747_, _35746_, _03622_);
  or (_35748_, _35747_, _35745_);
  and (_35749_, _35748_, _35554_);
  or (_35750_, _35749_, _03790_);
  nand (_35752_, _35650_, _03790_);
  and (_35753_, _35752_, _34895_);
  and (_35754_, _35753_, _35750_);
  or (_35755_, _35576_, \oc8051_golden_model_1.PSW [7]);
  or (_35756_, _11529_, _07871_);
  and (_35757_, _35756_, _11337_);
  and (_35758_, _35757_, _35755_);
  or (_35759_, _35758_, _11864_);
  or (_35760_, _35759_, _35754_);
  or (_35761_, _35546_, _11335_);
  and (_35763_, _35761_, _08459_);
  and (_35764_, _35763_, _35760_);
  nor (_35765_, _35650_, _08459_);
  or (_35766_, _35765_, _03624_);
  or (_35767_, _35766_, _35764_);
  and (_35768_, _35767_, _35553_);
  or (_35769_, _35768_, _03785_);
  nand (_35770_, _35650_, _03785_);
  and (_35771_, _35770_, _35120_);
  and (_35772_, _35771_, _35769_);
  or (_35774_, _35576_, _07871_);
  or (_35775_, _11529_, \oc8051_golden_model_1.PSW [7]);
  and (_35776_, _35775_, _11880_);
  and (_35777_, _35776_, _35774_);
  or (_35778_, _35777_, _11885_);
  or (_35779_, _35778_, _35772_);
  or (_35780_, _35546_, _11330_);
  and (_35781_, _35780_, _08507_);
  and (_35782_, _35781_, _35779_);
  nor (_35783_, _35650_, _08507_);
  or (_35785_, _35783_, _08587_);
  or (_35786_, _35785_, _35782_);
  and (_35787_, _35786_, _35551_);
  or (_35788_, _35787_, _03798_);
  nand (_35789_, _04875_, _03798_);
  and (_35790_, _35789_, _35477_);
  and (_35791_, _35790_, _35788_);
  or (_35792_, _35566_, _11908_);
  or (_35793_, _11394_, _09854_);
  and (_35794_, _35793_, _03621_);
  and (_35796_, _35794_, _35792_);
  or (_35797_, _35796_, _11907_);
  or (_35798_, _35797_, _35791_);
  or (_35799_, _35546_, _11328_);
  and (_35800_, _35799_, _08702_);
  and (_35801_, _35800_, _35798_);
  nor (_35802_, _35650_, _08702_);
  or (_35803_, _35802_, _08732_);
  or (_35804_, _35803_, _35801_);
  and (_35805_, _35804_, _35550_);
  or (_35807_, _35805_, _03515_);
  nand (_35808_, _04875_, _03515_);
  and (_35809_, _35808_, _23212_);
  and (_35810_, _35809_, _35807_);
  or (_35811_, _35566_, _09854_);
  nand (_35812_, _11395_, _09854_);
  and (_35813_, _35812_, _35811_);
  and (_35814_, _35813_, _03628_);
  or (_35815_, _35814_, _11934_);
  or (_35816_, _35815_, _35810_);
  or (_35818_, _35546_, _11933_);
  and (_35819_, _35818_, _35816_);
  or (_35820_, _35819_, _03815_);
  nand (_35821_, _35650_, _03815_);
  and (_35822_, _35821_, _11940_);
  and (_35823_, _35822_, _35820_);
  nor (_35824_, _35549_, _11940_);
  or (_35825_, _35824_, _03629_);
  or (_35826_, _35825_, _35823_);
  nand (_35827_, _03904_, _03629_);
  and (_35829_, _35827_, _35186_);
  and (_35830_, _35829_, _35826_);
  and (_35831_, _35813_, _03453_);
  or (_35832_, _35831_, _11958_);
  or (_35833_, _35832_, _35830_);
  and (_35834_, _35833_, _35548_);
  or (_35835_, _35834_, _03447_);
  nand (_35836_, _35650_, _03447_);
  and (_35837_, _35836_, _11964_);
  and (_35838_, _35837_, _35835_);
  nor (_35840_, _35549_, _11964_);
  or (_35841_, _35840_, _03631_);
  or (_35842_, _35841_, _35838_);
  nand (_35843_, _03904_, _03631_);
  and (_35844_, _35843_, _24553_);
  and (_35845_, _35844_, _35842_);
  or (_35846_, _35845_, _35547_);
  or (_35847_, _35846_, _43004_);
  or (_35848_, _43000_, \oc8051_golden_model_1.PC [10]);
  and (_35849_, _35848_, _41806_);
  and (_43679_, _35849_, _35847_);
  nor (_35851_, _11320_, \oc8051_golden_model_1.PC [11]);
  nor (_35852_, _35851_, _11321_);
  nor (_35853_, _35852_, _11328_);
  nor (_35854_, _35852_, _11330_);
  nor (_35855_, _35852_, _11335_);
  nor (_35856_, _35852_, _11851_);
  nor (_35857_, _35852_, _11345_);
  nor (_35858_, _11533_, _05894_);
  and (_35859_, _11399_, _03222_);
  and (_35861_, _11399_, _10061_);
  nor (_35862_, _35562_, _11396_);
  and (_35863_, _35862_, _11403_);
  nor (_35864_, _35862_, _11403_);
  nor (_35865_, _35864_, _35863_);
  nor (_35866_, _35865_, _10061_);
  or (_35867_, _35866_, _35861_);
  and (_35868_, _35867_, _03604_);
  and (_35869_, _11399_, _11685_);
  not (_35870_, _35865_);
  and (_35872_, _35870_, _10018_);
  or (_35873_, _35872_, _35869_);
  nor (_35874_, _35873_, _09920_);
  and (_35875_, _11533_, _03729_);
  nor (_35876_, _11360_, _11533_);
  and (_35877_, _11400_, _11369_);
  and (_35878_, _35865_, _11367_);
  or (_35879_, _35878_, _04081_);
  or (_35880_, _35879_, _35877_);
  and (_35881_, _11504_, _11533_);
  not (_35883_, _35881_);
  nor (_35884_, _35573_, _11530_);
  and (_35885_, _35884_, _11537_);
  nor (_35886_, _35884_, _11537_);
  nor (_35887_, _35886_, _35885_);
  nor (_35888_, _35887_, _11504_);
  nor (_35889_, _35888_, _06072_);
  and (_35890_, _35889_, _35883_);
  nor (_35891_, _35852_, _11643_);
  and (_35892_, _11534_, _03980_);
  and (_35894_, _11534_, _03979_);
  nor (_35895_, _04409_, \oc8051_golden_model_1.PC [11]);
  and (_35896_, _35895_, _11634_);
  nor (_35897_, _35896_, _35894_);
  nor (_35898_, _35897_, _11632_);
  nor (_35899_, _35898_, _35892_);
  nor (_35900_, _35899_, _11631_);
  nor (_35901_, _35900_, _35891_);
  nor (_35902_, _35901_, _06073_);
  or (_35903_, _35902_, _33523_);
  or (_35905_, _35903_, _35890_);
  and (_35906_, _35905_, _35880_);
  or (_35907_, _35906_, _35265_);
  not (_35908_, _35852_);
  or (_35909_, _35908_, _11653_);
  and (_35910_, _35909_, _11360_);
  and (_35911_, _35910_, _35907_);
  nor (_35912_, _35911_, _35876_);
  nor (_35913_, _35912_, _11660_);
  nor (_35914_, _35852_, _11659_);
  nor (_35916_, _35914_, _03729_);
  not (_35917_, _35916_);
  nor (_35918_, _35917_, _35913_);
  nor (_35919_, _35918_, _35875_);
  nor (_35920_, _35919_, _11668_);
  nor (_35921_, _35908_, _11666_);
  nor (_35922_, _35921_, _11673_);
  not (_35923_, _35922_);
  or (_35924_, _35923_, _35920_);
  nor (_35925_, _11672_, _11533_);
  nor (_35927_, _35925_, _09917_);
  and (_35928_, _35927_, _35924_);
  or (_35929_, _35870_, _09969_);
  nand (_35930_, _11400_, _09969_);
  and (_35931_, _35930_, _09917_);
  and (_35932_, _35931_, _35929_);
  or (_35933_, _35932_, _09919_);
  nor (_35934_, _35933_, _35928_);
  or (_35935_, _35934_, _35874_);
  or (_35936_, _35935_, _03615_);
  and (_35938_, _11399_, _09876_);
  nor (_35939_, _35865_, _09876_);
  nor (_35940_, _35939_, _35938_);
  or (_35941_, _35940_, _04107_);
  and (_35942_, _35941_, _35936_);
  nor (_35943_, _35942_, _03604_);
  or (_35944_, _35943_, _35868_);
  nand (_35945_, _35944_, _11358_);
  and (_35946_, _35852_, _10025_);
  not (_35947_, _35946_);
  and (_35949_, _35947_, _11720_);
  nand (_35950_, _35949_, _35945_);
  nor (_35951_, _11720_, _11533_);
  nor (_35952_, _35951_, _11356_);
  nand (_35953_, _35952_, _35950_);
  not (_35954_, _11729_);
  nor (_35955_, _35908_, _11355_);
  nor (_35956_, _35955_, _35954_);
  and (_35957_, _35956_, _35953_);
  or (_35958_, _11729_, _11533_);
  nand (_35960_, _35958_, _11350_);
  or (_35961_, _35960_, _35957_);
  nor (_35962_, _35908_, _11350_);
  nor (_35963_, _35962_, _08187_);
  nand (_35964_, _35963_, _35961_);
  nor (_35965_, _11533_, _08186_);
  nor (_35966_, _35965_, _07912_);
  nand (_35967_, _35966_, _35964_);
  nor (_35968_, _35908_, _03248_);
  nor (_35969_, _35968_, _11741_);
  nand (_35971_, _35969_, _35967_);
  nor (_35972_, _11740_, _11533_);
  nor (_35973_, _35972_, _03625_);
  nand (_35974_, _35973_, _35971_);
  and (_35975_, _11399_, _03625_);
  nor (_35976_, _35975_, _33299_);
  nand (_35977_, _35976_, _35974_);
  nor (_35978_, _11749_, _11533_);
  nor (_35979_, _35978_, _03222_);
  and (_35980_, _35979_, _35977_);
  or (_35982_, _35980_, _35859_);
  nand (_35983_, _35982_, _11756_);
  nor (_35984_, _35908_, _11756_);
  nor (_35985_, _35984_, _11761_);
  nand (_35986_, _35985_, _35983_);
  nor (_35987_, _11760_, _11533_);
  nor (_35988_, _35987_, _11764_);
  nand (_35989_, _35988_, _35986_);
  nor (_35990_, _35887_, _11765_);
  nor (_35991_, _35990_, _06168_);
  and (_35993_, _35991_, _35989_);
  or (_35994_, _35993_, _35858_);
  nand (_35995_, _35994_, _05886_);
  and (_35996_, _11400_, _03601_);
  nor (_35997_, _35996_, _08363_);
  and (_35998_, _35997_, _35995_);
  and (_35999_, _11533_, _08363_);
  or (_36000_, _35999_, _35998_);
  nand (_36001_, _36000_, _11348_);
  nor (_36002_, _11806_, \oc8051_golden_model_1.DPH [3]);
  not (_36004_, _36002_);
  nor (_36005_, _11807_, _11348_);
  and (_36006_, _36005_, _36004_);
  nor (_36007_, _36006_, _11816_);
  nand (_36008_, _36007_, _36001_);
  nor (_36009_, _11815_, _11533_);
  nor (_36010_, _36009_, _11819_);
  nand (_36011_, _36010_, _36008_);
  and (_36012_, _11533_, _08786_);
  nor (_36013_, _35887_, _08786_);
  or (_36015_, _36013_, _36012_);
  and (_36016_, _36015_, _11819_);
  nor (_36017_, _36016_, _11824_);
  and (_36018_, _36017_, _36011_);
  or (_36019_, _36018_, _35857_);
  nand (_36020_, _36019_, _11341_);
  nor (_36021_, _11533_, _11341_);
  nor (_36022_, _36021_, _03600_);
  nand (_36023_, _36022_, _36020_);
  not (_36024_, _11838_);
  and (_36026_, _11399_, _03600_);
  nor (_36027_, _36026_, _36024_);
  nand (_36028_, _36027_, _36023_);
  nor (_36029_, _11838_, _11533_);
  nor (_36030_, _36029_, _11841_);
  nand (_36031_, _36030_, _36028_);
  nand (_36032_, _35887_, _08786_);
  or (_36033_, _11533_, _08786_);
  and (_36034_, _36033_, _11841_);
  and (_36035_, _36034_, _36032_);
  nor (_36037_, _36035_, _11853_);
  and (_36038_, _36037_, _36031_);
  or (_36039_, _36038_, _35856_);
  nand (_36040_, _36039_, _08430_);
  nor (_36041_, _11533_, _08430_);
  nor (_36042_, _36041_, _03622_);
  nand (_36043_, _36042_, _36040_);
  and (_36044_, _11399_, _03622_);
  nor (_36045_, _36044_, _10754_);
  and (_36046_, _36045_, _36043_);
  nor (_36048_, _11534_, _11337_);
  nor (_36049_, _36048_, _24116_);
  or (_36050_, _36049_, _36046_);
  and (_36051_, _11533_, \oc8051_golden_model_1.PSW [7]);
  nor (_36052_, _35887_, \oc8051_golden_model_1.PSW [7]);
  or (_36053_, _36052_, _36051_);
  and (_36054_, _36053_, _11337_);
  nor (_36055_, _36054_, _11864_);
  and (_36056_, _36055_, _36050_);
  or (_36057_, _36056_, _35855_);
  nand (_36059_, _36057_, _08459_);
  nor (_36060_, _11533_, _08459_);
  nor (_36061_, _36060_, _03624_);
  nand (_36062_, _36061_, _36059_);
  not (_36063_, _11877_);
  and (_36064_, _11399_, _03624_);
  nor (_36065_, _36064_, _36063_);
  and (_36066_, _36065_, _36062_);
  nor (_36067_, _11880_, _11534_);
  nor (_36068_, _36067_, _24239_);
  or (_36070_, _36068_, _36066_);
  and (_36071_, _35887_, \oc8051_golden_model_1.PSW [7]);
  nor (_36072_, _11533_, \oc8051_golden_model_1.PSW [7]);
  nor (_36073_, _36072_, _11881_);
  not (_36074_, _36073_);
  nor (_36075_, _36074_, _36071_);
  nor (_36076_, _36075_, _11885_);
  and (_36077_, _36076_, _36070_);
  or (_36078_, _36077_, _35854_);
  nand (_36079_, _36078_, _08507_);
  nor (_36081_, _11533_, _08507_);
  nor (_36082_, _36081_, _08587_);
  and (_36083_, _36082_, _36079_);
  and (_36084_, _35852_, _08587_);
  or (_36085_, _36084_, _03798_);
  nor (_36086_, _36085_, _36083_);
  and (_36087_, _05005_, _03798_);
  or (_36088_, _36087_, _36086_);
  nand (_36089_, _36088_, _06399_);
  and (_36090_, _11534_, _03188_);
  nor (_36092_, _36090_, _03621_);
  nand (_36093_, _36092_, _36089_);
  and (_36094_, _35865_, _09854_);
  nor (_36095_, _11399_, _09854_);
  or (_36096_, _36095_, _11903_);
  nor (_36097_, _36096_, _36094_);
  nor (_36098_, _36097_, _11907_);
  and (_36099_, _36098_, _36093_);
  or (_36100_, _36099_, _35853_);
  nand (_36101_, _36100_, _08702_);
  nor (_36103_, _11533_, _08702_);
  nor (_36104_, _36103_, _08732_);
  and (_36105_, _36104_, _36101_);
  and (_36106_, _35852_, _08732_);
  or (_36107_, _36106_, _03515_);
  nor (_36108_, _36107_, _36105_);
  and (_36109_, _05005_, _03515_);
  or (_36110_, _36109_, _36108_);
  nand (_36111_, _36110_, _32165_);
  and (_36112_, _11534_, _03203_);
  nor (_36114_, _36112_, _03628_);
  nand (_36115_, _36114_, _36111_);
  nor (_36116_, _35870_, _09854_);
  and (_36117_, _11400_, _09854_);
  nor (_36118_, _36117_, _36116_);
  and (_36119_, _36118_, _03628_);
  nor (_36120_, _36119_, _11934_);
  nand (_36121_, _36120_, _36115_);
  nor (_36122_, _35852_, _11933_);
  nor (_36123_, _36122_, _03815_);
  nand (_36125_, _36123_, _36121_);
  and (_36126_, _11533_, _03815_);
  nor (_36127_, _36126_, _32765_);
  nand (_36128_, _36127_, _36125_);
  nor (_36129_, _35852_, _11940_);
  nor (_36130_, _36129_, _03629_);
  nand (_36131_, _36130_, _36128_);
  nor (_36132_, _11944_, _03581_);
  nor (_36133_, _36132_, _03198_);
  nand (_36134_, _36133_, _36131_);
  and (_36136_, _11534_, _03198_);
  nor (_36137_, _36136_, _03453_);
  nand (_36138_, _36137_, _36134_);
  and (_36139_, _36118_, _03453_);
  nor (_36140_, _36139_, _11958_);
  nand (_36141_, _36140_, _36138_);
  nor (_36142_, _35852_, _11957_);
  nor (_36143_, _36142_, _03447_);
  nand (_36144_, _36143_, _36141_);
  and (_36145_, _11533_, _03447_);
  nor (_36147_, _36145_, _33825_);
  nand (_36148_, _36147_, _36144_);
  nor (_36149_, _35852_, _11964_);
  nor (_36150_, _36149_, _03631_);
  nand (_36151_, _36150_, _36148_);
  nor (_36152_, _11968_, _03581_);
  nor (_36153_, _36152_, _03196_);
  and (_36154_, _36153_, _36151_);
  and (_36155_, _11534_, _03196_);
  nor (_36156_, _36155_, _36154_);
  and (_36158_, _36156_, _11976_);
  and (_36159_, _35852_, _11975_);
  or (_36160_, _36159_, _36158_);
  or (_36161_, _36160_, _43004_);
  or (_36162_, _43000_, \oc8051_golden_model_1.PC [11]);
  and (_36163_, _36162_, _41806_);
  and (_43682_, _36163_, _36161_);
  and (_36164_, _11525_, _08786_);
  and (_36165_, _11611_, _11608_);
  nor (_36166_, _36165_, _11612_);
  and (_36168_, _36166_, _11826_);
  or (_36169_, _36168_, _36164_);
  and (_36170_, _36169_, _11819_);
  and (_36171_, _11390_, _03222_);
  and (_36172_, _11390_, _11685_);
  and (_36173_, _11484_, _11481_);
  nor (_36174_, _36173_, _11485_);
  and (_36175_, _36174_, _10018_);
  or (_36176_, _36175_, _36172_);
  nor (_36177_, _36176_, _09920_);
  nor (_36179_, _11321_, \oc8051_golden_model_1.PC [12]);
  nor (_36180_, _36179_, _11322_);
  nor (_36181_, _36180_, _11653_);
  not (_36182_, _36180_);
  nor (_36183_, _36182_, _11643_);
  not (_36184_, _36183_);
  and (_36185_, _11525_, _04409_);
  and (_36186_, _09029_, \oc8051_golden_model_1.PC [12]);
  and (_36187_, _36186_, _33169_);
  nor (_36188_, _36187_, _36185_);
  not (_36190_, _36188_);
  and (_36191_, _36190_, _32816_);
  and (_36192_, _11525_, _03980_);
  nor (_36193_, _36192_, _06073_);
  not (_36194_, _36193_);
  nor (_36195_, _36194_, _36191_);
  and (_36196_, _36195_, _36184_);
  and (_36197_, _11504_, _11525_);
  and (_36198_, _36166_, _11624_);
  or (_36199_, _36198_, _36197_);
  nor (_36201_, _36199_, _06072_);
  nor (_36202_, _36201_, _36196_);
  nor (_36203_, _36202_, _33523_);
  and (_36204_, _11390_, _11369_);
  not (_36205_, _36204_);
  and (_36206_, _36174_, _11367_);
  nor (_36207_, _36206_, _04081_);
  and (_36208_, _36207_, _36205_);
  nor (_36209_, _36208_, _36203_);
  nor (_36210_, _36209_, _35265_);
  nor (_36212_, _36210_, _36181_);
  nor (_36213_, _36212_, _11652_);
  nor (_36214_, _11360_, _11525_);
  nor (_36215_, _36214_, _11660_);
  not (_36216_, _36215_);
  nor (_36217_, _36216_, _36213_);
  nor (_36218_, _36182_, _11659_);
  nor (_36219_, _36218_, _03729_);
  not (_36220_, _36219_);
  nor (_36221_, _36220_, _36217_);
  and (_36223_, _11526_, _03729_);
  nor (_36224_, _36223_, _11668_);
  not (_36225_, _36224_);
  or (_36226_, _36225_, _36221_);
  nor (_36227_, _36182_, _11666_);
  nor (_36228_, _36227_, _11673_);
  and (_36229_, _36228_, _36226_);
  nor (_36230_, _11672_, _11525_);
  or (_36231_, _36230_, _09917_);
  or (_36232_, _36231_, _36229_);
  and (_36234_, _11391_, _09969_);
  nor (_36235_, _36174_, _09969_);
  or (_36236_, _36235_, _09921_);
  or (_36237_, _36236_, _36234_);
  and (_36238_, _36237_, _09920_);
  and (_36239_, _36238_, _36232_);
  or (_36240_, _36239_, _03615_);
  or (_36241_, _36240_, _36177_);
  and (_36242_, _36174_, _11693_);
  and (_36243_, _11390_, _09876_);
  nor (_36245_, _36243_, _36242_);
  nor (_36246_, _36245_, _04107_);
  nor (_36247_, _36246_, _03604_);
  and (_36248_, _36247_, _36241_);
  nor (_36249_, _36174_, _10061_);
  and (_36250_, _11391_, _10061_);
  nor (_36251_, _36250_, _36249_);
  nor (_36252_, _36251_, _09856_);
  nor (_36253_, _36252_, _10025_);
  not (_36254_, _36253_);
  or (_36256_, _36254_, _36248_);
  and (_36257_, _36180_, _10025_);
  not (_36258_, _36257_);
  and (_36259_, _36258_, _11720_);
  nand (_36260_, _36259_, _36256_);
  nor (_36261_, _11720_, _11525_);
  nor (_36262_, _36261_, _11356_);
  nand (_36263_, _36262_, _36260_);
  nor (_36264_, _36182_, _11355_);
  nor (_36265_, _36264_, _35954_);
  nand (_36267_, _36265_, _36263_);
  nor (_36268_, _11729_, _11525_);
  not (_36269_, _36268_);
  and (_36270_, _36269_, _11350_);
  nand (_36271_, _36270_, _36267_);
  nor (_36272_, _36182_, _11350_);
  nor (_36273_, _36272_, _08187_);
  nand (_36274_, _36273_, _36271_);
  nor (_36275_, _11525_, _08186_);
  nor (_36276_, _36275_, _07912_);
  nand (_36278_, _36276_, _36274_);
  nor (_36279_, _36182_, _03248_);
  nor (_36280_, _36279_, _11741_);
  nand (_36281_, _36280_, _36278_);
  nor (_36282_, _11740_, _11525_);
  nor (_36283_, _36282_, _03625_);
  nand (_36284_, _36283_, _36281_);
  and (_36285_, _11390_, _03625_);
  nor (_36286_, _36285_, _33299_);
  nand (_36287_, _36286_, _36284_);
  nor (_36289_, _11749_, _11525_);
  nor (_36290_, _36289_, _03222_);
  and (_36291_, _36290_, _36287_);
  or (_36292_, _36291_, _36171_);
  nand (_36293_, _36292_, _11756_);
  nor (_36294_, _36182_, _11756_);
  nor (_36295_, _36294_, _11761_);
  nand (_36296_, _36295_, _36293_);
  nor (_36297_, _11760_, _11525_);
  nor (_36298_, _36297_, _11764_);
  nand (_36300_, _36298_, _36296_);
  and (_36301_, _36166_, _11764_);
  nor (_36302_, _36301_, _06168_);
  and (_36303_, _36302_, _36300_);
  nor (_36304_, _11526_, _03601_);
  nor (_36305_, _36304_, _05895_);
  or (_36306_, _36305_, _36303_);
  and (_36307_, _11390_, _03601_);
  nor (_36308_, _36307_, _08363_);
  nand (_36309_, _36308_, _36306_);
  and (_36311_, _11526_, _08363_);
  nor (_36312_, _36311_, _11347_);
  nand (_36313_, _36312_, _36309_);
  nor (_36314_, _11807_, \oc8051_golden_model_1.DPH [4]);
  nor (_36315_, _36314_, _11808_);
  and (_36316_, _36315_, _11347_);
  nor (_36317_, _36316_, _11816_);
  nand (_36318_, _36317_, _36313_);
  nor (_36319_, _11815_, _11525_);
  nor (_36320_, _36319_, _11819_);
  and (_36322_, _36320_, _36318_);
  or (_36323_, _36322_, _36170_);
  nand (_36324_, _36323_, _11345_);
  nor (_36325_, _36182_, _11345_);
  nor (_36326_, _36325_, _11342_);
  nand (_36327_, _36326_, _36324_);
  nor (_36328_, _11525_, _11341_);
  nor (_36329_, _36328_, _03600_);
  nand (_36330_, _36329_, _36327_);
  and (_36331_, _11390_, _03600_);
  nor (_36333_, _36331_, _36024_);
  nand (_36334_, _36333_, _36330_);
  nor (_36335_, _11838_, _11525_);
  nor (_36336_, _36335_, _11841_);
  nand (_36337_, _36336_, _36334_);
  nand (_36338_, _11525_, _11826_);
  nand (_36339_, _36166_, _08786_);
  and (_36340_, _36339_, _36338_);
  or (_36341_, _36340_, _11842_);
  nand (_36342_, _36341_, _36337_);
  nand (_36344_, _36342_, _11851_);
  nor (_36345_, _36182_, _11851_);
  nor (_36346_, _36345_, _08431_);
  nand (_36347_, _36346_, _36344_);
  nor (_36348_, _11525_, _08430_);
  nor (_36349_, _36348_, _03622_);
  nand (_36350_, _36349_, _36347_);
  and (_36351_, _11390_, _03622_);
  nor (_36352_, _36351_, _10754_);
  and (_36353_, _36352_, _36350_);
  nor (_36355_, _11526_, _11337_);
  nor (_36356_, _36355_, _24116_);
  nor (_36357_, _36356_, _36353_);
  and (_36358_, _11525_, \oc8051_golden_model_1.PSW [7]);
  and (_36359_, _36166_, _07871_);
  or (_36360_, _36359_, _36358_);
  and (_36361_, _36360_, _11337_);
  or (_36362_, _36361_, _36357_);
  nand (_36363_, _36362_, _11335_);
  nor (_36364_, _36182_, _11335_);
  nor (_36366_, _36364_, _08460_);
  nand (_36367_, _36366_, _36363_);
  nor (_36368_, _11525_, _08459_);
  nor (_36369_, _36368_, _03624_);
  nand (_36370_, _36369_, _36367_);
  and (_36371_, _11390_, _03624_);
  nor (_36372_, _36371_, _36063_);
  and (_36373_, _36372_, _36370_);
  nor (_36374_, _11880_, _11526_);
  nor (_36375_, _36374_, _24239_);
  or (_36377_, _36375_, _36373_);
  nand (_36378_, _11525_, _07871_);
  nand (_36379_, _36166_, \oc8051_golden_model_1.PSW [7]);
  and (_36380_, _36379_, _36378_);
  or (_36381_, _36380_, _11881_);
  nand (_36382_, _36381_, _36377_);
  nand (_36383_, _36382_, _11330_);
  nor (_36384_, _36182_, _11330_);
  nor (_36385_, _36384_, _08508_);
  nand (_36386_, _36385_, _36383_);
  nor (_36388_, _11525_, _08507_);
  nor (_36389_, _36388_, _08587_);
  and (_36390_, _36389_, _36386_);
  and (_36391_, _36180_, _08587_);
  or (_36392_, _36391_, _03798_);
  nor (_36393_, _36392_, _36390_);
  and (_36394_, _05777_, _03798_);
  or (_36395_, _36394_, _36393_);
  nand (_36396_, _36395_, _06399_);
  and (_36397_, _11526_, _03188_);
  nor (_36399_, _36397_, _03621_);
  and (_36400_, _36399_, _36396_);
  and (_36401_, _36174_, _09854_);
  nor (_36402_, _11391_, _09854_);
  nor (_36403_, _36402_, _36401_);
  nor (_36404_, _36403_, _11903_);
  or (_36405_, _36404_, _36400_);
  nand (_36406_, _36405_, _11328_);
  nor (_36407_, _36182_, _11328_);
  nor (_36408_, _36407_, _08703_);
  nand (_36410_, _36408_, _36406_);
  nor (_36411_, _11525_, _08702_);
  nor (_36412_, _36411_, _08732_);
  nand (_36413_, _36412_, _36410_);
  and (_36414_, _36180_, _08732_);
  nor (_36415_, _36414_, _03515_);
  nand (_36416_, _36415_, _36413_);
  and (_36417_, _05777_, _03515_);
  nor (_36418_, _36417_, _03203_);
  and (_36419_, _36418_, _36416_);
  and (_36421_, _11525_, _03203_);
  or (_36422_, _36421_, _03628_);
  or (_36423_, _36422_, _36419_);
  nor (_36424_, _36174_, _09854_);
  and (_36425_, _11391_, _09854_);
  nor (_36426_, _36425_, _36424_);
  nor (_36427_, _36426_, _03816_);
  nor (_36428_, _36427_, _11934_);
  nand (_36429_, _36428_, _36423_);
  nor (_36430_, _36182_, _11933_);
  nor (_36432_, _36430_, _03815_);
  nand (_36433_, _36432_, _36429_);
  and (_36434_, _11526_, _03815_);
  nor (_36435_, _36434_, _32765_);
  nand (_36436_, _36435_, _36433_);
  nor (_36437_, _36182_, _11940_);
  nor (_36438_, _36437_, _03629_);
  nand (_36439_, _36438_, _36436_);
  and (_36440_, _03486_, _03629_);
  nor (_36441_, _36440_, _03198_);
  and (_36443_, _36441_, _36439_);
  and (_36444_, _11525_, _03198_);
  or (_36445_, _36444_, _03453_);
  or (_36446_, _36445_, _36443_);
  nor (_36447_, _36426_, _03823_);
  nor (_36448_, _36447_, _11958_);
  nand (_36449_, _36448_, _36446_);
  nor (_36450_, _36182_, _11957_);
  nor (_36451_, _36450_, _03447_);
  nand (_36452_, _36451_, _36449_);
  and (_36454_, _11526_, _03447_);
  nor (_36455_, _36454_, _33825_);
  nand (_36456_, _36455_, _36452_);
  nor (_36457_, _36182_, _11964_);
  nor (_36458_, _36457_, _03631_);
  nand (_36459_, _36458_, _36456_);
  and (_36460_, _03486_, _03631_);
  nor (_36461_, _36460_, _03196_);
  nand (_36462_, _36461_, _36459_);
  and (_36463_, _11525_, _03196_);
  nor (_36465_, _36463_, _11975_);
  and (_36466_, _36465_, _36462_);
  and (_36467_, _36182_, _11975_);
  nor (_36468_, _36467_, _36466_);
  or (_36469_, _36468_, _43004_);
  or (_36470_, _43000_, \oc8051_golden_model_1.PC [12]);
  and (_36471_, _36470_, _41806_);
  and (_43683_, _36471_, _36469_);
  nor (_36472_, _11322_, \oc8051_golden_model_1.PC [13]);
  nor (_36473_, _36472_, _11323_);
  or (_36475_, _36473_, _11328_);
  or (_36476_, _36473_, _11330_);
  or (_36477_, _36473_, _11335_);
  or (_36478_, _11523_, _11522_);
  not (_36479_, _36478_);
  nor (_36480_, _36479_, _11613_);
  and (_36481_, _36479_, _11613_);
  or (_36482_, _36481_, _36480_);
  or (_36483_, _36482_, _08786_);
  or (_36484_, _11521_, _11826_);
  and (_36486_, _36484_, _11819_);
  and (_36487_, _36486_, _36483_);
  or (_36488_, _11521_, _05894_);
  and (_36489_, _11385_, _03222_);
  or (_36490_, _36473_, _11350_);
  and (_36491_, _36473_, _11356_);
  or (_36492_, _11388_, _11387_);
  not (_36493_, _36492_);
  nor (_36494_, _36493_, _11486_);
  and (_36495_, _36493_, _11486_);
  or (_36497_, _36495_, _36494_);
  or (_36498_, _36497_, _10061_);
  nand (_36499_, _11386_, _10061_);
  and (_36500_, _36499_, _03604_);
  and (_36501_, _36500_, _36498_);
  and (_36502_, _36497_, _10018_);
  and (_36503_, _11385_, _11685_);
  or (_36504_, _36503_, _36502_);
  or (_36505_, _36504_, _09920_);
  and (_36506_, _11521_, _03729_);
  or (_36508_, _11360_, _11521_);
  or (_36509_, _36497_, _11369_);
  or (_36510_, _11385_, _11367_);
  and (_36511_, _36510_, _03610_);
  and (_36512_, _36511_, _36509_);
  and (_36513_, _36482_, _11624_);
  and (_36514_, _11504_, _11521_);
  or (_36515_, _36514_, _06072_);
  or (_36516_, _36515_, _36513_);
  or (_36517_, _36473_, _11643_);
  or (_36519_, _11521_, _04763_);
  or (_36520_, _11521_, _35582_);
  or (_36521_, _04409_, \oc8051_golden_model_1.PC [13]);
  or (_36522_, _36521_, _04729_);
  nand (_36523_, _36522_, _36520_);
  nand (_36524_, _36523_, _32816_);
  and (_36525_, _36524_, _36519_);
  and (_36526_, _36525_, _36517_);
  or (_36527_, _36526_, _06073_);
  and (_36528_, _36527_, _11647_);
  and (_36530_, _36528_, _36516_);
  or (_36531_, _36530_, _36512_);
  and (_36532_, _36531_, _11362_);
  and (_36533_, _36473_, _11654_);
  or (_36534_, _36533_, _11652_);
  or (_36535_, _36534_, _36532_);
  and (_36536_, _36535_, _36508_);
  or (_36537_, _36536_, _11660_);
  or (_36538_, _36473_, _11659_);
  and (_36539_, _36538_, _03737_);
  and (_36541_, _36539_, _36537_);
  or (_36542_, _36541_, _36506_);
  and (_36543_, _36542_, _11666_);
  and (_36544_, _36473_, _11668_);
  or (_36545_, _36544_, _11673_);
  or (_36546_, _36545_, _36543_);
  or (_36547_, _11672_, _11521_);
  and (_36548_, _36547_, _09921_);
  and (_36549_, _36548_, _36546_);
  or (_36550_, _36497_, _09969_);
  nand (_36552_, _11386_, _09969_);
  and (_36553_, _36552_, _09917_);
  and (_36554_, _36553_, _36550_);
  or (_36555_, _36554_, _09919_);
  or (_36556_, _36555_, _36549_);
  and (_36557_, _36556_, _36505_);
  or (_36558_, _36557_, _03615_);
  and (_36559_, _36497_, _11693_);
  and (_36560_, _11385_, _09876_);
  or (_36561_, _36560_, _04107_);
  or (_36563_, _36561_, _36559_);
  and (_36564_, _36563_, _09856_);
  and (_36565_, _36564_, _36558_);
  or (_36566_, _36565_, _36501_);
  and (_36567_, _36566_, _11358_);
  nand (_36568_, _36473_, _10025_);
  nand (_36569_, _36568_, _11720_);
  or (_36570_, _36569_, _36567_);
  or (_36571_, _11720_, _11521_);
  and (_36572_, _36571_, _11355_);
  and (_36574_, _36572_, _36570_);
  or (_36575_, _36574_, _36491_);
  and (_36576_, _36575_, _11729_);
  nand (_36577_, _35954_, _11521_);
  nand (_36578_, _36577_, _11350_);
  or (_36579_, _36578_, _36576_);
  and (_36580_, _36579_, _36490_);
  or (_36581_, _36580_, _08187_);
  or (_36582_, _11521_, _08186_);
  and (_36583_, _36582_, _03248_);
  and (_36585_, _36583_, _36581_);
  nand (_36586_, _36473_, _07912_);
  nand (_36587_, _36586_, _11740_);
  or (_36588_, _36587_, _36585_);
  or (_36589_, _11740_, _11521_);
  and (_36590_, _36589_, _08832_);
  and (_36591_, _36590_, _36588_);
  nand (_36592_, _11385_, _03625_);
  nand (_36593_, _36592_, _11749_);
  or (_36594_, _36593_, _36591_);
  or (_36596_, _11749_, _11521_);
  and (_36597_, _36596_, _03589_);
  and (_36598_, _36597_, _36594_);
  or (_36599_, _36598_, _36489_);
  and (_36600_, _36599_, _11756_);
  and (_36601_, _36473_, _11758_);
  or (_36602_, _36601_, _11761_);
  or (_36603_, _36602_, _36600_);
  or (_36604_, _11760_, _11521_);
  and (_36605_, _36604_, _11765_);
  and (_36607_, _36605_, _36603_);
  and (_36608_, _36482_, _11764_);
  or (_36609_, _36608_, _06168_);
  or (_36610_, _36609_, _36607_);
  and (_36611_, _36610_, _36488_);
  or (_36612_, _36611_, _03601_);
  or (_36613_, _11385_, _05886_);
  and (_36614_, _36613_, _08364_);
  and (_36615_, _36614_, _36612_);
  and (_36616_, _11521_, _08363_);
  or (_36618_, _36616_, _36615_);
  and (_36619_, _36618_, _11348_);
  or (_36620_, _11808_, \oc8051_golden_model_1.DPH [5]);
  nor (_36621_, _11809_, _11348_);
  and (_36622_, _36621_, _36620_);
  or (_36623_, _36622_, _11816_);
  or (_36624_, _36623_, _36619_);
  or (_36625_, _11815_, _11521_);
  and (_36626_, _36625_, _11820_);
  and (_36627_, _36626_, _36624_);
  or (_36629_, _36627_, _36487_);
  and (_36630_, _36629_, _11345_);
  and (_36631_, _36473_, _11824_);
  or (_36632_, _36631_, _11342_);
  or (_36633_, _36632_, _36630_);
  or (_36634_, _11521_, _11341_);
  and (_36635_, _36634_, _07766_);
  and (_36636_, _36635_, _36633_);
  nand (_36637_, _11385_, _03600_);
  nand (_36638_, _36637_, _11838_);
  or (_36640_, _36638_, _36636_);
  or (_36641_, _11838_, _11521_);
  and (_36642_, _36641_, _11842_);
  and (_36643_, _36642_, _36640_);
  or (_36644_, _36482_, _11826_);
  or (_36645_, _11521_, _08786_);
  and (_36646_, _36645_, _11841_);
  and (_36647_, _36646_, _36644_);
  or (_36648_, _36647_, _36643_);
  and (_36649_, _36648_, _11851_);
  and (_36651_, _36473_, _11853_);
  or (_36652_, _36651_, _08431_);
  or (_36653_, _36652_, _36649_);
  or (_36654_, _11521_, _08430_);
  and (_36655_, _36654_, _07777_);
  and (_36656_, _36655_, _36653_);
  nand (_36657_, _11385_, _03622_);
  nand (_36658_, _36657_, _10753_);
  or (_36659_, _36658_, _36656_);
  and (_36660_, _11521_, _11338_);
  or (_36662_, _36660_, _24116_);
  and (_36663_, _36662_, _36659_);
  or (_36664_, _36482_, \oc8051_golden_model_1.PSW [7]);
  or (_36665_, _11521_, _07871_);
  and (_36666_, _36665_, _11337_);
  and (_36667_, _36666_, _36664_);
  or (_36668_, _36667_, _11864_);
  or (_36669_, _36668_, _36663_);
  and (_36670_, _36669_, _36477_);
  or (_36671_, _36670_, _08460_);
  or (_36673_, _11521_, _08459_);
  and (_36674_, _36673_, _07795_);
  and (_36675_, _36674_, _36671_);
  nand (_36676_, _11385_, _03624_);
  nand (_36677_, _36676_, _11877_);
  or (_36678_, _36677_, _36675_);
  and (_36679_, _11881_, _11521_);
  or (_36680_, _36679_, _24239_);
  and (_36681_, _36680_, _36678_);
  or (_36682_, _36482_, _07871_);
  or (_36684_, _11521_, \oc8051_golden_model_1.PSW [7]);
  and (_36685_, _36684_, _11880_);
  and (_36686_, _36685_, _36682_);
  or (_36687_, _36686_, _11885_);
  or (_36688_, _36687_, _36681_);
  and (_36689_, _36688_, _36476_);
  or (_36690_, _36689_, _08508_);
  or (_36691_, _11521_, _08507_);
  and (_36692_, _36691_, _08588_);
  and (_36693_, _36692_, _36690_);
  and (_36695_, _36473_, _08587_);
  or (_36696_, _36695_, _03798_);
  or (_36697_, _36696_, _36693_);
  nand (_36698_, _05469_, _03798_);
  and (_36699_, _36698_, _36697_);
  or (_36700_, _36699_, _03188_);
  or (_36701_, _11521_, _06399_);
  and (_36702_, _36701_, _11903_);
  and (_36703_, _36702_, _36700_);
  or (_36704_, _36497_, _11908_);
  or (_36706_, _11385_, _09854_);
  and (_36707_, _36706_, _03621_);
  and (_36708_, _36707_, _36704_);
  or (_36709_, _36708_, _11907_);
  or (_36710_, _36709_, _36703_);
  and (_36711_, _36710_, _36475_);
  or (_36712_, _36711_, _08703_);
  or (_36713_, _11521_, _08702_);
  and (_36714_, _36713_, _08733_);
  and (_36715_, _36714_, _36712_);
  and (_36717_, _36473_, _08732_);
  or (_36718_, _36717_, _03515_);
  or (_36719_, _36718_, _36715_);
  nand (_36720_, _05469_, _03515_);
  and (_36721_, _36720_, _36719_);
  or (_36722_, _36721_, _03203_);
  or (_36723_, _11521_, _32165_);
  and (_36724_, _36723_, _03816_);
  and (_36725_, _36724_, _36722_);
  nand (_36726_, _11386_, _09854_);
  or (_36728_, _36497_, _09854_);
  and (_36729_, _36728_, _36726_);
  and (_36730_, _36729_, _03628_);
  or (_36731_, _36730_, _11934_);
  or (_36732_, _36731_, _36725_);
  or (_36733_, _36473_, _11933_);
  and (_36734_, _36733_, _04246_);
  and (_36735_, _36734_, _36732_);
  nand (_36736_, _11521_, _03815_);
  nand (_36737_, _36736_, _11940_);
  or (_36739_, _36737_, _36735_);
  or (_36740_, _36473_, _11940_);
  and (_36741_, _36740_, _11944_);
  and (_36742_, _36741_, _36739_);
  nor (_36743_, _03860_, _11944_);
  or (_36744_, _36743_, _03198_);
  or (_36745_, _36744_, _36742_);
  or (_36746_, _11521_, _12371_);
  and (_36747_, _36746_, _03823_);
  and (_36748_, _36747_, _36745_);
  and (_36750_, _36729_, _03453_);
  or (_36751_, _36750_, _11958_);
  or (_36752_, _36751_, _36748_);
  or (_36753_, _36473_, _11957_);
  and (_36754_, _36753_, _03514_);
  and (_36755_, _36754_, _36752_);
  nand (_36756_, _11521_, _03447_);
  nand (_36757_, _36756_, _11964_);
  or (_36758_, _36757_, _36755_);
  or (_36759_, _36473_, _11964_);
  and (_36761_, _36759_, _11968_);
  and (_36762_, _36761_, _36758_);
  nor (_36763_, _03860_, _11968_);
  or (_36764_, _36763_, _03196_);
  or (_36765_, _36764_, _36762_);
  not (_36766_, _11521_);
  nand (_36767_, _36766_, _03196_);
  and (_36768_, _36767_, _11976_);
  and (_36769_, _36768_, _36765_);
  and (_36770_, _36473_, _11975_);
  or (_36772_, _36770_, _36769_);
  or (_36773_, _36772_, _43004_);
  or (_36774_, _43000_, \oc8051_golden_model_1.PC [13]);
  and (_36775_, _36774_, _41806_);
  and (_43684_, _36775_, _36773_);
  nor (_36776_, _11323_, \oc8051_golden_model_1.PC [14]);
  nor (_36777_, _36776_, _11324_);
  nor (_36778_, _36777_, _08733_);
  nor (_36779_, _11877_, _11515_);
  nor (_36780_, _11515_, _10753_);
  nor (_36782_, _11838_, _11515_);
  nor (_36783_, _11815_, _11515_);
  and (_36784_, _11488_, _11383_);
  nor (_36785_, _36784_, _11489_);
  or (_36786_, _36785_, _11685_);
  or (_36787_, _11378_, _10018_);
  and (_36788_, _36787_, _09919_);
  and (_36789_, _36788_, _36786_);
  and (_36790_, _36777_, _11668_);
  nor (_36791_, _36777_, _11659_);
  or (_36793_, _36785_, _11369_);
  or (_36794_, _11378_, _11367_);
  and (_36795_, _36794_, _36793_);
  nor (_36796_, _36795_, _04081_);
  and (_36797_, _11615_, _11519_);
  nor (_36798_, _36797_, _11616_);
  nand (_36799_, _36798_, _11624_);
  or (_36800_, _11624_, _11515_);
  and (_36801_, _36800_, _06073_);
  nand (_36802_, _36801_, _36799_);
  nor (_36804_, _36777_, _11642_);
  nor (_36805_, _11632_, \oc8051_golden_model_1.PC [14]);
  and (_36806_, _36805_, _09029_);
  and (_36807_, _36806_, _33169_);
  nor (_36808_, _36807_, _36804_);
  nor (_36809_, _36808_, _03980_);
  not (_36810_, _36809_);
  nor (_36811_, _03980_, _04409_);
  nor (_36812_, _36811_, _11514_);
  nor (_36813_, _36812_, _11631_);
  and (_36815_, _36813_, _36810_);
  not (_36816_, _36777_);
  nor (_36817_, _36816_, _11630_);
  nor (_36818_, _36817_, _06073_);
  not (_36819_, _36818_);
  nor (_36820_, _36819_, _36815_);
  nor (_36821_, _36820_, _04422_);
  nand (_36822_, _36821_, _36802_);
  and (_36823_, _36777_, _04422_);
  nor (_36824_, _36823_, _03610_);
  and (_36826_, _36824_, _36822_);
  or (_36827_, _36826_, _36796_);
  nand (_36828_, _36827_, _11362_);
  nor (_36829_, _36777_, _11362_);
  nor (_36830_, _36829_, _11652_);
  nand (_36831_, _36830_, _36828_);
  nor (_36832_, _11360_, _11515_);
  nor (_36833_, _36832_, _11660_);
  and (_36834_, _36833_, _36831_);
  or (_36835_, _36834_, _36791_);
  nand (_36837_, _36835_, _03737_);
  nor (_36838_, _11514_, _03737_);
  nor (_36839_, _36838_, _11668_);
  and (_36840_, _36839_, _36837_);
  or (_36841_, _36840_, _36790_);
  nand (_36842_, _36841_, _11672_);
  nor (_36843_, _11672_, _11515_);
  nor (_36844_, _36843_, _09917_);
  nand (_36845_, _36844_, _36842_);
  and (_36846_, _11378_, _09969_);
  not (_36848_, _36785_);
  nor (_36849_, _36848_, _09969_);
  or (_36850_, _36849_, _36846_);
  nor (_36851_, _36850_, _09921_);
  nor (_36852_, _36851_, _09919_);
  and (_36853_, _36852_, _36845_);
  or (_36854_, _36853_, _03615_);
  or (_36855_, _36854_, _36789_);
  and (_36856_, _11378_, _09876_);
  nor (_36857_, _36848_, _09876_);
  or (_36859_, _36857_, _04107_);
  or (_36860_, _36859_, _36856_);
  and (_36861_, _36860_, _09856_);
  nand (_36862_, _36861_, _36855_);
  and (_36863_, _11379_, _10061_);
  nor (_36864_, _36785_, _10061_);
  or (_36865_, _36864_, _09856_);
  or (_36866_, _36865_, _36863_);
  and (_36867_, _36866_, _11358_);
  and (_36868_, _36867_, _36862_);
  nor (_36870_, _36777_, _11358_);
  or (_36871_, _36870_, _36868_);
  and (_36872_, _36871_, _11720_);
  nor (_36873_, _11720_, _11514_);
  or (_36874_, _36873_, _36872_);
  nand (_36875_, _36874_, _11355_);
  nor (_36876_, _36777_, _11355_);
  nor (_36877_, _36876_, _35954_);
  and (_36878_, _36877_, _36875_);
  nor (_36879_, _11729_, _11515_);
  nor (_36881_, _36879_, _36878_);
  nand (_36882_, _36881_, _11350_);
  nor (_36883_, _36777_, _11350_);
  nor (_36884_, _36883_, _08187_);
  nand (_36885_, _36884_, _36882_);
  nor (_36886_, _11515_, _08186_);
  nor (_36887_, _36886_, _07912_);
  nand (_36888_, _36887_, _36885_);
  nor (_36889_, _36777_, _03248_);
  nor (_36890_, _36889_, _11741_);
  nand (_36892_, _36890_, _36888_);
  nor (_36893_, _11740_, _11515_);
  nor (_36894_, _36893_, _03625_);
  nand (_36895_, _36894_, _36892_);
  nor (_36896_, _11378_, _08832_);
  nor (_36897_, _36896_, _33299_);
  nand (_36898_, _36897_, _36895_);
  nor (_36899_, _11749_, _11515_);
  nor (_36900_, _36899_, _03222_);
  nand (_36901_, _36900_, _36898_);
  nor (_36903_, _11378_, _03589_);
  nor (_36904_, _36903_, _11758_);
  nand (_36905_, _36904_, _36901_);
  and (_36906_, _36777_, _11758_);
  nor (_36907_, _36906_, _11761_);
  nand (_36908_, _36907_, _36905_);
  nor (_36909_, _11760_, _11514_);
  nor (_36910_, _36909_, _11764_);
  and (_36911_, _36910_, _36908_);
  and (_36912_, _36798_, _11764_);
  nor (_36914_, _36912_, _36911_);
  or (_36915_, _36914_, _06168_);
  or (_36916_, _11515_, _05894_);
  and (_36917_, _36916_, _05886_);
  nand (_36918_, _36917_, _36915_);
  nor (_36919_, _11378_, _05886_);
  nor (_36920_, _36919_, _08363_);
  nand (_36921_, _36920_, _36918_);
  and (_36922_, _11514_, _08363_);
  nor (_36923_, _36922_, _11347_);
  nand (_36925_, _36923_, _36921_);
  nor (_36926_, _11809_, \oc8051_golden_model_1.DPH [6]);
  nor (_36927_, _36926_, _11810_);
  nor (_36928_, _36927_, _11348_);
  nor (_36929_, _36928_, _11816_);
  and (_36930_, _36929_, _36925_);
  or (_36931_, _36930_, _36783_);
  nand (_36932_, _36931_, _11820_);
  and (_36933_, _11514_, _08786_);
  and (_36934_, _36798_, _11826_);
  or (_36936_, _36934_, _36933_);
  and (_36937_, _36936_, _11819_);
  nor (_36938_, _36937_, _11824_);
  nand (_36939_, _36938_, _36932_);
  nor (_36940_, _36777_, _11345_);
  nor (_36941_, _36940_, _11342_);
  nand (_36942_, _36941_, _36939_);
  nor (_36943_, _11515_, _11341_);
  nor (_36944_, _36943_, _03600_);
  nand (_36945_, _36944_, _36942_);
  nor (_36947_, _11378_, _07766_);
  nor (_36948_, _36947_, _36024_);
  and (_36949_, _36948_, _36945_);
  or (_36950_, _36949_, _36782_);
  nand (_36951_, _36950_, _11842_);
  or (_36952_, _36798_, _11826_);
  or (_36953_, _11514_, _08786_);
  and (_36954_, _36953_, _11841_);
  and (_36955_, _36954_, _36952_);
  nor (_36956_, _36955_, _11853_);
  nand (_36958_, _36956_, _36951_);
  nor (_36959_, _36777_, _11851_);
  nor (_36960_, _36959_, _08431_);
  nand (_36961_, _36960_, _36958_);
  nor (_36962_, _11515_, _08430_);
  nor (_36963_, _36962_, _03622_);
  nand (_36964_, _36963_, _36961_);
  nor (_36965_, _11378_, _07777_);
  nor (_36966_, _36965_, _10754_);
  and (_36967_, _36966_, _36964_);
  or (_36969_, _36967_, _36780_);
  nand (_36970_, _36969_, _11338_);
  and (_36971_, _11514_, \oc8051_golden_model_1.PSW [7]);
  and (_36972_, _36798_, _07871_);
  or (_36973_, _36972_, _36971_);
  and (_36974_, _36973_, _11337_);
  nor (_36975_, _36974_, _11864_);
  nand (_36976_, _36975_, _36970_);
  nor (_36977_, _36777_, _11335_);
  nor (_36978_, _36977_, _08460_);
  nand (_36980_, _36978_, _36976_);
  nor (_36981_, _11515_, _08459_);
  nor (_36982_, _36981_, _03624_);
  nand (_36983_, _36982_, _36980_);
  nor (_36984_, _11378_, _07795_);
  nor (_36985_, _36984_, _36063_);
  and (_36986_, _36985_, _36983_);
  or (_36987_, _36986_, _36779_);
  nand (_36988_, _36987_, _11881_);
  nor (_36989_, _36798_, _07871_);
  nor (_36991_, _11514_, \oc8051_golden_model_1.PSW [7]);
  nor (_36992_, _36991_, _11881_);
  not (_36993_, _36992_);
  nor (_36994_, _36993_, _36989_);
  nor (_36995_, _36994_, _11885_);
  nand (_36996_, _36995_, _36988_);
  nor (_36997_, _36777_, _11330_);
  nor (_36998_, _36997_, _08508_);
  nand (_36999_, _36998_, _36996_);
  nor (_37000_, _11515_, _08507_);
  nor (_37002_, _37000_, _08587_);
  nand (_37003_, _37002_, _36999_);
  nor (_37004_, _36777_, _08588_);
  nor (_37005_, _37004_, _03798_);
  and (_37006_, _37005_, _37003_);
  nor (_37007_, _05363_, _10652_);
  or (_37008_, _37007_, _03188_);
  or (_37009_, _37008_, _37006_);
  nor (_37010_, _11514_, _06399_);
  nor (_37011_, _37010_, _03621_);
  nand (_37013_, _37011_, _37009_);
  nor (_37014_, _11378_, _09854_);
  and (_37015_, _36848_, _09854_);
  or (_37016_, _37015_, _11903_);
  or (_37017_, _37016_, _37014_);
  and (_37018_, _37017_, _11328_);
  nand (_37019_, _37018_, _37013_);
  nor (_37020_, _36777_, _11328_);
  nor (_37021_, _37020_, _08703_);
  nand (_37022_, _37021_, _37019_);
  nor (_37024_, _11515_, _08702_);
  nor (_37025_, _37024_, _08732_);
  and (_37026_, _37025_, _37022_);
  or (_37027_, _37026_, _36778_);
  nand (_37028_, _37027_, _03516_);
  and (_37029_, _05363_, _03515_);
  nor (_37030_, _37029_, _03203_);
  and (_37031_, _37030_, _37028_);
  and (_37032_, _11514_, _03203_);
  or (_37033_, _37032_, _03628_);
  nor (_37035_, _37033_, _37031_);
  and (_37036_, _11379_, _09854_);
  nor (_37037_, _36785_, _09854_);
  nor (_37038_, _37037_, _37036_);
  nor (_37039_, _37038_, _03816_);
  or (_37040_, _37039_, _37035_);
  and (_37041_, _37040_, _11933_);
  nor (_37042_, _36777_, _11933_);
  or (_37043_, _37042_, _37041_);
  nand (_37044_, _37043_, _04246_);
  nor (_37046_, _11514_, _04246_);
  nor (_37047_, _37046_, _32765_);
  nand (_37048_, _37047_, _37044_);
  nor (_37049_, _36816_, _11940_);
  nor (_37050_, _37049_, _03629_);
  nand (_37051_, _37050_, _37048_);
  and (_37052_, _03629_, _03549_);
  nor (_37053_, _37052_, _03198_);
  nand (_37054_, _37053_, _37051_);
  and (_37055_, _11514_, _03198_);
  nor (_37057_, _37055_, _03453_);
  nand (_37058_, _37057_, _37054_);
  nor (_37059_, _37038_, _03823_);
  nor (_37060_, _37059_, _11958_);
  nand (_37061_, _37060_, _37058_);
  nor (_37062_, _36816_, _11957_);
  nor (_37063_, _37062_, _03447_);
  nand (_37064_, _37063_, _37061_);
  nor (_37065_, _11514_, _03514_);
  nor (_37066_, _37065_, _33825_);
  nand (_37068_, _37066_, _37064_);
  nor (_37069_, _36816_, _11964_);
  nor (_37070_, _37069_, _03631_);
  nand (_37071_, _37070_, _37068_);
  and (_37072_, _03631_, _03549_);
  nor (_37073_, _37072_, _03196_);
  nand (_37074_, _37073_, _37071_);
  and (_37075_, _11514_, _03196_);
  nor (_37076_, _37075_, _11975_);
  and (_37077_, _37076_, _37074_);
  nor (_37079_, _36777_, _11976_);
  nor (_37080_, _37079_, _37077_);
  or (_37081_, _37080_, _43004_);
  or (_37082_, _43000_, \oc8051_golden_model_1.PC [14]);
  and (_37083_, _37082_, _41806_);
  and (_43685_, _37083_, _37081_);
  and (_37084_, _43004_, \oc8051_golden_model_1.P0INREG [0]);
  or (_37085_, _37084_, _01169_);
  and (_43686_, _37085_, _41806_);
  and (_37086_, _43004_, \oc8051_golden_model_1.P0INREG [1]);
  or (_37088_, _37086_, _01153_);
  and (_43687_, _37088_, _41806_);
  and (_37089_, _43004_, \oc8051_golden_model_1.P0INREG [2]);
  or (_37090_, _37089_, _01186_);
  and (_43688_, _37090_, _41806_);
  and (_37091_, _43004_, \oc8051_golden_model_1.P0INREG [3]);
  or (_37092_, _37091_, _01202_);
  and (_43689_, _37092_, _41806_);
  and (_37093_, _43004_, \oc8051_golden_model_1.P0INREG [4]);
  or (_37094_, _37093_, _01162_);
  and (_43690_, _37094_, _41806_);
  and (_37096_, _43004_, \oc8051_golden_model_1.P0INREG [5]);
  or (_37097_, _37096_, _01146_);
  and (_43691_, _37097_, _41806_);
  and (_37098_, _43004_, \oc8051_golden_model_1.P0INREG [6]);
  or (_37099_, _37098_, _01179_);
  and (_43692_, _37099_, _41806_);
  and (_37100_, _43004_, \oc8051_golden_model_1.P1INREG [0]);
  or (_37101_, _37100_, _01133_);
  and (_43695_, _37101_, _41806_);
  and (_37103_, _43004_, \oc8051_golden_model_1.P1INREG [1]);
  or (_37104_, _37103_, _01083_);
  and (_43696_, _37104_, _41806_);
  and (_37105_, _43004_, \oc8051_golden_model_1.P1INREG [2]);
  or (_37106_, _37105_, _01117_);
  and (_43697_, _37106_, _41806_);
  and (_37107_, _43004_, \oc8051_golden_model_1.P1INREG [3]);
  or (_37108_, _37107_, _01099_);
  and (_43698_, _37108_, _41806_);
  and (_37109_, _43004_, \oc8051_golden_model_1.P1INREG [4]);
  or (_37111_, _37109_, _01126_);
  and (_43699_, _37111_, _41806_);
  and (_37112_, _43004_, \oc8051_golden_model_1.P1INREG [5]);
  or (_37113_, _37112_, _01076_);
  and (_43702_, _37113_, _41806_);
  and (_37114_, _43004_, \oc8051_golden_model_1.P1INREG [6]);
  or (_37115_, _37114_, _01110_);
  and (_43703_, _37115_, _41806_);
  and (_37116_, _43004_, \oc8051_golden_model_1.P2INREG [0]);
  or (_37117_, _37116_, _00899_);
  and (_43704_, _37117_, _41806_);
  and (_37119_, _43004_, \oc8051_golden_model_1.P2INREG [1]);
  or (_37120_, _37119_, _00926_);
  and (_43705_, _37120_, _41806_);
  and (_37121_, _43004_, \oc8051_golden_model_1.P2INREG [2]);
  or (_37122_, _37121_, _00874_);
  and (_43706_, _37122_, _41806_);
  and (_37123_, _43004_, \oc8051_golden_model_1.P2INREG [3]);
  or (_37124_, _37123_, _00916_);
  and (_43707_, _37124_, _41806_);
  and (_37126_, _43004_, \oc8051_golden_model_1.P2INREG [4]);
  or (_37127_, _37126_, _00891_);
  and (_43708_, _37127_, _41806_);
  and (_37128_, _43004_, \oc8051_golden_model_1.P2INREG [5]);
  or (_37129_, _37128_, _00933_);
  and (_43709_, _37129_, _41806_);
  and (_37130_, _43004_, \oc8051_golden_model_1.P2INREG [6]);
  or (_37131_, _37130_, _00881_);
  and (_43710_, _37131_, _41806_);
  and (_37132_, _43004_, \oc8051_golden_model_1.P3INREG [0]);
  or (_37134_, _37132_, _01019_);
  and (_43713_, _37134_, _41806_);
  and (_37135_, _43004_, \oc8051_golden_model_1.P3INREG [1]);
  or (_37136_, _37135_, _01045_);
  and (_43714_, _37136_, _41806_);
  and (_37137_, _43004_, \oc8051_golden_model_1.P3INREG [2]);
  or (_37138_, _37137_, _00996_);
  and (_43715_, _37138_, _41806_);
  and (_37139_, _43004_, \oc8051_golden_model_1.P3INREG [3]);
  or (_37140_, _37139_, _01035_);
  and (_43716_, _37140_, _41806_);
  and (_37142_, _43004_, \oc8051_golden_model_1.P3INREG [4]);
  or (_37143_, _37142_, _01012_);
  and (_43717_, _37143_, _41806_);
  and (_37144_, _43004_, \oc8051_golden_model_1.P3INREG [5]);
  or (_37145_, _37144_, _01052_);
  and (_43718_, _37145_, _41806_);
  and (_37146_, _43004_, \oc8051_golden_model_1.P3INREG [6]);
  or (_37147_, _37146_, _01003_);
  and (_43719_, _37147_, _41806_);
  nor (_00005_[6], _01004_, rst);
  nor (_00005_[5], _01053_, rst);
  nor (_00005_[4], _01013_, rst);
  nor (_00005_[3], _01036_, rst);
  nor (_00005_[2], _00997_, rst);
  nor (_00005_[1], _01046_, rst);
  nor (_00005_[0], _01020_, rst);
  nor (_00004_[6], _00882_, rst);
  nor (_00004_[5], _00934_, rst);
  nor (_00004_[4], _00892_, rst);
  nor (_00004_[3], _00917_, rst);
  nor (_00004_[2], _00875_, rst);
  nor (_00004_[1], _00927_, rst);
  nor (_00004_[0], _00900_, rst);
  nor (_00003_[6], _01111_, rst);
  nor (_00003_[5], _01077_, rst);
  nor (_00003_[4], _01127_, rst);
  nor (_00003_[3], _01100_, rst);
  nor (_00003_[2], _01118_, rst);
  nor (_00003_[1], _01084_, rst);
  nor (_00003_[0], _01134_, rst);
  nor (_00002_[6], _01180_, rst);
  nor (_00002_[5], _01147_, rst);
  nor (_00002_[4], _01163_, rst);
  nor (_00002_[3], _01203_, rst);
  nor (_00002_[2], _01187_, rst);
  nor (_00002_[1], _01154_, rst);
  nor (_00002_[0], _01170_, rst);
  or (_37151_, _10641_, _09230_);
  nor (_37152_, _37151_, _10903_);
  not (_37154_, _28767_);
  and (_37155_, _37154_, _28534_);
  nor (_37156_, _29111_, _28997_);
  and (_37157_, _37156_, _37155_);
  nor (_37158_, _27118_, _27001_);
  nor (_37159_, _27463_, _27349_);
  and (_37160_, _37159_, _37158_);
  nor (_37161_, _19863_, _19634_);
  nor (_37162_, _26885_, _19976_);
  and (_37163_, _37162_, _37161_);
  and (_37165_, _37163_, _37160_);
  and (_37166_, _37165_, _37157_);
  nor (_37167_, _11230_, _11148_);
  nor (_37168_, _18722_, _11311_);
  and (_37169_, _37168_, _37167_);
  nor (_37170_, _10533_, _10452_);
  nor (_37171_, _11066_, _10985_);
  and (_37172_, _37171_, _37170_);
  and (_37173_, _37172_, _37169_);
  not (_37174_, _26774_);
  nor (_37176_, _37174_, _19517_);
  not (_37177_, _28423_);
  nor (_37178_, _28650_, _37177_);
  nand (_37179_, _37178_, _37176_);
  nor (_37180_, _37179_, _18954_);
  and (_37181_, _37180_, _37173_);
  nor (_37182_, _19068_, _18839_);
  nor (_37183_, _19400_, _19182_);
  and (_37184_, _37183_, _37182_);
  or (_37185_, _31193_, _29972_);
  nor (_37187_, _37185_, _31800_);
  or (_37188_, _11764_, _03165_);
  nor (_37189_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor (_37190_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor (_37191_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and (_37192_, _37191_, _37190_);
  and (_37193_, _37192_, _37189_);
  nor (_37194_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_37195_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and (_37196_, _37195_, _37194_);
  nor (_37198_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor (_37199_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and (_37200_, _37199_, _37198_);
  and (_37201_, _37200_, _37196_);
  and (_37202_, _37201_, _37193_);
  nor (_37203_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor (_37204_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and (_37205_, _37204_, _37203_);
  nor (_37206_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor (_37207_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and (_37209_, _37207_, _37206_);
  and (_37210_, _37209_, _37205_);
  nor (_37211_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_37212_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and (_37213_, _37212_, _37211_);
  nor (_37214_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor (_37215_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and (_37216_, _37215_, _37214_);
  and (_37217_, _37216_, _37213_);
  and (_37218_, _37217_, _37210_);
  and (_37220_, _37218_, _37202_);
  nor (_37221_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_37222_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and (_37223_, _37222_, _37221_);
  nor (_37224_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor (_37225_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and (_37226_, _37225_, _37224_);
  and (_37227_, _37226_, _37223_);
  nor (_37228_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  nor (_37229_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  and (_37231_, _37229_, _37228_);
  nor (_37232_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor (_37233_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and (_37234_, _37233_, _37232_);
  and (_37235_, _37234_, _37231_);
  and (_37236_, _37235_, _37227_);
  nor (_37237_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_37238_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and (_37239_, _37238_, _37237_);
  nor (_37240_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  nor (_37242_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  and (_37243_, _37242_, _37240_);
  and (_37244_, _37243_, _37239_);
  nor (_37245_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor (_37246_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and (_37247_, _37246_, _37245_);
  nor (_37248_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor (_37249_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and (_37250_, _37249_, _37248_);
  and (_37251_, _37250_, _37247_);
  and (_37253_, _37251_, _37244_);
  and (_37254_, _37253_, _37236_);
  nor (_37255_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and (_37256_, _37255_, op0_cnst);
  nor (_37257_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor (_37258_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and (_37259_, _37258_, _37257_);
  nor (_37260_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor (_37261_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and (_37262_, _37261_, _37260_);
  and (_37264_, _37262_, _37259_);
  and (_37265_, _37264_, _37256_);
  nor (_37266_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_37267_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and (_37268_, _37267_, _37266_);
  nor (_37269_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor (_37270_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and (_37271_, _37270_, _37269_);
  and (_37272_, _37271_, _37268_);
  and (_37273_, \oc8051_golden_model_1.TCON [1], _28320_);
  nor (_37275_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and (_37276_, _37275_, _37273_);
  nor (_37277_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor (_37278_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and (_37279_, _37278_, _37277_);
  and (_37280_, _37279_, _37276_);
  and (_37281_, _37280_, _37272_);
  and (_37282_, _37281_, _37265_);
  and (_37283_, _37282_, _37254_);
  and (_37284_, _37283_, _37220_);
  nand (_37286_, _37284_, _37188_);
  nor (_37287_, _37286_, _25536_);
  nor (_37288_, _29192_, _26140_);
  and (_37289_, _37288_, _37287_);
  nor (_37290_, _26316_, _25712_);
  and (_37291_, _37290_, _37289_);
  and (_37292_, _37291_, _37187_);
  nor (_37293_, _26227_, _25623_);
  and (_37294_, _37293_, _37292_);
  nor (_37295_, _29884_, _29454_);
  nor (_37297_, _30586_, _30058_);
  and (_37298_, _37297_, _37295_);
  nor (_37299_, _30398_, _29799_);
  nor (_37300_, _31624_, _31016_);
  nand (_37301_, _37300_, _37299_);
  nor (_37302_, _37301_, _25798_);
  nor (_37303_, _29368_, _26403_);
  and (_37304_, _37303_, _37302_);
  and (_37305_, _37304_, _37298_);
  and (_37306_, _37305_, _37294_);
  nor (_37308_, _30497_, _29279_);
  nor (_37309_, _31711_, _31104_);
  nand (_37310_, _37309_, _37308_);
  nor (_37311_, _37310_, _19289_);
  and (_37312_, _37311_, _37306_);
  nor (_37313_, _29629_, _26666_);
  nor (_37314_, _30233_, _29716_);
  and (_37315_, _37314_, _37313_);
  or (_37316_, _31280_, _30672_);
  or (_37317_, _37316_, _31886_);
  nor (_37319_, _37317_, _25973_);
  nor (_37320_, _26579_, _26059_);
  and (_37321_, _37320_, _37319_);
  and (_37322_, _37321_, _37315_);
  and (_37323_, _37322_, _37312_);
  or (_37324_, _31369_, _30760_);
  nor (_37325_, _37324_, _31975_);
  nor (_37326_, _26492_, _25886_);
  nor (_37327_, _30146_, _29543_);
  and (_37328_, _37327_, _37326_);
  and (_37330_, _37328_, _37325_);
  and (_37331_, _37330_, _37323_);
  or (_37332_, _32061_, _31542_);
  nor (_37333_, _37332_, _32147_);
  nor (_37334_, _30846_, _30319_);
  nor (_37335_, _31456_, _30933_);
  and (_37336_, _37335_, _37334_);
  nand (_37337_, _37336_, _37333_);
  or (_37338_, _37337_, _18494_);
  nor (_37339_, _37338_, _18606_);
  and (_37341_, _37339_, _37331_);
  and (_37342_, _37341_, _37184_);
  and (_37343_, _37342_, _37181_);
  or (_37344_, _27234_, _19749_);
  or (_37345_, _37344_, _28882_);
  nor (_37346_, _37345_, _09123_);
  and (_37347_, _37346_, _37343_);
  and (_37348_, _37347_, _37166_);
  and (_37349_, _37348_, _37152_);
  and (_37350_, _37349_, _43000_);
  and (_37352_, _37350_, _41806_);
  nor (_37353_, _10796_, _38443_);
  and (_37354_, _10796_, _38443_);
  or (_37355_, _37354_, _37353_);
  and (_37356_, _28315_, _38487_);
  nor (_37357_, _28315_, _38487_);
  or (_37358_, _37357_, _37356_);
  and (_37359_, _28181_, _38481_);
  or (_37360_, _27548_, _40411_);
  nand (_37361_, _27548_, _40411_);
  and (_37363_, _37361_, _37360_);
  or (_37364_, _27668_, _38457_);
  nand (_37365_, _27668_, _38457_);
  and (_37366_, _37365_, _37364_);
  or (_37367_, _37366_, _37363_);
  and (_37368_, _27790_, _38463_);
  nor (_37369_, _27790_, _38463_);
  or (_37370_, _37369_, _37368_);
  or (_37371_, _37370_, _37367_);
  or (_37372_, _37371_, _37359_);
  nor (_37374_, _27912_, _38469_);
  and (_37375_, _27912_, _38469_);
  or (_37376_, _37375_, _37374_);
  or (_37377_, _28046_, _40511_);
  nand (_37378_, _28046_, _40511_);
  and (_37379_, _37378_, _37377_);
  nor (_37380_, _28181_, _38481_);
  or (_37381_, _37380_, _37379_);
  or (_37382_, _37381_, _37376_);
  or (_37383_, _37382_, _37372_);
  or (_37385_, _37383_, _37358_);
  or (_37386_, _37385_, _37355_);
  and (_00007_, _37386_, _37352_);
  nor (_37387_, _25047_, _40277_);
  and (_37388_, _25047_, _40277_);
  or (_37389_, _37388_, _37387_);
  and (_37390_, _25164_, _38949_);
  nor (_37391_, _25164_, _38949_);
  or (_37392_, _37391_, _37390_);
  or (_37393_, _37392_, _37389_);
  nor (_37395_, _24693_, _38864_);
  and (_37396_, _24693_, _38864_);
  or (_37397_, _37396_, _37395_);
  not (_37398_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_37399_, _25279_, _37398_);
  and (_37400_, _25279_, _37398_);
  or (_37401_, _37400_, _37399_);
  or (_37402_, _37401_, _37397_);
  or (_37403_, _37402_, _37393_);
  and (_37404_, _25455_, _31066_);
  nor (_37406_, _25455_, _31066_);
  or (_37407_, _37406_, _37404_);
  or (_37408_, _37407_, _37403_);
  and (_37409_, _24932_, _38901_);
  nor (_37410_, _24932_, _38901_);
  or (_37411_, _37410_, _37409_);
  or (_37412_, _37411_, _37408_);
  and (_37413_, _10371_, _38839_);
  nor (_37414_, _10371_, _38839_);
  or (_37415_, _37414_, _37413_);
  or (_37417_, _37415_, _37412_);
  and (_00006_, _37417_, _37352_);
  or (_00001_, _37349_, rst);
  nor (_00005_[7], _01029_, rst);
  nor (_00004_[7], _00909_, rst);
  nor (_00003_[7], _01093_, rst);
  nor (_00002_[7], _01196_, rst);
  and (_37418_, _37349_, inst_finished_r);
  nor (_37419_, _38443_, \oc8051_golden_model_1.SP [7]);
  and (_37420_, _38443_, \oc8051_golden_model_1.SP [7]);
  or (_37422_, _37420_, _37419_);
  nor (_37423_, _38487_, \oc8051_golden_model_1.SP [6]);
  and (_37424_, _38487_, \oc8051_golden_model_1.SP [6]);
  or (_37425_, _37424_, _37423_);
  nor (_37426_, _38481_, \oc8051_golden_model_1.SP [5]);
  and (_37427_, _38481_, \oc8051_golden_model_1.SP [5]);
  or (_37428_, _37427_, _37426_);
  nor (_37429_, _38469_, \oc8051_golden_model_1.SP [3]);
  and (_37430_, _38469_, \oc8051_golden_model_1.SP [3]);
  or (_37431_, _37430_, _37429_);
  and (_37433_, _38457_, \oc8051_golden_model_1.SP [1]);
  nor (_37434_, _38451_, \oc8051_golden_model_1.SP [0]);
  and (_37435_, _38451_, \oc8051_golden_model_1.SP [0]);
  or (_37436_, _37435_, _37434_);
  nor (_37437_, _38457_, \oc8051_golden_model_1.SP [1]);
  or (_37438_, _37437_, _37436_);
  or (_37439_, _37438_, _37433_);
  nor (_37440_, _38463_, \oc8051_golden_model_1.SP [2]);
  and (_37441_, _38463_, \oc8051_golden_model_1.SP [2]);
  or (_37442_, _37441_, _37440_);
  or (_37444_, _37442_, _37439_);
  or (_37445_, _37444_, _37431_);
  nor (_37446_, _38475_, \oc8051_golden_model_1.SP [4]);
  and (_37447_, _38475_, \oc8051_golden_model_1.SP [4]);
  or (_37448_, _37447_, _37446_);
  or (_37449_, _37448_, _37445_);
  or (_37450_, _37449_, _37428_);
  or (_37451_, _37450_, _37425_);
  or (_37452_, _37451_, _37422_);
  and (_37453_, _37452_, property_invalid_sp_1_r);
  and (property_invalid_sp, _37453_, _37418_);
  and (_37455_, _25052_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_37456_, \oc8051_golden_model_1.PSW [4], _38949_);
  or (_37457_, _37456_, _37455_);
  and (_37458_, _05018_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_37459_, \oc8051_golden_model_1.PSW [3], _40277_);
  or (_37460_, _37459_, _37458_);
  or (_37461_, _37460_, _37457_);
  and (_37462_, _24593_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_37463_, \oc8051_golden_model_1.PSW [1], _38864_);
  or (_37465_, _37463_, _37462_);
  nand (_37466_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_37467_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_37468_, _37467_, _37466_);
  or (_37469_, _37468_, _37465_);
  or (_37470_, _37469_, _37461_);
  and (_37471_, _07871_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_37472_, \oc8051_golden_model_1.PSW [7], _38839_);
  or (_37473_, _37472_, _37471_);
  and (_37474_, _25169_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_37476_, \oc8051_golden_model_1.PSW [5], _37398_);
  or (_37477_, _37476_, _37474_);
  nand (_37478_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_37479_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_37480_, _37479_, _37478_);
  or (_37481_, _37480_, _37477_);
  or (_37482_, _37481_, _37473_);
  or (_37483_, _37482_, _37470_);
  and (_37484_, _37483_, property_invalid_psw_1_r);
  and (property_invalid_psw, _37484_, _37418_);
  nand (_37486_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_37487_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_37488_, _37487_, _37486_);
  and (_37489_, _22590_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_37490_, \oc8051_golden_model_1.P3 [2], _39721_);
  or (_37491_, _37490_, _37489_);
  or (_37492_, _37491_, _37488_);
  and (_37493_, \oc8051_golden_model_1.P3 [0], _39688_);
  and (_37494_, _22373_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_37495_, _37494_, _37493_);
  and (_37497_, _22487_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_37498_, \oc8051_golden_model_1.P3 [1], _39701_);
  or (_37499_, _37498_, _37497_);
  or (_37500_, _37499_, _37495_);
  or (_37501_, _37500_, _37492_);
  or (_37502_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_37503_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_37504_, _37503_, _37502_);
  or (_37505_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_37506_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_37508_, _37506_, _37505_);
  or (_37509_, _37508_, _37504_);
  and (_37510_, _09553_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_37511_, \oc8051_golden_model_1.P3 [7], _39241_);
  or (_37512_, _37511_, _37510_);
  nand (_37513_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_37514_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_37515_, _37514_, _37513_);
  or (_37516_, _37515_, _37512_);
  or (_37517_, _37516_, _37509_);
  or (_37519_, _37517_, _37501_);
  and (property_invalid_p3, _37519_, _37418_);
  nand (_37520_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_37521_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_37522_, _37521_, _37520_);
  and (_37523_, _21818_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_37524_, \oc8051_golden_model_1.P2 [2], _39619_);
  or (_37525_, _37524_, _37523_);
  or (_37526_, _37525_, _37522_);
  and (_37527_, \oc8051_golden_model_1.P2 [0], _39592_);
  and (_37529_, _21602_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_37530_, _37529_, _37527_);
  and (_37531_, _21716_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_37532_, \oc8051_golden_model_1.P2 [1], _39605_);
  or (_37533_, _37532_, _37531_);
  or (_37534_, _37533_, _37530_);
  or (_37535_, _37534_, _37526_);
  or (_37536_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_37537_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_37538_, _37537_, _37536_);
  or (_37540_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_37541_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_37542_, _37541_, _37540_);
  or (_37543_, _37542_, _37538_);
  and (_37544_, _09450_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_37545_, \oc8051_golden_model_1.P2 [7], _39183_);
  or (_37546_, _37545_, _37544_);
  nand (_37547_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_37548_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_37549_, _37548_, _37547_);
  or (_37551_, _37549_, _37546_);
  or (_37552_, _37551_, _37543_);
  or (_37553_, _37552_, _37535_);
  and (property_invalid_p2, _37553_, _37418_);
  nand (_37554_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_37555_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_37556_, _37555_, _37554_);
  and (_37557_, _21045_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_37558_, \oc8051_golden_model_1.P1 [2], _39528_);
  or (_37559_, _37558_, _37557_);
  or (_37561_, _37559_, _37556_);
  and (_37562_, \oc8051_golden_model_1.P1 [0], _39502_);
  and (_37563_, _20834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_37564_, _37563_, _37562_);
  and (_37565_, _20944_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_37566_, \oc8051_golden_model_1.P1 [1], _39515_);
  or (_37567_, _37566_, _37565_);
  or (_37568_, _37567_, _37564_);
  or (_37569_, _37568_, _37561_);
  or (_37570_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_37572_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_37573_, _37572_, _37570_);
  or (_37574_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_37575_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_37576_, _37575_, _37574_);
  or (_37577_, _37576_, _37573_);
  and (_37578_, _09348_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_37579_, \oc8051_golden_model_1.P1 [7], _39165_);
  or (_37580_, _37579_, _37578_);
  nand (_37581_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_37583_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_37584_, _37583_, _37581_);
  or (_37585_, _37584_, _37580_);
  or (_37586_, _37585_, _37577_);
  or (_37587_, _37586_, _37569_);
  and (property_invalid_p1, _37587_, _37418_);
  nand (_37588_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_37589_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_37590_, _37589_, _37588_);
  and (_37591_, _20223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_37593_, \oc8051_golden_model_1.P0 [2], _39438_);
  or (_37594_, _37593_, _37591_);
  or (_37595_, _37594_, _37590_);
  and (_37596_, \oc8051_golden_model_1.P0 [0], _39327_);
  and (_37597_, _19980_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_37598_, _37597_, _37596_);
  and (_37599_, _20107_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_37600_, \oc8051_golden_model_1.P0 [1], _39422_);
  or (_37601_, _37600_, _37599_);
  or (_37602_, _37601_, _37598_);
  or (_37604_, _37602_, _37595_);
  or (_37605_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_37606_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_37607_, _37606_, _37605_);
  or (_37608_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand (_37609_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_37610_, _37609_, _37608_);
  or (_37611_, _37610_, _37607_);
  and (_37612_, _09234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_37613_, \oc8051_golden_model_1.P0 [7], _39151_);
  or (_37615_, _37613_, _37612_);
  nand (_37616_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_37617_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_37618_, _37617_, _37616_);
  or (_37619_, _37618_, _37615_);
  or (_37620_, _37619_, _37611_);
  or (_37621_, _37620_, _37604_);
  and (property_invalid_p0, _37621_, _37418_);
  or (_37622_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nand (_37623_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_37625_, _37623_, _37622_);
  or (_37626_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_37627_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_37628_, _37627_, _37626_);
  or (_37629_, _37628_, _37625_);
  and (_37630_, \oc8051_golden_model_1.IRAM[0] [0], _40890_);
  and (_37631_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_37632_, _37631_, _37630_);
  and (_37633_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_37634_, \oc8051_golden_model_1.IRAM[0] [1], _40903_);
  or (_37636_, _37634_, _37633_);
  or (_37637_, _37636_, _37632_);
  or (_37638_, _37637_, _37629_);
  or (_37639_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand (_37640_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_37641_, _37640_, _37639_);
  or (_37642_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand (_37643_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_37644_, _37643_, _37642_);
  or (_37645_, _37644_, _37641_);
  or (_37647_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_37648_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_37649_, _37648_, _37647_);
  or (_37650_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand (_37651_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_37652_, _37651_, _37650_);
  or (_37653_, _37652_, _37649_);
  or (_37654_, _37653_, _37645_);
  or (_37655_, _37654_, _37638_);
  or (_37656_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_37658_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_37659_, _37658_, _37656_);
  or (_37660_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_37661_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_37662_, _37661_, _37660_);
  or (_37663_, _37662_, _37659_);
  or (_37664_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand (_37665_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_37666_, _37665_, _37664_);
  or (_37667_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nand (_37669_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_37670_, _37669_, _37667_);
  or (_37671_, _37670_, _37666_);
  or (_37672_, _37671_, _37663_);
  and (_37673_, _05723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_37674_, \oc8051_golden_model_1.IRAM[1] [4], _40974_);
  or (_37675_, _37674_, _37673_);
  and (_37676_, \oc8051_golden_model_1.IRAM[1] [5], _40978_);
  and (_37677_, _05415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_37678_, _37677_, _37676_);
  or (_37680_, _37678_, _37675_);
  or (_37681_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand (_37682_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_37683_, _37682_, _37681_);
  or (_37684_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nand (_37685_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_37686_, _37685_, _37684_);
  or (_37687_, _37686_, _37683_);
  or (_37688_, _37687_, _37680_);
  or (_37689_, _37688_, _37672_);
  or (_37691_, _37689_, _37655_);
  or (_37692_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand (_37693_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_37694_, _37693_, _37692_);
  or (_37695_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand (_37696_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_37697_, _37696_, _37695_);
  or (_37698_, _37697_, _37694_);
  or (_37699_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nand (_37700_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_37702_, _37700_, _37699_);
  and (_37703_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_37704_, \oc8051_golden_model_1.IRAM[2] [2], _40993_);
  or (_37705_, _37704_, _37703_);
  or (_37706_, _37705_, _37702_);
  or (_37707_, _37706_, _37698_);
  and (_37708_, _05729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_37709_, \oc8051_golden_model_1.IRAM[2] [4], _40998_);
  or (_37710_, _37709_, _37708_);
  and (_37711_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_37713_, \oc8051_golden_model_1.IRAM[2] [5], _41001_);
  or (_37714_, _37713_, _37711_);
  or (_37715_, _37714_, _37710_);
  or (_37716_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nand (_37717_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_37718_, _37717_, _37716_);
  and (_37719_, \oc8051_golden_model_1.IRAM[2] [7], _41006_);
  and (_37720_, _05152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_37721_, _37720_, _37719_);
  or (_37722_, _37721_, _37718_);
  or (_37724_, _37722_, _37715_);
  or (_37725_, _37724_, _37707_);
  and (_37726_, \oc8051_golden_model_1.IRAM[3] [2], _41016_);
  and (_37727_, _04825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_37728_, _37727_, _37726_);
  nand (_37729_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_37730_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_37731_, _37730_, _37729_);
  or (_37732_, _37731_, _37728_);
  and (_37733_, _04569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_37735_, \oc8051_golden_model_1.IRAM[3] [0], _41010_);
  or (_37736_, _37735_, _37733_);
  and (_37737_, \oc8051_golden_model_1.IRAM[3] [1], _41013_);
  and (_37738_, _04352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_37739_, _37738_, _37737_);
  or (_37740_, _37739_, _37736_);
  or (_37741_, _37740_, _37732_);
  or (_37742_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nand (_37743_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_37744_, _37743_, _37742_);
  and (_37746_, _05150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_37747_, \oc8051_golden_model_1.IRAM[3] [7], _40758_);
  or (_37748_, _37747_, _37746_);
  or (_37749_, _37748_, _37744_);
  or (_37750_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_37751_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_37752_, _37751_, _37750_);
  or (_37753_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_37754_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_37755_, _37754_, _37753_);
  or (_37757_, _37755_, _37752_);
  or (_37758_, _37757_, _37749_);
  or (_37759_, _37758_, _37741_);
  or (_37760_, _37759_, _37725_);
  or (_37761_, _37760_, _37691_);
  and (_37762_, _04584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_37763_, \oc8051_golden_model_1.IRAM[4] [0], _41033_);
  or (_37764_, _37763_, _37762_);
  and (_37765_, \oc8051_golden_model_1.IRAM[4] [1], _41036_);
  and (_37766_, _04368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_37768_, _37766_, _37765_);
  or (_37769_, _37768_, _37764_);
  or (_37770_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand (_37771_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_37772_, _37771_, _37770_);
  nand (_37773_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_37774_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_37775_, _37774_, _37773_);
  or (_37776_, _37775_, _37772_);
  or (_37777_, _37776_, _37769_);
  or (_37779_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand (_37780_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_37781_, _37780_, _37779_);
  or (_37782_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand (_37783_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_37784_, _37783_, _37782_);
  or (_37785_, _37784_, _37781_);
  or (_37786_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand (_37787_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_37788_, _37787_, _37786_);
  nand (_37790_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_37791_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_37792_, _37791_, _37790_);
  or (_37793_, _37792_, _37788_);
  or (_37794_, _37793_, _37785_);
  or (_37795_, _37794_, _37777_);
  or (_37796_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand (_37797_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_37798_, _37797_, _37796_);
  nand (_37799_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_37801_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_37802_, _37801_, _37799_);
  or (_37803_, _37802_, _37798_);
  or (_37804_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_37805_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_37806_, _37805_, _37804_);
  or (_37807_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_37808_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_37809_, _37808_, _37807_);
  or (_37810_, _37809_, _37806_);
  or (_37812_, _37810_, _37803_);
  or (_37813_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand (_37814_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_37815_, _37814_, _37813_);
  nand (_37816_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_37817_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_37818_, _37817_, _37816_);
  or (_37819_, _37818_, _37815_);
  and (_37820_, _05743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_37821_, \oc8051_golden_model_1.IRAM[5] [4], _41063_);
  or (_37823_, _37821_, _37820_);
  and (_37824_, _05435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_37825_, \oc8051_golden_model_1.IRAM[5] [5], _41066_);
  or (_37826_, _37825_, _37824_);
  or (_37827_, _37826_, _37823_);
  or (_37828_, _37827_, _37819_);
  or (_37829_, _37828_, _37812_);
  or (_37830_, _37829_, _37795_);
  nand (_37831_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_37832_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_37834_, _37832_, _37831_);
  and (_37835_, \oc8051_golden_model_1.IRAM[6] [2], _41080_);
  and (_37836_, _04835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_37837_, _37836_, _37835_);
  or (_37838_, _37837_, _37834_);
  or (_37839_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand (_37840_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_37841_, _37840_, _37839_);
  or (_37842_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand (_37843_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_37845_, _37843_, _37842_);
  or (_37846_, _37845_, _37841_);
  or (_37847_, _37846_, _37838_);
  and (_37848_, _05160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_37849_, \oc8051_golden_model_1.IRAM[6] [7], _41094_);
  or (_37850_, _37849_, _37848_);
  nand (_37851_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_37852_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_37853_, _37852_, _37851_);
  or (_37854_, _37853_, _37850_);
  and (_37856_, _05737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_37857_, \oc8051_golden_model_1.IRAM[6] [4], _41085_);
  or (_37858_, _37857_, _37856_);
  and (_37859_, \oc8051_golden_model_1.IRAM[6] [5], _41088_);
  and (_37860_, _05429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_37861_, _37860_, _37859_);
  or (_37862_, _37861_, _37858_);
  or (_37863_, _37862_, _37854_);
  or (_37864_, _37863_, _37847_);
  and (_37865_, _04362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37867_, \oc8051_golden_model_1.IRAM[7] [1], _41101_);
  or (_37868_, _37867_, _37865_);
  and (_37869_, _04578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_37870_, \oc8051_golden_model_1.IRAM[7] [0], _41098_);
  or (_37871_, _37870_, _37869_);
  or (_37872_, _37871_, _37868_);
  and (_37873_, _04833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_37874_, \oc8051_golden_model_1.IRAM[7] [2], _41104_);
  or (_37875_, _37874_, _37873_);
  nand (_37876_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_37878_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_37879_, _37878_, _37876_);
  or (_37880_, _37879_, _37875_);
  or (_37881_, _37880_, _37872_);
  or (_37882_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_37883_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_37884_, _37883_, _37882_);
  or (_37885_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_37886_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_37887_, _37886_, _37885_);
  or (_37889_, _37887_, _37884_);
  nand (_37890_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_37891_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_37892_, _37891_, _37890_);
  and (_37893_, _05158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_37894_, \oc8051_golden_model_1.IRAM[7] [7], _40794_);
  or (_37895_, _37894_, _37893_);
  or (_37896_, _37895_, _37892_);
  or (_37897_, _37896_, _37889_);
  or (_37898_, _37897_, _37881_);
  or (_37900_, _37898_, _37864_);
  or (_37901_, _37900_, _37830_);
  or (_37902_, _37901_, _37761_);
  and (_37903_, _04599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_37904_, \oc8051_golden_model_1.IRAM[8] [0], _41121_);
  or (_37905_, _37904_, _37903_);
  and (_37906_, \oc8051_golden_model_1.IRAM[8] [1], _41124_);
  and (_37907_, _04385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_37908_, _37907_, _37906_);
  or (_37909_, _37908_, _37905_);
  or (_37911_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand (_37912_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_37913_, _37912_, _37911_);
  nand (_37914_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_37915_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_37916_, _37915_, _37914_);
  or (_37917_, _37916_, _37913_);
  or (_37918_, _37917_, _37909_);
  or (_37919_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nand (_37920_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_37922_, _37920_, _37919_);
  or (_37923_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nand (_37924_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_37925_, _37924_, _37923_);
  or (_37926_, _37925_, _37922_);
  or (_37927_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_37928_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_37929_, _37928_, _37927_);
  nand (_37930_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_37931_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_37933_, _37931_, _37930_);
  or (_37934_, _37933_, _37929_);
  or (_37935_, _37934_, _37926_);
  or (_37936_, _37935_, _37918_);
  or (_37937_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand (_37938_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_37939_, _37938_, _37937_);
  nand (_37940_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_37941_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_37942_, _37941_, _37940_);
  or (_37944_, _37942_, _37939_);
  or (_37945_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand (_37946_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_37947_, _37946_, _37945_);
  or (_37948_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nand (_37949_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_37950_, _37949_, _37948_);
  or (_37951_, _37950_, _37947_);
  or (_37952_, _37951_, _37944_);
  and (_37953_, _05449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_37955_, \oc8051_golden_model_1.IRAM[9] [5], _41155_);
  or (_37956_, _37955_, _37953_);
  and (_37957_, _05757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_37958_, \oc8051_golden_model_1.IRAM[9] [4], _41152_);
  or (_37959_, _37958_, _37957_);
  or (_37960_, _37959_, _37956_);
  or (_37961_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand (_37962_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_37963_, _37962_, _37961_);
  nand (_37964_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_37966_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_37967_, _37966_, _37964_);
  or (_37968_, _37967_, _37963_);
  or (_37969_, _37968_, _37960_);
  or (_37970_, _37969_, _37952_);
  or (_37971_, _37970_, _37936_);
  and (_37972_, _04851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_37973_, \oc8051_golden_model_1.IRAM[10] [2], _41168_);
  or (_37974_, _37973_, _37972_);
  nand (_37975_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_37976_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_37977_, _37976_, _37975_);
  or (_37978_, _37977_, _37974_);
  or (_37979_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nand (_37980_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_37981_, _37980_, _37979_);
  or (_37982_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nand (_37983_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_37984_, _37983_, _37982_);
  or (_37985_, _37984_, _37981_);
  or (_37987_, _37985_, _37978_);
  and (_37988_, \oc8051_golden_model_1.IRAM[10] [7], _40831_);
  and (_37989_, _05176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_37990_, _37989_, _37988_);
  nand (_37991_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_37992_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_37993_, _37992_, _37991_);
  or (_37994_, _37993_, _37990_);
  and (_37995_, _05752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_37996_, \oc8051_golden_model_1.IRAM[10] [4], _41174_);
  or (_37998_, _37996_, _37995_);
  and (_37999_, \oc8051_golden_model_1.IRAM[10] [5], _41177_);
  and (_38000_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_38001_, _38000_, _37999_);
  or (_38002_, _38001_, _37998_);
  or (_38003_, _38002_, _37994_);
  or (_38004_, _38003_, _37987_);
  and (_38005_, _04594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_38006_, \oc8051_golden_model_1.IRAM[11] [0], _41186_);
  or (_38007_, _38006_, _38005_);
  and (_38009_, \oc8051_golden_model_1.IRAM[11] [1], _41189_);
  and (_38010_, _04380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_38011_, _38010_, _38009_);
  or (_38012_, _38011_, _38007_);
  and (_38013_, \oc8051_golden_model_1.IRAM[11] [2], _41192_);
  and (_38014_, _04849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_38015_, _38014_, _38013_);
  nand (_38016_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_38017_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_38018_, _38017_, _38016_);
  or (_38020_, _38018_, _38015_);
  or (_38021_, _38020_, _38012_);
  or (_38022_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_38023_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_38024_, _38023_, _38022_);
  or (_38025_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_38026_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_38027_, _38026_, _38025_);
  or (_38028_, _38027_, _38024_);
  and (_38029_, _05174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_38031_, \oc8051_golden_model_1.IRAM[11] [7], _41204_);
  or (_38032_, _38031_, _38029_);
  nand (_38033_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_38034_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_38035_, _38034_, _38033_);
  or (_38036_, _38035_, _38032_);
  or (_38037_, _38036_, _38028_);
  or (_38038_, _38037_, _38021_);
  or (_38039_, _38038_, _38004_);
  or (_38040_, _38039_, _37971_);
  or (_38042_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand (_38043_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_38044_, _38043_, _38042_);
  nand (_38045_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_38046_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_38047_, _38046_, _38045_);
  or (_38048_, _38047_, _38044_);
  and (_38049_, \oc8051_golden_model_1.IRAM[12] [1], _41217_);
  and (_38050_, _04397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_38051_, _38050_, _38049_);
  and (_38053_, _04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_38054_, \oc8051_golden_model_1.IRAM[12] [0], _41210_);
  or (_38055_, _38054_, _38053_);
  or (_38056_, _38055_, _38051_);
  or (_38057_, _38056_, _38048_);
  or (_38058_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_38059_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_38060_, _38059_, _38058_);
  nand (_38061_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_38062_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_38064_, _38062_, _38061_);
  or (_38065_, _38064_, _38060_);
  or (_38066_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nand (_38067_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_38068_, _38067_, _38066_);
  or (_38069_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nand (_38070_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_38071_, _38070_, _38069_);
  or (_38072_, _38071_, _38068_);
  or (_38073_, _38072_, _38065_);
  or (_38075_, _38073_, _38057_);
  or (_38076_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand (_38077_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_38078_, _38077_, _38076_);
  or (_38079_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nand (_38080_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_38081_, _38080_, _38079_);
  or (_38082_, _38081_, _38078_);
  or (_38083_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand (_38084_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_38086_, _38084_, _38083_);
  nand (_38087_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_38088_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_38089_, _38088_, _38087_);
  or (_38090_, _38089_, _38086_);
  or (_38091_, _38090_, _38082_);
  and (_38092_, _05769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_38093_, \oc8051_golden_model_1.IRAM[13] [4], _41267_);
  or (_38094_, _38093_, _38092_);
  and (_38095_, \oc8051_golden_model_1.IRAM[13] [5], _41270_);
  and (_38097_, _05461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_38098_, _38097_, _38095_);
  or (_38099_, _38098_, _38094_);
  or (_38100_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand (_38101_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_38102_, _38101_, _38100_);
  nand (_38103_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_38104_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_38105_, _38104_, _38103_);
  or (_38106_, _38105_, _38102_);
  or (_38108_, _38106_, _38099_);
  or (_38109_, _38108_, _38091_);
  or (_38110_, _38109_, _38075_);
  or (_38111_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nand (_38112_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_38113_, _38112_, _38111_);
  or (_38114_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nand (_38115_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_38116_, _38115_, _38114_);
  or (_38117_, _38116_, _38113_);
  and (_38119_, \oc8051_golden_model_1.IRAM[14] [2], _41283_);
  and (_38120_, _04863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_38121_, _38120_, _38119_);
  nand (_38122_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_38123_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_38124_, _38123_, _38122_);
  or (_38125_, _38124_, _38121_);
  or (_38126_, _38125_, _38117_);
  and (_38127_, \oc8051_golden_model_1.IRAM[14] [5], _41292_);
  and (_38128_, _05456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_38130_, _38128_, _38127_);
  and (_38131_, _05764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_38132_, \oc8051_golden_model_1.IRAM[14] [4], _41289_);
  or (_38133_, _38132_, _38131_);
  or (_38134_, _38133_, _38130_);
  and (_38135_, _05190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_38136_, \oc8051_golden_model_1.IRAM[14] [7], _40842_);
  or (_38137_, _38136_, _38135_);
  nand (_38138_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_38139_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_38141_, _38139_, _38138_);
  or (_38142_, _38141_, _38137_);
  or (_38143_, _38142_, _38134_);
  or (_38144_, _38143_, _38126_);
  and (_38145_, _04861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_38146_, \oc8051_golden_model_1.IRAM[15] [2], _41306_);
  or (_38147_, _38146_, _38145_);
  nand (_38148_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_38149_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_38150_, _38149_, _38148_);
  or (_38152_, _38150_, _38147_);
  and (_38153_, _04606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_38154_, \oc8051_golden_model_1.IRAM[15] [0], _41300_);
  or (_38155_, _38154_, _38153_);
  and (_38156_, _04392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_38157_, \oc8051_golden_model_1.IRAM[15] [1], _41303_);
  or (_38158_, _38157_, _38156_);
  or (_38159_, _38158_, _38155_);
  or (_38160_, _38159_, _38152_);
  and (_38161_, \oc8051_golden_model_1.IRAM[15] [7], _40873_);
  and (_38163_, _05188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_38164_, _38163_, _38161_);
  nand (_38165_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_38166_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_38167_, _38166_, _38165_);
  or (_38168_, _38167_, _38164_);
  or (_38169_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_38170_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_38171_, _38170_, _38169_);
  or (_38172_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_38174_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_38175_, _38174_, _38172_);
  or (_38176_, _38175_, _38171_);
  or (_38177_, _38176_, _38168_);
  or (_38178_, _38177_, _38160_);
  or (_38179_, _38178_, _38144_);
  or (_38180_, _38179_, _38110_);
  or (_38181_, _38180_, _38040_);
  or (_38182_, _38181_, _37902_);
  and (property_invalid_iram, _38182_, _37418_);
  nand (_38184_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38185_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_38186_, _38185_, _38184_);
  and (_38187_, _17923_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_38188_, _17923_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38189_, _38188_, _38187_);
  or (_38190_, _38189_, _38186_);
  nor (_38191_, _17740_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_38192_, _17740_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38193_, _38192_, _38191_);
  and (_38195_, _17829_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_38196_, _17829_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38197_, _38196_, _38195_);
  or (_38198_, _38197_, _38193_);
  or (_38199_, _38198_, _38190_);
  or (_38200_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_38201_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_38202_, _38201_, _38200_);
  or (_38203_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_38204_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_38206_, _38204_, _38203_);
  or (_38207_, _38206_, _38202_);
  and (_38208_, _08918_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_38209_, _08918_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38210_, _38209_, _38208_);
  nand (_38211_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38212_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_38213_, _38212_, _38211_);
  or (_38214_, _38213_, _38210_);
  or (_38215_, _38214_, _38207_);
  or (_38217_, _38215_, _38199_);
  and (property_invalid_dph, _38217_, _37418_);
  nand (_38218_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_38219_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38220_, _38219_, _38218_);
  and (_38221_, _17271_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38222_, \oc8051_golden_model_1.DPL [2], _38799_);
  or (_38223_, _38222_, _38221_);
  or (_38224_, _38223_, _38220_);
  and (_38225_, \oc8051_golden_model_1.DPL [0], _38791_);
  and (_38227_, _17089_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_38228_, _38227_, _38225_);
  and (_38229_, _17177_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38230_, \oc8051_golden_model_1.DPL [1], _38795_);
  or (_38231_, _38230_, _38229_);
  or (_38232_, _38231_, _38228_);
  or (_38233_, _38232_, _38224_);
  or (_38234_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_38235_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38236_, _38235_, _38234_);
  or (_38238_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_38239_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38240_, _38239_, _38238_);
  or (_38241_, _38240_, _38236_);
  and (_38242_, _08821_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38243_, \oc8051_golden_model_1.DPL [7], _38590_);
  or (_38244_, _38243_, _38242_);
  nand (_38245_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_38246_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38247_, _38246_, _38245_);
  or (_38249_, _38247_, _38244_);
  or (_38250_, _38249_, _38241_);
  or (_38251_, _38250_, _38233_);
  and (property_invalid_dpl, _38251_, _37418_);
  nand (_38252_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_38253_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_38254_, _38253_, _38252_);
  and (_38255_, _07426_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_38256_, \oc8051_golden_model_1.B [2], _30599_);
  or (_38257_, _38256_, _38255_);
  or (_38259_, _38257_, _38254_);
  and (_38260_, \oc8051_golden_model_1.B [0], _29264_);
  and (_38261_, _07418_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_38262_, _38261_, _38260_);
  and (_38263_, _07412_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_38264_, \oc8051_golden_model_1.B [1], _29926_);
  or (_38265_, _38264_, _38263_);
  or (_38266_, _38265_, _38262_);
  or (_38267_, _38266_, _38259_);
  or (_38268_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_38270_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_38271_, _38270_, _38268_);
  or (_38272_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_38273_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_38274_, _38273_, _38272_);
  or (_38275_, _38274_, _38271_);
  and (_38276_, _06826_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_38277_, \oc8051_golden_model_1.B [7], _28098_);
  or (_38278_, _38277_, _38276_);
  nand (_38279_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_38281_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_38282_, _38281_, _38279_);
  or (_38283_, _38282_, _38278_);
  or (_38284_, _38283_, _38275_);
  or (_38285_, _38284_, _38267_);
  and (property_invalid_b_reg, _38285_, _37418_);
  nand (_38286_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38287_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38288_, _38287_, _38286_);
  and (_38289_, _07584_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_38291_, \oc8051_golden_model_1.ACC [2], _39082_);
  or (_38292_, _38291_, _38289_);
  or (_38293_, _38292_, _38288_);
  nor (_38294_, _03274_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38295_, _03274_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_38296_, _38295_, _38294_);
  and (_38297_, _03335_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38298_, _03335_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_38299_, _38298_, _38297_);
  or (_38300_, _38299_, _38296_);
  or (_38302_, _38300_, _38293_);
  or (_38303_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38304_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38305_, _38304_, _38303_);
  or (_38306_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_38307_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38308_, _38307_, _38306_);
  or (_38309_, _38308_, _38305_);
  and (_38310_, _07433_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_38311_, _07433_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_38313_, _38311_, _38310_);
  nand (_38314_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38315_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_38316_, _38315_, _38314_);
  or (_38317_, _38316_, _38313_);
  or (_38318_, _38317_, _38309_);
  or (_38319_, _38318_, _38302_);
  and (property_invalid_acc, _38319_, _37418_);
  and (_38320_, _32793_, _43931_);
  nor (_38321_, _32793_, _43931_);
  and (_38323_, _33139_, _43935_);
  nor (_38324_, _33139_, _43935_);
  and (_38325_, _33488_, _43939_);
  and (_38326_, _35539_, _38549_);
  nor (_38327_, _35539_, _38549_);
  nor (_38328_, _11981_, _38571_);
  nor (_38329_, _36772_, _38535_);
  and (_38330_, _11981_, _38571_);
  or (_38331_, _38330_, _38329_);
  or (_38332_, _38331_, _38328_);
  nand (_38334_, _35205_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_38335_, _35205_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38336_, _38335_, _38334_);
  nor (_38337_, _36160_, _38539_);
  and (_38338_, _35846_, _38554_);
  nor (_38339_, _35846_, _38554_);
  and (_38340_, _36468_, _38560_);
  nand (_38341_, _32414_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_38342_, _32414_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_38343_, _38342_, _38341_);
  nor (_38345_, _36468_, _38560_);
  or (_38346_, _38345_, _38343_);
  or (_38347_, _38346_, _38340_);
  and (_38348_, _37080_, _38566_);
  nor (_38349_, _37080_, _38566_);
  or (_38350_, _38349_, _38348_);
  or (_38351_, _38350_, _38347_);
  or (_38352_, _38351_, _38339_);
  or (_38353_, _38352_, _38338_);
  or (_38354_, _38353_, _38337_);
  and (_38356_, _36160_, _38539_);
  and (_38357_, _36772_, _38535_);
  or (_38358_, _38357_, _38356_);
  or (_38359_, _38358_, _38354_);
  or (_38360_, _38359_, _38336_);
  or (_38361_, _38360_, _38332_);
  or (_38362_, _38361_, _38327_);
  or (_38363_, _38362_, _38326_);
  or (_38364_, _38363_, _38325_);
  or (_38365_, _38364_, _38324_);
  or (_38367_, _38365_, _38323_);
  nor (_38368_, _34187_, _43947_);
  nor (_38369_, _34887_, _43955_);
  and (_38370_, _34187_, _43947_);
  or (_38371_, _38370_, _38369_);
  or (_38372_, _38371_, _38368_);
  nor (_38373_, _33488_, _43939_);
  and (_38374_, _33837_, _43943_);
  or (_38375_, _38374_, _38373_);
  nor (_38376_, _33837_, _43943_);
  and (_38378_, _34887_, _43955_);
  or (_38379_, _38378_, _38376_);
  or (_38380_, _38379_, _38375_);
  or (_38381_, _38380_, _38372_);
  or (_38382_, _38381_, _38367_);
  nor (_38383_, _34533_, _43951_);
  and (_38384_, _34533_, _43951_);
  or (_38385_, _38384_, _38383_);
  or (_38386_, _38385_, _38382_);
  or (_38387_, _38386_, _38321_);
  or (_38389_, _38387_, _38320_);
  and (property_invalid_pc, _38389_, _37350_);
  buf (_01429_, _41806_);
  buf (_01480_, _41806_);
  buf (_01532_, _41806_);
  buf (_01584_, _41806_);
  buf (_01629_, _41806_);
  buf (_01675_, _41806_);
  buf (_01728_, _41806_);
  buf (_01779_, _41806_);
  buf (_01831_, _41806_);
  buf (_01883_, _41806_);
  buf (_01935_, _41806_);
  buf (_01987_, _41806_);
  buf (_02039_, _41806_);
  buf (_02091_, _41806_);
  buf (_02143_, _41806_);
  buf (_02195_, _41806_);
  buf (_38916_, _38813_);
  buf (_38917_, _38814_);
  buf (_38930_, _38813_);
  buf (_38931_, _38814_);
  buf (_39244_, _38832_);
  buf (_39245_, _38834_);
  buf (_39246_, _38835_);
  buf (_39247_, _38836_);
  buf (_39248_, _38837_);
  buf (_39249_, _38838_);
  buf (_39250_, _38840_);
  buf (_39252_, _38841_);
  buf (_39253_, _38842_);
  buf (_39254_, _38843_);
  buf (_39255_, _38844_);
  buf (_39256_, _38846_);
  buf (_39257_, _38847_);
  buf (_39258_, _38848_);
  buf (_39310_, _38832_);
  buf (_39311_, _38834_);
  buf (_39312_, _38835_);
  buf (_39313_, _38836_);
  buf (_39314_, _38837_);
  buf (_39315_, _38838_);
  buf (_39316_, _38840_);
  buf (_39317_, _38841_);
  buf (_39318_, _38842_);
  buf (_39319_, _38843_);
  buf (_39320_, _38844_);
  buf (_39321_, _38846_);
  buf (_39322_, _38847_);
  buf (_39323_, _38848_);
  buf (_39651_, _39617_);
  buf (_39766_, _39617_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (property_invalid_psw_1_r, _00006_);
  dff (property_invalid_sp_1_r, _00007_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _01433_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _01437_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _01441_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _01444_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _01448_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _01452_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _01456_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _01426_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _01429_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _01484_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _01488_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _01492_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _01496_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _01500_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _01504_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _01508_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _01477_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _01480_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _01939_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _01943_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _01947_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _01951_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _01955_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _01959_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _01963_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _01932_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _01935_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _01991_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _01995_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _01999_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _02003_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _02007_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _02011_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _02015_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _01984_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _01987_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _02043_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _02047_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _02051_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _02055_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _02059_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _02063_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _02067_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _02036_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _02039_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _02095_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _02099_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _02103_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _02107_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _02111_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _02115_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _02119_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _02088_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _02091_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _02147_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _02151_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _02155_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _02159_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _02163_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _02167_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _02171_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _02140_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _02143_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _02199_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _02203_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _02207_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _02211_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _02215_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _02219_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _02223_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _02192_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _02195_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _01536_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _01540_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _01544_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _01548_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _01552_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _01555_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _01559_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _01529_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _01532_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _01588_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _01591_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _01595_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _01599_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _01603_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _01607_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _01611_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _01581_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _01584_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _01630_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _01631_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _01634_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _01638_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _01642_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _01646_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _01650_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _01628_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _01629_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _01679_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _01683_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _01687_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _01691_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _01695_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _01699_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _01703_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _01672_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _01675_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _01732_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _01736_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _01740_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _01743_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _01747_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _01751_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _01755_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _01725_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _01728_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _01783_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _01787_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _01791_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _01795_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _01799_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _01803_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _01807_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _01777_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _01779_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _01835_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _01839_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _01843_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _01847_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _01851_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _01854_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _01858_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _01828_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _01831_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _01887_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _01891_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _01895_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _01899_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _01903_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _01907_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _01910_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _01880_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _01883_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _40819_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _40821_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _40822_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _40823_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _40824_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _40825_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _40827_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40565_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _40807_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _40809_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _40810_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _40811_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _40812_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _40813_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _40815_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _40816_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _40795_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _40796_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _40798_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _40799_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _40800_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _40801_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _40802_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _40804_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40783_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40784_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40786_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40787_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40788_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40789_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40790_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40792_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40771_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40772_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40773_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40774_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40776_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40777_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40778_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40779_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40759_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40760_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40761_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40762_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40764_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40765_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40766_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40767_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40747_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40748_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40749_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40750_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40751_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40753_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40754_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40755_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40735_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40736_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40737_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40738_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40739_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40741_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40742_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40743_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40722_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40723_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40724_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40725_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40727_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40728_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40729_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40730_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40710_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40711_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40712_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40713_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40715_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40716_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40717_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40718_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40698_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40699_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40700_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40701_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40702_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40704_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40705_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40706_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40686_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40687_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40688_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40689_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40690_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40692_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40693_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40694_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40673_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40674_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40675_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40676_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40678_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40679_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40680_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40681_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40661_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40662_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40663_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40664_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40665_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40667_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40668_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40669_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40648_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40649_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40650_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40651_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40653_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40654_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40655_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40656_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40634_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40635_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40637_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40638_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40640_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40641_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40642_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40644_);
  dff (\oc8051_golden_model_1.B [0], _43480_);
  dff (\oc8051_golden_model_1.B [1], _43481_);
  dff (\oc8051_golden_model_1.B [2], _43482_);
  dff (\oc8051_golden_model_1.B [3], _43485_);
  dff (\oc8051_golden_model_1.B [4], _43486_);
  dff (\oc8051_golden_model_1.B [5], _43487_);
  dff (\oc8051_golden_model_1.B [6], _43488_);
  dff (\oc8051_golden_model_1.B [7], _40566_);
  dff (\oc8051_golden_model_1.ACC [0], _43491_);
  dff (\oc8051_golden_model_1.ACC [1], _43492_);
  dff (\oc8051_golden_model_1.ACC [2], _43493_);
  dff (\oc8051_golden_model_1.ACC [3], _43494_);
  dff (\oc8051_golden_model_1.ACC [4], _43495_);
  dff (\oc8051_golden_model_1.ACC [5], _43496_);
  dff (\oc8051_golden_model_1.ACC [6], _43497_);
  dff (\oc8051_golden_model_1.ACC [7], _40567_);
  dff (\oc8051_golden_model_1.DPL [0], _43498_);
  dff (\oc8051_golden_model_1.DPL [1], _43499_);
  dff (\oc8051_golden_model_1.DPL [2], _43500_);
  dff (\oc8051_golden_model_1.DPL [3], _43501_);
  dff (\oc8051_golden_model_1.DPL [4], _43502_);
  dff (\oc8051_golden_model_1.DPL [5], _43505_);
  dff (\oc8051_golden_model_1.DPL [6], _43506_);
  dff (\oc8051_golden_model_1.DPL [7], _40568_);
  dff (\oc8051_golden_model_1.DPH [0], _43507_);
  dff (\oc8051_golden_model_1.DPH [1], _43510_);
  dff (\oc8051_golden_model_1.DPH [2], _43511_);
  dff (\oc8051_golden_model_1.DPH [3], _43512_);
  dff (\oc8051_golden_model_1.DPH [4], _43513_);
  dff (\oc8051_golden_model_1.DPH [5], _43514_);
  dff (\oc8051_golden_model_1.DPH [6], _43515_);
  dff (\oc8051_golden_model_1.DPH [7], _40569_);
  dff (\oc8051_golden_model_1.IE [0], _43516_);
  dff (\oc8051_golden_model_1.IE [1], _43517_);
  dff (\oc8051_golden_model_1.IE [2], _43518_);
  dff (\oc8051_golden_model_1.IE [3], _43519_);
  dff (\oc8051_golden_model_1.IE [4], _43520_);
  dff (\oc8051_golden_model_1.IE [5], _43521_);
  dff (\oc8051_golden_model_1.IE [6], _43522_);
  dff (\oc8051_golden_model_1.IE [7], _40571_);
  dff (\oc8051_golden_model_1.IP [0], _43525_);
  dff (\oc8051_golden_model_1.IP [1], _43526_);
  dff (\oc8051_golden_model_1.IP [2], _43527_);
  dff (\oc8051_golden_model_1.IP [3], _43530_);
  dff (\oc8051_golden_model_1.IP [4], _43531_);
  dff (\oc8051_golden_model_1.IP [5], _43532_);
  dff (\oc8051_golden_model_1.IP [6], _43533_);
  dff (\oc8051_golden_model_1.IP [7], _40572_);
  dff (\oc8051_golden_model_1.P0 [0], _43534_);
  dff (\oc8051_golden_model_1.P0 [1], _43535_);
  dff (\oc8051_golden_model_1.P0 [2], _43536_);
  dff (\oc8051_golden_model_1.P0 [3], _43537_);
  dff (\oc8051_golden_model_1.P0 [4], _43538_);
  dff (\oc8051_golden_model_1.P0 [5], _43539_);
  dff (\oc8051_golden_model_1.P0 [6], _43540_);
  dff (\oc8051_golden_model_1.P0 [7], _40573_);
  dff (\oc8051_golden_model_1.P1 [0], _43543_);
  dff (\oc8051_golden_model_1.P1 [1], _43544_);
  dff (\oc8051_golden_model_1.P1 [2], _43545_);
  dff (\oc8051_golden_model_1.P1 [3], _43546_);
  dff (\oc8051_golden_model_1.P1 [4], _43547_);
  dff (\oc8051_golden_model_1.P1 [5], _43550_);
  dff (\oc8051_golden_model_1.P1 [6], _43551_);
  dff (\oc8051_golden_model_1.P1 [7], _40574_);
  dff (\oc8051_golden_model_1.P2 [0], _43552_);
  dff (\oc8051_golden_model_1.P2 [1], _43553_);
  dff (\oc8051_golden_model_1.P2 [2], _43554_);
  dff (\oc8051_golden_model_1.P2 [3], _43555_);
  dff (\oc8051_golden_model_1.P2 [4], _43556_);
  dff (\oc8051_golden_model_1.P2 [5], _43557_);
  dff (\oc8051_golden_model_1.P2 [6], _43558_);
  dff (\oc8051_golden_model_1.P2 [7], _40575_);
  dff (\oc8051_golden_model_1.P3 [0], _43561_);
  dff (\oc8051_golden_model_1.P3 [1], _43562_);
  dff (\oc8051_golden_model_1.P3 [2], _43563_);
  dff (\oc8051_golden_model_1.P3 [3], _43564_);
  dff (\oc8051_golden_model_1.P3 [4], _43565_);
  dff (\oc8051_golden_model_1.P3 [5], _43566_);
  dff (\oc8051_golden_model_1.P3 [6], _43567_);
  dff (\oc8051_golden_model_1.P3 [7], _40577_);
  dff (\oc8051_golden_model_1.PSW [0], _43570_);
  dff (\oc8051_golden_model_1.PSW [1], _43571_);
  dff (\oc8051_golden_model_1.PSW [2], _43572_);
  dff (\oc8051_golden_model_1.PSW [3], _43573_);
  dff (\oc8051_golden_model_1.PSW [4], _43574_);
  dff (\oc8051_golden_model_1.PSW [5], _43575_);
  dff (\oc8051_golden_model_1.PSW [6], _43576_);
  dff (\oc8051_golden_model_1.PSW [7], _40578_);
  dff (\oc8051_golden_model_1.PCON [0], _43579_);
  dff (\oc8051_golden_model_1.PCON [1], _43580_);
  dff (\oc8051_golden_model_1.PCON [2], _43581_);
  dff (\oc8051_golden_model_1.PCON [3], _43582_);
  dff (\oc8051_golden_model_1.PCON [4], _43583_);
  dff (\oc8051_golden_model_1.PCON [5], _43584_);
  dff (\oc8051_golden_model_1.PCON [6], _43585_);
  dff (\oc8051_golden_model_1.PCON [7], _40579_);
  dff (\oc8051_golden_model_1.SBUF [0], _43588_);
  dff (\oc8051_golden_model_1.SBUF [1], _43589_);
  dff (\oc8051_golden_model_1.SBUF [2], _43590_);
  dff (\oc8051_golden_model_1.SBUF [3], _43591_);
  dff (\oc8051_golden_model_1.SBUF [4], _43592_);
  dff (\oc8051_golden_model_1.SBUF [5], _43594_);
  dff (\oc8051_golden_model_1.SBUF [6], _43595_);
  dff (\oc8051_golden_model_1.SBUF [7], _40580_);
  dff (\oc8051_golden_model_1.SCON [0], _43596_);
  dff (\oc8051_golden_model_1.SCON [1], _43599_);
  dff (\oc8051_golden_model_1.SCON [2], _43600_);
  dff (\oc8051_golden_model_1.SCON [3], _43601_);
  dff (\oc8051_golden_model_1.SCON [4], _43602_);
  dff (\oc8051_golden_model_1.SCON [5], _43603_);
  dff (\oc8051_golden_model_1.SCON [6], _43604_);
  dff (\oc8051_golden_model_1.SCON [7], _40581_);
  dff (\oc8051_golden_model_1.SP [0], _43606_);
  dff (\oc8051_golden_model_1.SP [1], _43607_);
  dff (\oc8051_golden_model_1.SP [2], _43608_);
  dff (\oc8051_golden_model_1.SP [3], _43609_);
  dff (\oc8051_golden_model_1.SP [4], _43610_);
  dff (\oc8051_golden_model_1.SP [5], _43611_);
  dff (\oc8051_golden_model_1.SP [6], _43612_);
  dff (\oc8051_golden_model_1.SP [7], _40583_);
  dff (\oc8051_golden_model_1.TCON [0], _43613_);
  dff (\oc8051_golden_model_1.TCON [1], _43614_);
  dff (\oc8051_golden_model_1.TCON [2], _43615_);
  dff (\oc8051_golden_model_1.TCON [3], _43618_);
  dff (\oc8051_golden_model_1.TCON [4], _43619_);
  dff (\oc8051_golden_model_1.TCON [5], _43620_);
  dff (\oc8051_golden_model_1.TCON [6], _43621_);
  dff (\oc8051_golden_model_1.TCON [7], _40584_);
  dff (\oc8051_golden_model_1.TH0 [0], _43624_);
  dff (\oc8051_golden_model_1.TH0 [1], _43625_);
  dff (\oc8051_golden_model_1.TH0 [2], _43626_);
  dff (\oc8051_golden_model_1.TH0 [3], _43627_);
  dff (\oc8051_golden_model_1.TH0 [4], _43628_);
  dff (\oc8051_golden_model_1.TH0 [5], _43629_);
  dff (\oc8051_golden_model_1.TH0 [6], _43630_);
  dff (\oc8051_golden_model_1.TH0 [7], _40585_);
  dff (\oc8051_golden_model_1.TH1 [0], _43631_);
  dff (\oc8051_golden_model_1.TH1 [1], _43632_);
  dff (\oc8051_golden_model_1.TH1 [2], _43633_);
  dff (\oc8051_golden_model_1.TH1 [3], _43634_);
  dff (\oc8051_golden_model_1.TH1 [4], _43635_);
  dff (\oc8051_golden_model_1.TH1 [5], _43638_);
  dff (\oc8051_golden_model_1.TH1 [6], _43639_);
  dff (\oc8051_golden_model_1.TH1 [7], _40586_);
  dff (\oc8051_golden_model_1.TL0 [0], _43640_);
  dff (\oc8051_golden_model_1.TL0 [1], _43643_);
  dff (\oc8051_golden_model_1.TL0 [2], _43644_);
  dff (\oc8051_golden_model_1.TL0 [3], _43645_);
  dff (\oc8051_golden_model_1.TL0 [4], _43646_);
  dff (\oc8051_golden_model_1.TL0 [5], _43647_);
  dff (\oc8051_golden_model_1.TL0 [6], _43648_);
  dff (\oc8051_golden_model_1.TL0 [7], _40587_);
  dff (\oc8051_golden_model_1.TL1 [0], _43649_);
  dff (\oc8051_golden_model_1.TL1 [1], _43650_);
  dff (\oc8051_golden_model_1.TL1 [2], _43651_);
  dff (\oc8051_golden_model_1.TL1 [3], _43652_);
  dff (\oc8051_golden_model_1.TL1 [4], _43653_);
  dff (\oc8051_golden_model_1.TL1 [5], _43654_);
  dff (\oc8051_golden_model_1.TL1 [6], _43655_);
  dff (\oc8051_golden_model_1.TL1 [7], _40589_);
  dff (\oc8051_golden_model_1.TMOD [0], _43658_);
  dff (\oc8051_golden_model_1.TMOD [1], _43659_);
  dff (\oc8051_golden_model_1.TMOD [2], _43660_);
  dff (\oc8051_golden_model_1.TMOD [3], _43663_);
  dff (\oc8051_golden_model_1.TMOD [4], _43664_);
  dff (\oc8051_golden_model_1.TMOD [5], _43665_);
  dff (\oc8051_golden_model_1.TMOD [6], _43666_);
  dff (\oc8051_golden_model_1.TMOD [7], _40590_);
  dff (\oc8051_golden_model_1.PC [0], _43667_);
  dff (\oc8051_golden_model_1.PC [1], _43670_);
  dff (\oc8051_golden_model_1.PC [2], _43671_);
  dff (\oc8051_golden_model_1.PC [3], _43672_);
  dff (\oc8051_golden_model_1.PC [4], _43673_);
  dff (\oc8051_golden_model_1.PC [5], _43674_);
  dff (\oc8051_golden_model_1.PC [6], _43675_);
  dff (\oc8051_golden_model_1.PC [7], _43676_);
  dff (\oc8051_golden_model_1.PC [8], _43677_);
  dff (\oc8051_golden_model_1.PC [9], _43678_);
  dff (\oc8051_golden_model_1.PC [10], _43679_);
  dff (\oc8051_golden_model_1.PC [11], _43682_);
  dff (\oc8051_golden_model_1.PC [12], _43683_);
  dff (\oc8051_golden_model_1.PC [13], _43684_);
  dff (\oc8051_golden_model_1.PC [14], _43685_);
  dff (\oc8051_golden_model_1.PC [15], _40591_);
  dff (\oc8051_golden_model_1.P0INREG [0], _43686_);
  dff (\oc8051_golden_model_1.P0INREG [1], _43687_);
  dff (\oc8051_golden_model_1.P0INREG [2], _43688_);
  dff (\oc8051_golden_model_1.P0INREG [3], _43689_);
  dff (\oc8051_golden_model_1.P0INREG [4], _43690_);
  dff (\oc8051_golden_model_1.P0INREG [5], _43691_);
  dff (\oc8051_golden_model_1.P0INREG [6], _43692_);
  dff (\oc8051_golden_model_1.P0INREG [7], _40592_);
  dff (\oc8051_golden_model_1.P1INREG [0], _43695_);
  dff (\oc8051_golden_model_1.P1INREG [1], _43696_);
  dff (\oc8051_golden_model_1.P1INREG [2], _43697_);
  dff (\oc8051_golden_model_1.P1INREG [3], _43698_);
  dff (\oc8051_golden_model_1.P1INREG [4], _43699_);
  dff (\oc8051_golden_model_1.P1INREG [5], _43702_);
  dff (\oc8051_golden_model_1.P1INREG [6], _43703_);
  dff (\oc8051_golden_model_1.P1INREG [7], _40593_);
  dff (\oc8051_golden_model_1.P2INREG [0], _43704_);
  dff (\oc8051_golden_model_1.P2INREG [1], _43705_);
  dff (\oc8051_golden_model_1.P2INREG [2], _43706_);
  dff (\oc8051_golden_model_1.P2INREG [3], _43707_);
  dff (\oc8051_golden_model_1.P2INREG [4], _43708_);
  dff (\oc8051_golden_model_1.P2INREG [5], _43709_);
  dff (\oc8051_golden_model_1.P2INREG [6], _43710_);
  dff (\oc8051_golden_model_1.P2INREG [7], _40595_);
  dff (\oc8051_golden_model_1.P3INREG [0], _43713_);
  dff (\oc8051_golden_model_1.P3INREG [1], _43714_);
  dff (\oc8051_golden_model_1.P3INREG [2], _43715_);
  dff (\oc8051_golden_model_1.P3INREG [3], _43716_);
  dff (\oc8051_golden_model_1.P3INREG [4], _43717_);
  dff (\oc8051_golden_model_1.P3INREG [5], _43718_);
  dff (\oc8051_golden_model_1.P3INREG [6], _43719_);
  dff (\oc8051_golden_model_1.P3INREG [7], _40596_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03014_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03025_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03046_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03068_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03089_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00893_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03100_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00862_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03111_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03122_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03133_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03144_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03155_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03166_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03177_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00914_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02465_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22434_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02660_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02854_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03057_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03268_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03469_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03670_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03871_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04072_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04173_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04274_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04375_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04476_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04577_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04678_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04779_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24620_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38825_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38826_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38827_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38828_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38829_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38830_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38831_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38811_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38832_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38834_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38835_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38836_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38837_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38838_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38840_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38813_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38841_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38842_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38843_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38844_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38846_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38847_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38848_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38814_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _30468_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06011_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _30471_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _06014_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _30473_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _30475_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _06017_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _30477_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _30479_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _06020_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _30481_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _06023_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _30483_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _30485_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _30487_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _06026_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _30489_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _06029_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _06032_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _06091_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _06093_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _05996_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _06096_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _06099_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _05999_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _06102_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _06002_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _06105_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _06108_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _06111_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _06114_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _06117_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _06120_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _06123_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _06005_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _06008_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39617_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38985_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38986_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38987_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38989_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38990_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38991_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38992_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38993_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38994_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38995_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38996_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38997_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38998_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39000_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39001_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38872_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39005_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39006_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39007_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39008_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39009_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39010_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39011_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39012_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39013_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39014_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39015_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39016_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39017_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39018_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39019_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38874_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39209_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39213_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39216_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39217_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39219_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39222_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39223_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39224_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39226_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39227_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39228_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39230_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38938_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39231_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39232_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39233_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38913_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39237_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39238_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39239_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39240_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39242_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39243_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38914_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39244_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39245_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39246_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39247_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39248_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39249_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39250_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39252_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39253_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39254_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39255_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39256_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39257_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39258_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38918_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39259_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39260_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39261_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39263_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39264_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39265_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39266_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38920_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39267_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39268_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39269_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39270_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39271_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39272_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39274_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39275_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39276_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39277_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39278_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39279_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39280_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39281_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39282_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38922_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39283_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39285_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39286_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39287_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39288_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39289_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39290_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39291_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39292_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39293_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39294_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39296_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39297_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39298_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39299_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38923_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38924_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38927_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38925_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39300_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39301_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39302_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39303_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39304_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39305_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39307_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38928_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39308_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39309_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39310_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39311_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39312_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39313_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39314_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39315_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39316_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38930_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39317_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39318_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39319_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39320_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39321_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39322_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39323_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38931_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _38932_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39324_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39325_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39326_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39328_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39329_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39330_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39331_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38934_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _38935_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39332_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39333_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39334_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38937_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39335_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39336_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39337_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39339_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39340_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39341_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39342_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39343_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39344_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39345_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39346_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39347_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39348_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39350_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39351_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39352_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39353_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39354_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39358_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39359_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39361_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39362_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39363_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39364_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39365_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39366_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39367_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39368_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38939_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39369_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39370_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39372_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39373_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39374_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39375_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39376_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38940_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38942_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39377_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39378_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39379_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39381_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39383_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39384_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39385_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39386_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39387_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39388_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39389_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39390_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39391_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39392_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38944_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38945_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38946_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39394_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39395_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39396_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39397_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39398_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39399_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39400_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39401_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39402_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39403_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39405_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39406_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39407_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39408_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38948_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39764_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39783_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39784_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39785_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39786_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39787_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39788_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39789_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39765_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39766_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39790_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39791_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _43133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _43139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _43145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _43151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _43157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _43163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _43169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _43172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _43413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _43417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _43421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _43425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _43429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _43433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _43437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _43440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _43180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _43184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _43188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _43192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _43196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _43200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _43204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _43207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _43378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _43382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _43386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _43390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _43394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _43398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _43402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _43405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _43346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _43350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _43354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _43358_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _43362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _43366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _43370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _43373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _43315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _43319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _43322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _43326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _43330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _43334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _43338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _43341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _43283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _43287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _43291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _43295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _43299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _43303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _43307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _43310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _43248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _43252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _43256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _43260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _43264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _43268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _43272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _43275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _43215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _43219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _43223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _43227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _43231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _43235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _43239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _43242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _43445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _43449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _43453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _43457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _43461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _43465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _43469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _43472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _43796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _43800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _43804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _43808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _43812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _43816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _43820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _43823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _43764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _43768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _43772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _43776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _43780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _43784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _43788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _43791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _43732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _43736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _43740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _43744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _43748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _43752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _43756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _43759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _43617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _43637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _43657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _43669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _43694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _43712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _43723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _43726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _43477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _43484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _43504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _43524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _43542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _43560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _43578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _43593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _43826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _43829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _43833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _43837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _43841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _43844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _43847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _42875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _01406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _01408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _01410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _01412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _01414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _01416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _01418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _42863_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39648_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39649_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39713_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39714_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39715_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39716_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39717_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39718_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39719_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39650_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24186_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24198_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24210_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24222_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24246_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22313_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08932_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08943_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08965_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08976_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08998_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06695_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13631_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13670_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13679_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13688_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13708_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12723_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _41806_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _42729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _42731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42733_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _42734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _42736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _42738_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41804_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _42742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _41802_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _41800_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _42744_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _42746_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _41798_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _42748_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _42750_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _41796_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _42752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41795_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _42754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _41761_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _41759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _41757_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _41755_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _42756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _42758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _42760_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _41753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _42762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _42764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _42766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _42768_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _42770_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _42772_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _42774_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _41751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _42776_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _42778_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _42780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _42782_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _42784_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _42786_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _42788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _41748_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41207_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41213_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41214_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41216_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41218_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35484_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41220_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41227_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41228_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41230_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35507_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41232_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41235_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41240_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35530_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41244_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41251_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41252_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35552_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21479_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21490_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21502_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21514_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21526_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21538_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09544_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10712_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10723_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10745_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09564_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1264 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1281 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1341 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1382 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1437 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1567 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1603 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1636 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1785 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1802 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1917 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1934 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2066 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2083 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2209 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2450 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2480 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2576 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2694 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2834 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2875 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2892 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0988 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n0988 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n0988 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0988 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0988 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n0988 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n0988 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0989 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0990 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0991 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0992 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0993 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0995 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0996 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1003 , \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1011 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1011 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1011 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1011 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1011 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1011 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1011 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1017 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1018 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1019 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1026 , \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.n1027 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1027 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1027 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1027 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1027 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1043 , \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.n1044 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1044 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1044 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1044 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1044 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1044 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1044 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1137 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1137 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1137 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1137 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1139 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1141 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1141 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1142 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1142 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1142 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1143 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1144 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1144 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1145 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1145 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1146 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1146 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1194 , \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n1239 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1240 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1240 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1240 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1240 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1240 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1240 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1240 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1241 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1241 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1241 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1241 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1241 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1241 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1241 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1241 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1241 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1242 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1242 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1242 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1242 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1242 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1242 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1242 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1242 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1243 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1244 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1244 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1244 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1247 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1247 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1247 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1247 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1247 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1247 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1247 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1247 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1248 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1248 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1248 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1248 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1248 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1248 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1248 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1249 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1251 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1252 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1253 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1254 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1255 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1256 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1264 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1264 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1280 , \oc8051_golden_model_1.n1281 [0]);
  buf(\oc8051_golden_model_1.n1281 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1281 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1281 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1281 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1281 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1281 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1281 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1323 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1323 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1323 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1323 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1323 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1323 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1323 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1323 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1323 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1323 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1323 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1323 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1323 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1323 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1323 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1323 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1325 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1325 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1325 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1325 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1325 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1325 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1325 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1327 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1328 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1329 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1330 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1331 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1332 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1340 , \oc8051_golden_model_1.n1341 [0]);
  buf(\oc8051_golden_model_1.n1341 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1341 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1341 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1341 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1341 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1341 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1343 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1347 [8], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1349 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1349 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1349 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1349 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1350 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1354 [4], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1356 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1356 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1356 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1356 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1356 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1356 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1356 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1356 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1356 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1364 , \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1365 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1365 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1365 [2], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1365 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1365 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1365 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1365 [6], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1365 [7], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1366 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1366 [6], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1381 , \oc8051_golden_model_1.n1382 [0]);
  buf(\oc8051_golden_model_1.n1382 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1382 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1382 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1382 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1404 [8], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1405 , \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1410 [4], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1411 , \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1419 , \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1420 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1420 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1420 [2], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1420 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1420 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1420 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1420 [6], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1420 [7], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1421 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1421 [1], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1421 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1421 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1421 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1421 [5], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1421 [6], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1436 , \oc8051_golden_model_1.n1437 [0]);
  buf(\oc8051_golden_model_1.n1437 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1437 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1437 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1437 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1439 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1439 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1439 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1439 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1439 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1439 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1439 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1439 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1439 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1441 [8], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1442 , \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1443 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1443 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1443 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1443 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1444 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1444 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1444 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1444 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1444 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1446 [4], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1447 , \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1448 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1448 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1448 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1448 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1448 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1448 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1448 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1448 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1448 [8], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1455 , \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1456 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1456 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1456 [2], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1456 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1456 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1456 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1456 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1456 [7], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1457 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1457 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1457 [6], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1472 , \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.n1473 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.n1473 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1473 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1473 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1473 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1473 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1476 [8], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1477 , \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1484 , \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1485 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1485 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1485 [2], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1485 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1485 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1485 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1485 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1485 [7], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1486 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1486 [1], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1486 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1486 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1486 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1486 [5], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1486 [6], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1487 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1487 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1487 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1487 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1489 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1489 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1489 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1489 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1489 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1489 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1489 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1489 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1489 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1491 [8], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1493 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1493 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1495 [4], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1496 , \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1497 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1497 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1497 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1497 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1497 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1497 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1497 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1497 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1497 [8], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1504 , \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1521 , \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1522 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1524 [4], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1525 , \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1526 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1527 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1527 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1527 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1527 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1527 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1527 [5], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1527 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1528 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1528 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1528 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1528 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1528 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1528 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1530 [8], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1531 , \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1538 , \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1539 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1539 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1539 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1539 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1539 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1539 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1539 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1539 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1540 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1540 [1], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1540 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1540 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1540 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1540 [5], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1540 [6], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1541 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1541 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1541 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1541 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1541 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1541 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1541 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1543 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1543 [1], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1543 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1543 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1543 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1543 [5], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1543 [6], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1544 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1544 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1544 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1547 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1547 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1548 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1548 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1548 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1549 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1549 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1549 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1549 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1549 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1549 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1549 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1549 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1550 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1550 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1550 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1550 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1550 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1550 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1550 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1550 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1551 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1551 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1551 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1551 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1551 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1551 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1551 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1552 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1553 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1555 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1557 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1559 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1566 , \oc8051_golden_model_1.n1567 [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1571 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [8], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1575 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1575 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [4], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1585 , \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1586 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1586 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1586 [2], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1586 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1586 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1586 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1586 [6], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1586 [7], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1587 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1602 , \oc8051_golden_model_1.n1603 [0]);
  buf(\oc8051_golden_model_1.n1603 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1603 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1603 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1603 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [8], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1608 , \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1610 [4], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1611 , \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1618 , \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1619 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1619 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1619 [2], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1619 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1619 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1619 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1619 [6], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1619 [7], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1620 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1620 [1], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1620 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1620 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1620 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1620 [5], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1620 [6], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1635 , \oc8051_golden_model_1.n1636 [0]);
  buf(\oc8051_golden_model_1.n1636 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1636 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1636 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1636 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [8], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1641 , \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1643 [4], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1644 , \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1651 , \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1652 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1652 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1652 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1652 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1652 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1652 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1652 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1652 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1653 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1653 [1], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1653 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1653 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1653 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1653 [5], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1653 [6], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1668 , \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.n1669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [8], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1674 , \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1676 [4], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1677 , \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1684 , \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1685 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1685 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1685 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1685 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1685 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1685 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1685 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1685 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1686 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1686 [1], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1686 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1686 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1686 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1686 [5], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1686 [6], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1701 , \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.n1702 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1702 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1702 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1702 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1727 [1], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.n1727 [2], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.n1727 [3], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.n1727 [4], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.n1727 [5], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.n1727 [6], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.n1727 [7], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.n1728 [0], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.n1728 [1], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.n1728 [2], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.n1728 [3], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.n1728 [4], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.n1728 [5], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.n1728 [6], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.n1729 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1784 , \oc8051_golden_model_1.n1785 [0]);
  buf(\oc8051_golden_model_1.n1785 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1785 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1785 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1785 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1785 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1785 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1785 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1801 , \oc8051_golden_model_1.n1802 [0]);
  buf(\oc8051_golden_model_1.n1802 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1802 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1802 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1802 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1802 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1802 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1802 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1818 , \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.n1819 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1819 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1819 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1819 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1819 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1819 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1819 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1835 , \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.n1836 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1836 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1836 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1836 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1836 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1836 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1836 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1859 [1], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.n1859 [2], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.n1859 [3], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.n1859 [4], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.n1859 [5], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.n1859 [6], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.n1859 [7], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.n1860 [0], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.n1860 [1], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.n1860 [2], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.n1860 [3], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.n1860 [4], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.n1860 [5], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.n1860 [6], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.n1861 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1916 , \oc8051_golden_model_1.n1917 [0]);
  buf(\oc8051_golden_model_1.n1917 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1917 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1917 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1917 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1917 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1917 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1917 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1933 , \oc8051_golden_model_1.n1934 [0]);
  buf(\oc8051_golden_model_1.n1934 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1934 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1934 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1934 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1934 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1934 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1934 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1950 , \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.n1951 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1951 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1951 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1951 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1951 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1951 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1951 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1967 , \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.n1968 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1968 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1968 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1968 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1968 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1968 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1968 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2065 , \oc8051_golden_model_1.n2066 [0]);
  buf(\oc8051_golden_model_1.n2066 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2066 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2066 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2066 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2066 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2066 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2066 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2082 , \oc8051_golden_model_1.n2083 [0]);
  buf(\oc8051_golden_model_1.n2083 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2083 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2083 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2083 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2083 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2083 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2083 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2099 , \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.n2100 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2100 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2100 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2100 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2100 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2100 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2116 , \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.n2117 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2117 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2117 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2117 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2117 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2117 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2117 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2121 , \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2122 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2122 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2122 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2122 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2122 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2122 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2122 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2123 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2123 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2123 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2123 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2123 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2123 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2123 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2123 [7], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2124 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2124 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2124 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2124 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2124 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2124 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2124 [6], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2125 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2125 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2125 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2125 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2125 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2125 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2125 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2140 , \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.n2141 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2141 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2141 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2141 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2141 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2141 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2180 , \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2181 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2181 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2181 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2181 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2181 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2181 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2181 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2181 [7], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2182 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2182 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2182 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2182 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2182 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2182 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2182 [6], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2183 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2183 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2183 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2183 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2183 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2183 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2183 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2190 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2190 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2190 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2190 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2191 , \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2192 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2192 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2192 [2], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2192 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2192 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2192 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2192 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2192 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2193 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2193 [1], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2193 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2193 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2193 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2193 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2193 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2208 , \oc8051_golden_model_1.n2209 [0]);
  buf(\oc8051_golden_model_1.n2209 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2209 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2209 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2209 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2209 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2209 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2421 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2424 , \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2426 , \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2432 , \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2433 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2433 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2433 [2], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2433 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2433 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2433 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2433 [6], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2433 [7], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2434 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2434 [1], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2434 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2434 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2434 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2434 [5], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2434 [6], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2449 , \oc8051_golden_model_1.n2450 [0]);
  buf(\oc8051_golden_model_1.n2450 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2450 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2450 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2450 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 , \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2456 , \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2462 , \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2463 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2463 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2463 [2], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2463 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2463 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2463 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2463 [6], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2463 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2464 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2464 [1], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2464 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2464 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2464 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2464 [5], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2464 [6], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2479 , \oc8051_golden_model_1.n2480 [0]);
  buf(\oc8051_golden_model_1.n2480 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2480 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2480 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2480 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 , \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2486 , \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2492 , \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2493 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2493 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2493 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2493 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2494 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2494 [1], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2494 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2494 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2494 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2494 [5], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2494 [6], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2509 , \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.n2510 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2510 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2510 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2510 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 , \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2516 , \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2522 , \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2523 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2523 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2523 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2523 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2523 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2523 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2523 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2523 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2524 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2524 [1], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2524 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2524 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2524 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2524 [5], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2524 [6], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2539 , \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.n2540 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2540 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2540 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2540 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2545 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2545 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2545 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2545 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2545 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2545 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2545 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [7], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n2547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2547 [6], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n2548 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2548 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2548 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2552 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2552 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2552 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2552 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2552 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2552 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2552 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2552 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2552 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2558 , \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2559 [2], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2559 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2559 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2560 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2575 , \oc8051_golden_model_1.n2576 [0]);
  buf(\oc8051_golden_model_1.n2576 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2576 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2576 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2576 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2576 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2576 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2579 , \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [7], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2581 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2581 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2581 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2581 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2581 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2581 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2581 [6], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2582 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2582 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2582 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2582 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2582 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2582 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2582 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2614 , \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2615 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2615 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2615 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2615 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2615 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2615 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2615 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2615 [7], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2616 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2616 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2616 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2616 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2616 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2616 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2616 [6], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2617 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2617 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2617 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2617 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2617 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2617 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2617 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2622 , \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2623 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2623 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2623 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2623 [7], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2624 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2624 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2624 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2624 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2624 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2624 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2624 [6], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2625 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2625 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2625 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2625 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2625 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2625 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2625 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2630 , \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2631 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2631 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2631 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2631 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2631 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2631 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2631 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2631 [7], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2632 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2632 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2632 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2632 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2632 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2632 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2632 [6], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2633 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2633 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2633 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2633 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2633 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2633 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2633 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2638 , \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2639 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2639 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2639 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2640 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2640 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2640 [6], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2641 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2641 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2641 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2641 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2641 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2641 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2641 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2646 , \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2647 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2647 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2647 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2647 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2647 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2647 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2647 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2647 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2648 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2648 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2648 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2648 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2648 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2648 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2648 [6], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2649 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2649 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2649 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2649 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2649 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2649 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2649 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2674 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2674 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2674 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2674 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2674 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2674 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2675 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2675 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2675 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2675 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2675 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2675 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2675 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2676 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2676 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2676 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2676 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2676 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2676 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2676 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2676 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2677 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2677 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2677 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2677 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2678 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2678 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2678 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2678 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2678 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2678 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2678 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2678 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2679 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2680 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2681 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2682 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2683 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2684 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2685 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2686 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2693 , \oc8051_golden_model_1.n2694 [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2715 [0], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2715 [1], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2715 [2], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2715 [3], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2715 [4], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2715 [5], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2715 [6], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2731 [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2731 [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2731 [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2731 [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2731 [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2731 [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2731 [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2732 , \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n2733 , \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n2734 , \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n2735 , \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n2736 , \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n2737 , \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n2738 , \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n2739 , \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n2746 , \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.n2747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2747 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2747 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2747 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2762 , \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.n2763 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2763 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2763 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2763 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2763 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2763 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2763 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2795 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2795 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2795 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2795 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2795 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2795 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2795 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2795 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2796 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2796 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2796 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2796 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2796 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2796 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2796 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2797 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2797 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2797 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2797 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2797 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2797 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2797 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2797 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 , \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2818 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2818 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2818 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2818 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2818 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2818 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2818 [6], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2833 , \oc8051_golden_model_1.n2834 [0]);
  buf(\oc8051_golden_model_1.n2834 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2834 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2834 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2834 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2834 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2834 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2838 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2839 [0], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n2839 [1], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n2839 [2], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n2839 [3], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n2840 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2840 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2840 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2840 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2841 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2842 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2843 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2844 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2855 , \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.n2856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2874 , \oc8051_golden_model_1.n2875 [0]);
  buf(\oc8051_golden_model_1.n2875 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2875 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2875 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2875 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2875 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2875 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2875 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2891 , \oc8051_golden_model_1.n2892 [0]);
  buf(\oc8051_golden_model_1.n2892 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2892 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2892 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2892 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2892 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2892 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2892 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
