
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_jc, ABINPUT, ABINPUT000, ABINPUT000000);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  input [8:0] ABINPUT;
  input [16:0] ABINPUT000;
  input [16:0] ABINPUT000000;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [16:0] \oc8051_top_1.ABINPUT000 ;
  wire [16:0] \oc8051_top_1.ABINPUT000000 ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT000 ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire \oc8051_top_1.oc8051_alu1.divOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.mulOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_jc;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not _13496_ (_05141_, rst);
  not _13497_ (_05142_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  not _13498_ (_05143_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _13499_ (_05144_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05143_);
  and _13500_ (_05145_, _05144_, _05142_);
  and _13501_ (_05146_, _05145_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _13502_ (_05147_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  not _13503_ (_05148_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _13504_ (_05149_, _05145_, _05148_);
  and _13505_ (_05150_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _13506_ (_05151_, _05150_, _05147_);
  not _13507_ (_05152_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  not _13508_ (_05153_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nand _13509_ (_05154_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  or _13510_ (_05155_, _05154_, _05153_);
  and _13511_ (_05156_, _05155_, _05152_);
  and _13512_ (_05157_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05143_);
  and _13513_ (_05158_, _05157_, _05148_);
  and _13514_ (_05159_, _05158_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  or _13515_ (_05160_, _05155_, _05152_);
  nand _13516_ (_05161_, _05160_, _05159_);
  or _13517_ (_05162_, _05161_, _05156_);
  nor _13518_ (_05163_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nor _13519_ (_05164_, _05163_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _13520_ (_05165_, _05164_, _05144_);
  nand _13521_ (_05166_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  not _13522_ (_05167_, _05158_);
  nor _13523_ (_05168_, _05167_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  nand _13524_ (_05169_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and _13525_ (_05170_, _05169_, _05166_);
  and _13526_ (_05171_, _05170_, _05162_);
  and _13527_ (_05172_, _05171_, _05151_);
  not _13528_ (_05173_, _05172_);
  and _13529_ (_05174_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and _13530_ (_05175_, _05174_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _13531_ (_05176_, _05154_, _05153_);
  nor _13532_ (_05177_, _05176_, _05175_);
  and _13533_ (_05178_, _05177_, _05159_);
  and _13534_ (_05179_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _13535_ (_05180_, _05179_, _05178_);
  and _13536_ (_05181_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand _13537_ (_05182_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  nand _13538_ (_05183_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  nand _13539_ (_05184_, _05183_, _05182_);
  nor _13540_ (_05185_, _05184_, _05181_);
  and _13541_ (_05186_, _05185_, _05180_);
  and _13542_ (_05187_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _13543_ (_05188_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _13544_ (_05189_, _05188_, _05187_);
  and _13545_ (_05190_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not _13546_ (_05191_, _05190_);
  not _13547_ (_05192_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _13548_ (_05193_, _05159_, _05192_);
  and _13549_ (_05194_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _13550_ (_05195_, _05194_, _05193_);
  and _13551_ (_05196_, _05195_, _05191_);
  and _13552_ (_05197_, _05196_, _05189_);
  nor _13553_ (_05198_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _13554_ (_05199_, _05198_, _05174_);
  and _13555_ (_05200_, _05199_, _05159_);
  and _13556_ (_05201_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _13557_ (_05202_, _05201_, _05200_);
  and _13558_ (_05203_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand _13559_ (_05204_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nand _13560_ (_05205_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  nand _13561_ (_05206_, _05205_, _05204_);
  nor _13562_ (_05207_, _05206_, _05203_);
  and _13563_ (_05208_, _05207_, _05202_);
  and _13564_ (_05209_, _05208_, _05197_);
  and _13565_ (_05210_, _05209_, _05186_);
  and _13566_ (_05211_, _05210_, _05173_);
  not _13567_ (_05212_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _13568_ (_05213_, _05160_, _05212_);
  and _13569_ (_05214_, _05213_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nand _13570_ (_05215_, _05214_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  or _13571_ (_05216_, _05214_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _13572_ (_05217_, _05216_, _05159_);
  nand _13573_ (_05218_, _05217_, _05215_);
  nand _13574_ (_05219_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _13575_ (_05220_, _05144_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nand _13576_ (_05221_, _05220_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _13577_ (_05222_, _05221_, _05219_);
  nand _13578_ (_05223_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nand _13579_ (_05224_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _13580_ (_05225_, _05224_, _05223_);
  and _13581_ (_05226_, _05225_, _05222_);
  and _13582_ (_05227_, _05226_, _05218_);
  not _13583_ (_05228_, _05227_);
  nand _13584_ (_05229_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or _13585_ (_05230_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand _13586_ (_05231_, _05230_, _05229_);
  nand _13587_ (_05232_, _05231_, _05159_);
  nand _13588_ (_05233_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _13589_ (_05234_, _05233_, _05221_);
  nand _13590_ (_05236_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nand _13591_ (_05237_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _13592_ (_05239_, _05237_, _05236_);
  and _13593_ (_05240_, _05239_, _05234_);
  nand _13594_ (_05241_, _05240_, _05232_);
  nor _13595_ (_05242_, _05241_, _05228_);
  not _13596_ (_05243_, _05159_);
  and _13597_ (_05244_, _05160_, _05212_);
  or _13598_ (_05245_, _05244_, _05243_);
  or _13599_ (_05246_, _05245_, _05213_);
  nand _13600_ (_05247_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _13601_ (_05248_, _05247_, _05221_);
  nand _13602_ (_05249_, _05165_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nand _13603_ (_05250_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  and _13604_ (_05252_, _05250_, _05249_);
  nand _13605_ (_05253_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _13606_ (_05254_, _05253_, _05252_);
  and _13607_ (_05255_, _05254_, _05248_);
  and _13608_ (_05256_, _05255_, _05246_);
  or _13609_ (_05257_, _05213_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _13610_ (_05258_, _05214_, _05243_);
  nand _13611_ (_05259_, _05258_, _05257_);
  nand _13612_ (_05260_, _05149_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _13613_ (_05261_, _05260_, _05221_);
  nand _13614_ (_05262_, _05168_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  nand _13615_ (_05263_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _13616_ (_05264_, _05263_, _05262_);
  and _13617_ (_05265_, _05264_, _05261_);
  and _13618_ (_05266_, _05265_, _05259_);
  and _13619_ (_05267_, _05266_, _05256_);
  and _13620_ (_05268_, _05267_, _05242_);
  and _13621_ (_05269_, _05268_, _05211_);
  not _13622_ (_05270_, _05269_);
  and _13623_ (_05271_, _05186_, _05172_);
  and _13624_ (_05272_, _05209_, _05271_);
  and _13625_ (_05273_, _05272_, _05268_);
  not _13626_ (_05274_, _05208_);
  nor _13627_ (_05275_, _05274_, _05197_);
  and _13628_ (_05276_, _05271_, _05275_);
  and _13629_ (_05277_, _05268_, _05276_);
  nor _13630_ (_05278_, _05277_, _05273_);
  and _13631_ (_05279_, _05278_, _05270_);
  not _13632_ (_05280_, _05266_);
  nor _13633_ (_05281_, _05280_, _05256_);
  and _13634_ (_05282_, _05281_, _05242_);
  and _13635_ (_05283_, _05282_, _05276_);
  and _13636_ (_05284_, _05211_, _05282_);
  nor _13637_ (_05285_, _05284_, _05283_);
  not _13638_ (_05286_, _05197_);
  and _13639_ (_05287_, _05186_, _05208_);
  and _13640_ (_05288_, _05287_, _05286_);
  and _13641_ (_05289_, _05288_, _05173_);
  and _13642_ (_05290_, _05289_, _05268_);
  and _13643_ (_05291_, _05272_, _05282_);
  nor _13644_ (_05292_, _05291_, _05290_);
  and _13645_ (_05293_, _05292_, _05285_);
  and _13646_ (_05294_, _05293_, _05279_);
  not _13647_ (_05295_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _13648_ (_05296_, _05143_, \oc8051_top_1.oc8051_decoder1.wr );
  and _13649_ (_05297_, _05296_, _05295_);
  nand _13650_ (_05298_, _05297_, _05279_);
  or _13651_ (_05299_, _05298_, _05294_);
  and _13652_ (_05300_, _05299_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  not _13653_ (_05301_, _05290_);
  nor _13654_ (_05302_, _05291_, _05283_);
  nand _13655_ (_05303_, _05302_, _05301_);
  and _13656_ (_05305_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _13657_ (_05306_, _05305_, _05303_);
  not _13658_ (_05307_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  not _13659_ (_05308_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or _13660_ (_05309_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _13661_ (_05310_, _05309_, _05308_);
  nor _13662_ (_05311_, _05310_, _05307_);
  not _13663_ (_05312_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nand _13664_ (_05313_, _05308_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _13665_ (_05314_, _05313_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor _13666_ (_05315_, _05314_, _05312_);
  nor _13667_ (_05316_, _05315_, _05311_);
  not _13668_ (_05317_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _13669_ (_05318_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _13670_ (_05319_, _05318_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor _13671_ (_05320_, _05319_, _05317_);
  not _13672_ (_05321_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _13673_ (_05322_, _05313_, _05321_);
  not _13674_ (_05323_, _05322_);
  and _13675_ (_05324_, _05323_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _13676_ (_05325_, _05324_, _05320_);
  and _13677_ (_05326_, _05325_, _05316_);
  nor _13678_ (_05327_, _05309_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  not _13679_ (_05328_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _13680_ (_05330_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05328_);
  nor _13681_ (_05331_, _05330_, ABINPUT[5]);
  nand _13682_ (_05332_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05328_);
  nor _13683_ (_05333_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor _13684_ (_05334_, _05333_, _05331_);
  and _13685_ (_05335_, _05334_, _05327_);
  and _13686_ (_05336_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _13687_ (_05337_, _05336_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _13688_ (_05338_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  not _13689_ (_05339_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _13690_ (_05341_, _05336_, _05321_);
  nor _13691_ (_05342_, _05341_, _05339_);
  nor _13692_ (_05343_, _05342_, _05338_);
  not _13693_ (_05344_, _05343_);
  nor _13694_ (_05345_, _05344_, _05335_);
  and _13695_ (_05346_, _05345_, _05326_);
  and _13696_ (_05347_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05143_);
  and _13697_ (_05348_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05143_);
  nor _13698_ (_05349_, _05348_, _05347_);
  not _13699_ (_05350_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or _13700_ (_05351_, _05350_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _13701_ (_05352_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _05143_);
  not _13702_ (_05353_, _05352_);
  and _13703_ (_05354_, _05353_, _05351_);
  and _13704_ (_05355_, _05354_, _05349_);
  not _13705_ (_05356_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _13706_ (_05357_, _05347_, _05356_);
  nand _13707_ (_05358_, _05357_, _05350_);
  nand _13708_ (_05359_, _05349_, _05352_);
  nand _13709_ (_05360_, _05359_, _05358_);
  nor _13710_ (_05361_, _05360_, _05355_);
  and _13711_ (_05362_, _05348_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _13712_ (_05363_, _05362_, _05350_);
  not _13713_ (_05364_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _13714_ (_05365_, _05348_, _05364_);
  not _13715_ (_05366_, _05365_);
  nor _13716_ (_05367_, _05366_, _05351_);
  nor _13717_ (_05368_, _05367_, _05363_);
  and _13718_ (_05370_, _05368_, _05361_);
  nor _13719_ (_05371_, _05370_, _05346_);
  not _13720_ (_05372_, _05371_);
  not _13721_ (_05373_, _05346_);
  and _13722_ (_05374_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _13723_ (_05375_, _05374_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _13724_ (_05376_, _05375_);
  or _13725_ (_05377_, _05330_, ABINPUT[0]);
  or _13726_ (_05378_, _05332_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _13727_ (_05379_, _05378_, _05377_);
  or _13728_ (_05380_, _05379_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and _13729_ (_05381_, _05380_, _05376_);
  not _13730_ (_05382_, _05381_);
  not _13731_ (_05383_, _05310_);
  and _13732_ (_05384_, _05383_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  not _13733_ (_05385_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _13734_ (_05386_, _05314_, _05385_);
  nor _13735_ (_05387_, _05386_, _05384_);
  not _13736_ (_05388_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _13737_ (_05389_, _05322_, _05388_);
  not _13738_ (_05390_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _13739_ (_05391_, _05319_, _05390_);
  nor _13740_ (_05392_, _05391_, _05389_);
  and _13741_ (_05393_, _05392_, _05387_);
  not _13742_ (_05394_, _05327_);
  or _13743_ (_05395_, _05330_, ABINPUT[4]);
  or _13744_ (_05396_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _13745_ (_05397_, _05396_, _05395_);
  or _13746_ (_05398_, _05397_, _05394_);
  not _13747_ (_05399_, _05341_);
  and _13748_ (_05400_, _05399_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _13749_ (_05401_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor _13750_ (_05402_, _05401_, _05400_);
  and _13751_ (_05403_, _05402_, _05398_);
  and _13752_ (_05404_, _05403_, _05393_);
  not _13753_ (_05405_, _05404_);
  not _13754_ (_05406_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or _13755_ (_05407_, _05314_, _05406_);
  not _13756_ (_05408_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  or _13757_ (_05409_, _05310_, _05408_);
  and _13758_ (_05410_, _05409_, _05407_);
  not _13759_ (_05411_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _13760_ (_05412_, _05319_, _05411_);
  nand _13761_ (_05413_, _05323_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _13762_ (_05414_, _05413_, _05412_);
  and _13763_ (_05415_, _05414_, _05410_);
  or _13764_ (_05416_, _05330_, ABINPUT[1]);
  or _13765_ (_05417_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _13766_ (_05418_, _05417_, _05416_);
  or _13767_ (_05419_, _05418_, _05394_);
  not _13768_ (_05420_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _13769_ (_05421_, _05341_, _05420_);
  nand _13770_ (_05422_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and _13771_ (_05423_, _05422_, _05421_);
  and _13772_ (_05424_, _05423_, _05419_);
  and _13773_ (_05425_, _05424_, _05415_);
  or _13774_ (_05426_, _05330_, ABINPUT[2]);
  or _13775_ (_05427_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _13776_ (_05428_, _05427_, _05426_);
  or _13777_ (_05429_, _05428_, _05394_);
  not _13778_ (_05430_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or _13779_ (_05431_, _05314_, _05430_);
  not _13780_ (_05432_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or _13781_ (_05433_, _05310_, _05432_);
  and _13782_ (_05434_, _05433_, _05431_);
  and _13783_ (_05435_, _05434_, _05429_);
  not _13784_ (_05436_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _13785_ (_05437_, _05319_, _05436_);
  not _13786_ (_05438_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _13787_ (_05439_, _05322_, _05438_);
  and _13788_ (_05440_, _05439_, _05437_);
  not _13789_ (_05441_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _13790_ (_05442_, _05341_, _05441_);
  nand _13791_ (_05443_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _13792_ (_05444_, _05443_, _05442_);
  and _13793_ (_05445_, _05444_, _05440_);
  and _13794_ (_05446_, _05445_, _05435_);
  not _13795_ (_05447_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _13796_ (_05448_, _05314_, _05447_);
  not _13797_ (_05449_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or _13798_ (_05450_, _05310_, _05449_);
  and _13799_ (_05452_, _05450_, _05448_);
  not _13800_ (_05453_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _13801_ (_05454_, _05322_, _05453_);
  not _13802_ (_05455_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _13803_ (_05456_, _05319_, _05455_);
  and _13804_ (_05457_, _05456_, _05454_);
  and _13805_ (_05458_, _05457_, _05452_);
  or _13806_ (_05459_, _05330_, ABINPUT[3]);
  or _13807_ (_05460_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _13808_ (_05461_, _05460_, _05459_);
  or _13809_ (_05462_, _05461_, _05394_);
  nand _13810_ (_05463_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not _13811_ (_05464_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _13812_ (_05465_, _05341_, _05464_);
  and _13813_ (_05466_, _05465_, _05463_);
  and _13814_ (_05467_, _05466_, _05462_);
  and _13815_ (_05469_, _05467_, _05458_);
  and _13816_ (_05470_, _05469_, _05446_);
  nand _13817_ (_05471_, _05470_, _05425_);
  or _13818_ (_05472_, _05471_, _05405_);
  or _13819_ (_05473_, _05472_, _05382_);
  or _13820_ (_05474_, _05446_, _05425_);
  nor _13821_ (_05475_, _05474_, _05469_);
  nand _13822_ (_05476_, _05475_, _05405_);
  or _13823_ (_05477_, _05476_, _05381_);
  nand _13824_ (_05478_, _05477_, _05473_);
  nand _13825_ (_05479_, _05478_, _05373_);
  nor _13826_ (_05480_, _05351_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _13827_ (_05481_, _05362_, _05480_);
  or _13828_ (_05482_, _05478_, _05373_);
  and _13829_ (_05483_, _05482_, _05481_);
  nand _13830_ (_05484_, _05483_, _05479_);
  and _13831_ (_05485_, _05365_, _05354_);
  nor _13832_ (_05486_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _13833_ (_05487_, _05486_, _05334_);
  not _13834_ (_05488_, _05487_);
  and _13835_ (_05489_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _13836_ (_05490_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not _13837_ (_05491_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _13838_ (_05492_, _05491_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _13839_ (_05493_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _13840_ (_05494_, _05493_, _05490_);
  and _13841_ (_05495_, _05494_, _05488_);
  nor _13842_ (_05496_, _05495_, _05346_);
  and _13843_ (_05497_, _05495_, _05346_);
  nor _13844_ (_05498_, _05497_, _05496_);
  nand _13845_ (_05499_, _05498_, _05485_);
  and _13846_ (_05500_, _05352_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _13847_ (_05501_, _05500_, _05357_);
  and _13848_ (_05503_, _05501_, _05496_);
  and _13849_ (_05504_, _05480_, _05357_);
  and _13850_ (_05505_, _05504_, _05346_);
  nor _13851_ (_05506_, _05505_, _05503_);
  and _13852_ (_05507_, _05382_, _05346_);
  not _13853_ (_05508_, _05507_);
  and _13854_ (_05509_, _05362_, _05500_);
  not _13855_ (_05510_, _05509_);
  and _13856_ (_05511_, _05495_, _05381_);
  nor _13857_ (_05512_, _05511_, _05510_);
  and _13858_ (_05513_, _05512_, _05508_);
  and _13859_ (_05514_, _05352_, _05350_);
  and _13860_ (_05515_, _05365_, _05514_);
  not _13861_ (_05516_, _05515_);
  nor _13862_ (_05517_, _05516_, _05497_);
  nor _13863_ (_05518_, _05517_, _05513_);
  and _13864_ (_05519_, _05518_, _05506_);
  and _13865_ (_05520_, _05519_, _05499_);
  and _13866_ (_05521_, _05520_, _05484_);
  nand _13867_ (_05522_, _05521_, _05372_);
  and _13868_ (_05523_, _05297_, _05284_);
  and _13869_ (_05524_, _05523_, _05522_);
  or _13870_ (_05525_, _05524_, _05306_);
  or _13871_ (_05526_, _05525_, _05300_);
  and _13872_ (_09109_, _05526_, _05141_);
  not _13873_ (_05527_, _05486_);
  or _13874_ (_05528_, _05527_, _05461_);
  and _13875_ (_05529_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and _13876_ (_05530_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _13877_ (_05531_, _05530_, _05529_);
  and _13878_ (_05532_, _05531_, _05528_);
  nor _13879_ (_05533_, _05532_, _05510_);
  not _13880_ (_05534_, _05469_);
  nand _13881_ (_05535_, _05424_, _05415_);
  and _13882_ (_05536_, _05535_, _05381_);
  nand _13883_ (_05537_, _05445_, _05435_);
  or _13884_ (_05538_, _05537_, _05382_);
  and _13885_ (_05539_, _05538_, _05474_);
  nor _13886_ (_05540_, _05539_, _05536_);
  nand _13887_ (_05541_, _05540_, _05534_);
  or _13888_ (_05542_, _05540_, _05534_);
  and _13889_ (_05543_, _05542_, _05481_);
  and _13890_ (_05544_, _05543_, _05541_);
  nor _13891_ (_05545_, _05544_, _05533_);
  nor _13892_ (_05546_, _05469_, _05370_);
  not _13893_ (_05547_, _05546_);
  nor _13894_ (_05548_, _05532_, _05469_);
  and _13895_ (_05549_, _05548_, _05501_);
  and _13896_ (_05550_, _05504_, _05469_);
  nor _13897_ (_05551_, _05550_, _05549_);
  and _13898_ (_05552_, _05532_, _05469_);
  nor _13899_ (_05553_, _05552_, _05548_);
  and _13900_ (_05554_, _05553_, _05485_);
  nor _13901_ (_05555_, _05552_, _05516_);
  nor _13902_ (_05556_, _05555_, _05554_);
  and _13903_ (_05557_, _05556_, _05551_);
  and _13904_ (_05559_, _05557_, _05547_);
  and _13905_ (_05560_, _05559_, _05545_);
  not _13906_ (_05561_, _05560_);
  and _13907_ (_05562_, _05561_, _05284_);
  or _13908_ (_05563_, _05303_, _05299_);
  and _13909_ (_05564_, _05563_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or _13910_ (_05565_, _05564_, _05562_);
  or _13911_ (_05566_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _13912_ (_05567_, _05566_, _05141_);
  and _13913_ (_10437_, _05567_, _05565_);
  not _13914_ (_05568_, _05291_);
  nand _13915_ (_05569_, _05568_, _05285_);
  and _13916_ (_05570_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _13917_ (_05571_, _05570_, _05569_);
  not _13918_ (_05572_, _05297_);
  nand _13919_ (_05573_, _05282_, _05287_);
  or _13920_ (_05574_, _05573_, _05572_);
  and _13921_ (_05575_, _05574_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _13922_ (_05576_, _05289_, _05282_);
  or _13923_ (_05577_, _05527_, _05418_);
  nand _13924_ (_05578_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nand _13925_ (_05579_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _13926_ (_05580_, _05579_, _05578_);
  and _13927_ (_05581_, _05580_, _05577_);
  and _13928_ (_05582_, _05581_, _05425_);
  not _13929_ (_05583_, _05485_);
  not _13930_ (_05584_, _05581_);
  and _13931_ (_05585_, _05584_, _05535_);
  or _13932_ (_05586_, _05585_, _05583_);
  and _13933_ (_05587_, _05586_, _05516_);
  or _13934_ (_05588_, _05587_, _05582_);
  not _13935_ (_05589_, _05501_);
  or _13936_ (_05590_, _05581_, _05425_);
  or _13937_ (_05591_, _05590_, _05589_);
  not _13938_ (_05592_, _05504_);
  or _13939_ (_05593_, _05592_, _05535_);
  and _13940_ (_05594_, _05593_, _05591_);
  or _13941_ (_05595_, _05581_, _05510_);
  not _13942_ (_05597_, _05481_);
  or _13943_ (_05598_, _05597_, _05535_);
  and _13944_ (_05600_, _05598_, _05595_);
  or _13945_ (_05601_, _05425_, _05370_);
  and _13946_ (_05602_, _05601_, _05600_);
  and _13947_ (_05603_, _05602_, _05594_);
  and _13948_ (_05604_, _05603_, _05588_);
  nor _13949_ (_05605_, _05604_, _05572_);
  and _13950_ (_05606_, _05605_, _05576_);
  or _13951_ (_05607_, _05606_, _05575_);
  or _13952_ (_05608_, _05607_, _05571_);
  and _13953_ (_00002_, _05608_, _05141_);
  and _13954_ (_05609_, _05292_, _05270_);
  not _13955_ (_05610_, _05609_);
  nand _13956_ (_05611_, _05268_, _05287_);
  and _13957_ (_05612_, _05611_, _05302_);
  nand _13958_ (_05613_, _05297_, _05278_);
  or _13959_ (_05614_, _05613_, _05612_);
  or _13960_ (_05615_, _05614_, _05610_);
  and _13961_ (_05616_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _13962_ (_05617_, _05297_, _05283_);
  and _13963_ (_05618_, _05617_, _05522_);
  or _13964_ (_05619_, _05618_, _05616_);
  and _13965_ (_02660_, _05619_, _05141_);
  and _13966_ (_05620_, _05605_, _05290_);
  not _13967_ (_05621_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _13968_ (_05622_, _05297_, _05290_);
  nor _13969_ (_05623_, _05622_, _05621_);
  or _13970_ (_05624_, _05623_, _05620_);
  and _13971_ (_06673_, _05624_, _05141_);
  nor _13972_ (_05625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _13973_ (_05626_, _05625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not _13974_ (_05627_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _13975_ (_05628_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _13976_ (_05629_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _13977_ (_05630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _13978_ (_05631_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _05630_);
  nor _13979_ (_05632_, _05631_, _05629_);
  nor _13980_ (_05633_, _05632_, _05628_);
  nor _13981_ (_05634_, _05633_, _05627_);
  and _13982_ (_05635_, _05630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _13983_ (_05636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or _13984_ (_05637_, _05636_, _05635_);
  and _13985_ (_05638_, _05637_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _13986_ (_05639_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _13987_ (_05640_, _05630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor _13988_ (_05641_, _05640_, _05639_);
  and _13989_ (_05642_, _05641_, _05638_);
  nand _13990_ (_05643_, _05642_, _05634_);
  and _13991_ (_05644_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor _13992_ (_05645_, _05644_, _05626_);
  and _13993_ (_05646_, _05296_, _05167_);
  and _13994_ (_05647_, _05646_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _13995_ (_05648_, _05241_, _05227_);
  and _13996_ (_05649_, _05648_, _05267_);
  nor _13997_ (_05650_, _05208_, _05197_);
  nor _13998_ (_05651_, _05186_, _05172_);
  and _13999_ (_05652_, _05651_, _05650_);
  and _14000_ (_05653_, _05652_, _05649_);
  and _14001_ (_05654_, _05653_, _05647_);
  or _14002_ (_05655_, _05654_, _05645_);
  and _14003_ (_05656_, _05480_, _05349_);
  not _14004_ (_05657_, _05656_);
  not _14005_ (_05658_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _14006_ (_05659_, _05310_, _05658_);
  not _14007_ (_05660_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _14008_ (_05661_, _05314_, _05660_);
  nor _14009_ (_05662_, _05661_, _05659_);
  not _14010_ (_05663_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _14011_ (_05664_, _05319_, _05663_);
  not _14012_ (_05665_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _14013_ (_05666_, _05322_, _05665_);
  nor _14014_ (_05667_, _05666_, _05664_);
  and _14015_ (_05668_, _05667_, _05662_);
  nor _14016_ (_05669_, _05330_, ABINPUT[8]);
  nor _14017_ (_05670_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor _14018_ (_05671_, _05670_, _05669_);
  and _14019_ (_05672_, _05671_, _05327_);
  not _14020_ (_05673_, _05672_);
  and _14021_ (_05674_, _05399_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _14022_ (_05675_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _14023_ (_05676_, _05675_, _05674_);
  and _14024_ (_05677_, _05676_, _05673_);
  and _14025_ (_05678_, _05677_, _05668_);
  and _14026_ (_05679_, _05671_, _05486_);
  not _14027_ (_05680_, _05679_);
  and _14028_ (_05681_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _14029_ (_05682_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _14030_ (_05683_, _05682_, _05681_);
  and _14031_ (_05684_, _05683_, _05680_);
  not _14032_ (_05685_, _05684_);
  and _14033_ (_05686_, _05685_, _05678_);
  nor _14034_ (_05688_, _05684_, _05678_);
  and _14035_ (_05689_, _05684_, _05678_);
  nor _14036_ (_05691_, _05689_, _05688_);
  not _14037_ (_05692_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _14038_ (_05693_, _05314_, _05692_);
  not _14039_ (_05694_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor _14040_ (_05695_, _05310_, _05694_);
  nor _14041_ (_05696_, _05695_, _05693_);
  and _14042_ (_05697_, _05323_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _14043_ (_05699_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _14044_ (_05700_, _05319_, _05699_);
  nor _14045_ (_05701_, _05700_, _05697_);
  and _14046_ (_05702_, _05701_, _05696_);
  nor _14047_ (_05703_, _05330_, ABINPUT[7]);
  nor _14048_ (_05704_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor _14049_ (_05705_, _05704_, _05703_);
  and _14050_ (_05706_, _05705_, _05327_);
  not _14051_ (_05708_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _14052_ (_05709_, _05341_, _05708_);
  and _14053_ (_05710_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor _14054_ (_05711_, _05710_, _05709_);
  not _14055_ (_05712_, _05711_);
  nor _14056_ (_05713_, _05712_, _05706_);
  and _14057_ (_05715_, _05713_, _05702_);
  not _14058_ (_05716_, _05715_);
  and _14059_ (_05718_, _05705_, _05486_);
  not _14060_ (_05719_, _05718_);
  and _14061_ (_05721_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _14062_ (_05722_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _14063_ (_05723_, _05722_, _05721_);
  and _14064_ (_05724_, _05723_, _05719_);
  and _14065_ (_05725_, _05724_, _05716_);
  nor _14066_ (_05727_, _05724_, _05715_);
  and _14067_ (_05728_, _05724_, _05715_);
  nor _14068_ (_05730_, _05728_, _05727_);
  not _14069_ (_05731_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _14070_ (_05733_, _05314_, _05731_);
  not _14071_ (_05734_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor _14072_ (_05736_, _05310_, _05734_);
  nor _14073_ (_05737_, _05736_, _05733_);
  not _14074_ (_05739_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _14075_ (_05740_, _05319_, _05739_);
  not _14076_ (_05742_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _14077_ (_05743_, _05322_, _05742_);
  nor _14078_ (_05745_, _05743_, _05740_);
  and _14079_ (_05746_, _05745_, _05737_);
  nor _14080_ (_05747_, _05330_, ABINPUT[6]);
  nor _14081_ (_05748_, _05332_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor _14082_ (_05749_, _05748_, _05747_);
  and _14083_ (_05750_, _05749_, _05327_);
  not _14084_ (_05751_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _14085_ (_05752_, _05341_, _05751_);
  and _14086_ (_05753_, _05337_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nor _14087_ (_05754_, _05753_, _05752_);
  not _14088_ (_05755_, _05754_);
  nor _14089_ (_05757_, _05755_, _05750_);
  and _14090_ (_05758_, _05757_, _05746_);
  not _14091_ (_05759_, _05758_);
  and _14092_ (_05761_, _05749_, _05486_);
  not _14093_ (_05762_, _05761_);
  and _14094_ (_05763_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _14095_ (_05765_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _14096_ (_05766_, _05765_, _05763_);
  and _14097_ (_05768_, _05766_, _05762_);
  and _14098_ (_05769_, _05768_, _05759_);
  not _14099_ (_05771_, _05495_);
  and _14100_ (_05772_, _05771_, _05346_);
  nor _14101_ (_05773_, _05768_, _05758_);
  and _14102_ (_05774_, _05768_, _05758_);
  nor _14103_ (_05775_, _05774_, _05773_);
  nor _14104_ (_05776_, _05775_, _05772_);
  nor _14105_ (_05777_, _05776_, _05769_);
  nor _14106_ (_05778_, _05777_, _05730_);
  nor _14107_ (_05779_, _05778_, _05725_);
  and _14108_ (_05781_, _05777_, _05730_);
  nor _14109_ (_05782_, _05781_, _05778_);
  and _14110_ (_05784_, _05775_, _05772_);
  nor _14111_ (_05785_, _05784_, _05776_);
  not _14112_ (_05786_, _05785_);
  not _14113_ (_05787_, _05498_);
  nor _14114_ (_05788_, _05527_, _05397_);
  not _14115_ (_05789_, _05788_);
  and _14116_ (_05791_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _14117_ (_05792_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _14118_ (_05794_, _05792_, _05791_);
  and _14119_ (_05795_, _05794_, _05789_);
  nor _14120_ (_05796_, _05795_, _05404_);
  and _14121_ (_05797_, _05795_, _05404_);
  nor _14122_ (_05798_, _05797_, _05796_);
  not _14123_ (_05799_, _05532_);
  nor _14124_ (_05800_, _05799_, _05469_);
  not _14125_ (_05801_, _05553_);
  and _14126_ (_05802_, _05584_, _05425_);
  or _14127_ (_05803_, _05527_, _05428_);
  nand _14128_ (_05804_, _05489_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand _14129_ (_05805_, _05492_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _14130_ (_05806_, _05805_, _05804_);
  and _14131_ (_05807_, _05806_, _05803_);
  and _14132_ (_05808_, _05807_, _05446_);
  nand _14133_ (_05809_, _05806_, _05803_);
  and _14134_ (_05810_, _05809_, _05537_);
  nor _14135_ (_05811_, _05810_, _05808_);
  or _14136_ (_05812_, _05811_, _05802_);
  or _14137_ (_05813_, _05809_, _05446_);
  nand _14138_ (_05814_, _05813_, _05812_);
  and _14139_ (_05815_, _05814_, _05801_);
  nor _14140_ (_05816_, _05815_, _05800_);
  nor _14141_ (_05817_, _05816_, _05798_);
  and _14142_ (_05818_, _05816_, _05798_);
  or _14143_ (_05819_, _05818_, _05817_);
  nor _14144_ (_05820_, _05814_, _05801_);
  or _14145_ (_05821_, _05820_, _05815_);
  and _14146_ (_05822_, _05811_, _05802_);
  not _14147_ (_05823_, _05822_);
  nand _14148_ (_05824_, _05823_, _05812_);
  nor _14149_ (_05825_, _05585_, _05582_);
  nor _14150_ (_05826_, _05825_, _05382_);
  and _14151_ (_05827_, _05826_, _05824_);
  and _14152_ (_05828_, _05827_, _05821_);
  and _14153_ (_05829_, _05828_, _05819_);
  not _14154_ (_05830_, _05795_);
  or _14155_ (_05831_, _05830_, _05404_);
  and _14156_ (_05832_, _05830_, _05404_);
  or _14157_ (_05833_, _05816_, _05832_);
  and _14158_ (_05834_, _05833_, _05831_);
  or _14159_ (_05835_, _05834_, _05829_);
  and _14160_ (_05836_, _05835_, _05787_);
  and _14161_ (_05837_, _05836_, _05786_);
  not _14162_ (_05838_, _05837_);
  nor _14163_ (_05839_, _05838_, _05782_);
  nor _14164_ (_05840_, _05839_, _05779_);
  nor _14165_ (_05841_, _05840_, _05691_);
  nor _14166_ (_05842_, _05841_, _05686_);
  or _14167_ (_05843_, _05842_, _05657_);
  and _14168_ (_05844_, _05514_, _05349_);
  not _14169_ (_05845_, _05844_);
  not _14170_ (_05846_, _05688_);
  not _14171_ (_05847_, _05548_);
  and _14172_ (_05848_, _05811_, _05585_);
  or _14173_ (_05849_, _05848_, _05810_);
  nand _14174_ (_05850_, _05849_, _05553_);
  nand _14175_ (_05851_, _05850_, _05847_);
  or _14176_ (_05852_, _05851_, _05798_);
  nand _14177_ (_05853_, _05851_, _05798_);
  and _14178_ (_05854_, _05853_, _05852_);
  and _14179_ (_05855_, _05825_, _05381_);
  and _14180_ (_05856_, _05855_, _05811_);
  or _14181_ (_05857_, _05849_, _05553_);
  and _14182_ (_05858_, _05857_, _05850_);
  and _14183_ (_05859_, _05858_, _05856_);
  and _14184_ (_05860_, _05859_, _05854_);
  not _14185_ (_05861_, _05797_);
  and _14186_ (_05862_, _05851_, _05861_);
  or _14187_ (_05863_, _05862_, _05796_);
  or _14188_ (_05864_, _05863_, _05860_);
  nand _14189_ (_05865_, _05864_, _05498_);
  and _14190_ (_05866_, _05775_, _05496_);
  nor _14191_ (_05867_, _05775_, _05496_);
  nor _14192_ (_05868_, _05867_, _05866_);
  not _14193_ (_05869_, _05868_);
  or _14194_ (_05870_, _05869_, _05865_);
  not _14195_ (_05871_, _05730_);
  nor _14196_ (_05872_, _05866_, _05773_);
  nor _14197_ (_05873_, _05872_, _05871_);
  and _14198_ (_05874_, _05872_, _05871_);
  nor _14199_ (_05875_, _05874_, _05873_);
  not _14200_ (_05876_, _05875_);
  or _14201_ (_05877_, _05876_, _05870_);
  nor _14202_ (_05878_, _05873_, _05727_);
  and _14203_ (_05879_, _05878_, _05877_);
  or _14204_ (_05880_, _05879_, _05689_);
  and _14205_ (_05881_, _05880_, _05846_);
  or _14206_ (_05882_, _05881_, _05845_);
  and _14207_ (_05883_, _05514_, _05357_);
  and _14208_ (_05884_, _05758_, _05715_);
  nor _14209_ (_05885_, _05884_, _05678_);
  and _14210_ (_05886_, _05885_, _05382_);
  nor _14211_ (_05887_, _05470_, _05404_);
  nor _14212_ (_05888_, _05885_, _05382_);
  or _14213_ (_05889_, _05888_, _05887_);
  or _14214_ (_05890_, _05889_, _05886_);
  and _14215_ (_05891_, _05890_, _05883_);
  and _14216_ (_05892_, _05365_, _05500_);
  not _14217_ (_05893_, _05892_);
  nor _14218_ (_05894_, _05678_, _05893_);
  and _14219_ (_05895_, _05379_, _05375_);
  and _14220_ (_05896_, _05365_, _05480_);
  and _14221_ (_05897_, _05501_, _05379_);
  nor _14222_ (_05898_, _05897_, _05896_);
  nor _14223_ (_05899_, _05898_, _05895_);
  nor _14224_ (_05900_, _05899_, _05894_);
  nor _14225_ (_05901_, _05381_, _05379_);
  and _14226_ (_05902_, _05379_, _05376_);
  nor _14227_ (_05903_, _05902_, _05583_);
  nor _14228_ (_05904_, _05903_, _05515_);
  nor _14229_ (_05905_, _05904_, _05901_);
  not _14230_ (_05906_, _05905_);
  and _14231_ (_05907_, _05362_, _05514_);
  and _14232_ (_05908_, _05535_, _05907_);
  and _14233_ (_05909_, _05362_, _05354_);
  not _14234_ (_05910_, _05379_);
  and _14235_ (_05911_, _05910_, _05909_);
  nor _14236_ (_05912_, _05911_, _05355_);
  and _14237_ (_05913_, _05912_, _05381_);
  nor _14238_ (_05914_, _05504_, _05381_);
  nor _14239_ (_05915_, _05914_, _05913_);
  nor _14240_ (_05916_, _05915_, _05908_);
  and _14241_ (_05917_, _05916_, _05906_);
  and _14242_ (_05918_, _05917_, _05900_);
  not _14243_ (_05919_, _05918_);
  nor _14244_ (_05920_, _05919_, _05891_);
  and _14245_ (_05921_, _05920_, _05882_);
  nand _14246_ (_05922_, _05921_, _05843_);
  nand _14247_ (_05923_, _05654_, _05922_);
  and _14248_ (_05924_, _05923_, _05655_);
  and _14249_ (_05925_, _05297_, _05167_);
  and _14250_ (_05926_, _05925_, _05211_);
  and _14251_ (_05927_, _05926_, _05649_);
  not _14252_ (_05928_, _05927_);
  nand _14253_ (_05929_, _05928_, _05924_);
  and _14254_ (_05930_, _05678_, _05382_);
  not _14255_ (_05931_, _05930_);
  and _14256_ (_05933_, _05684_, _05381_);
  nor _14257_ (_05934_, _05933_, _05510_);
  and _14258_ (_05935_, _05934_, _05931_);
  not _14259_ (_05936_, _05678_);
  nor _14260_ (_05937_, _05472_, _05373_);
  and _14261_ (_05938_, _05884_, _05937_);
  nor _14262_ (_05939_, _05938_, _05382_);
  nor _14263_ (_05940_, _05476_, _05346_);
  and _14264_ (_05941_, _05940_, _05759_);
  nand _14265_ (_05942_, _05941_, _05716_);
  and _14266_ (_05943_, _05942_, _05382_);
  nor _14267_ (_05944_, _05943_, _05939_);
  and _14268_ (_05945_, _05944_, _05936_);
  nor _14269_ (_05946_, _05944_, _05936_);
  nor _14270_ (_05947_, _05946_, _05945_);
  and _14271_ (_05948_, _05947_, _05481_);
  nor _14272_ (_05949_, _05948_, _05935_);
  and _14273_ (_05950_, _05691_, _05485_);
  and _14274_ (_05951_, _05688_, _05501_);
  nor _14275_ (_05952_, _05689_, _05516_);
  and _14276_ (_05953_, _05678_, _05504_);
  or _14277_ (_05954_, _05953_, _05952_);
  or _14278_ (_05955_, _05954_, _05951_);
  nor _14279_ (_05956_, _05955_, _05950_);
  nor _14280_ (_05957_, _05678_, _05370_);
  not _14281_ (_05958_, _05957_);
  and _14282_ (_05959_, _05958_, _05956_);
  and _14283_ (_05960_, _05959_, _05949_);
  nand _14284_ (_05961_, _05960_, _05927_);
  and _14285_ (_05962_, _05961_, _05141_);
  and _14286_ (_07206_, _05962_, _05929_);
  not _14287_ (_05963_, _05922_);
  and _14288_ (_05964_, _05651_, _05275_);
  and _14289_ (_05965_, _05964_, _05649_);
  and _14290_ (_05966_, _05965_, _05647_);
  nand _14291_ (_05967_, _05966_, _05963_);
  not _14292_ (_05968_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _14293_ (_05969_, _05968_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not _14294_ (_05970_, _05634_);
  nor _14295_ (_05971_, _05641_, _05628_);
  not _14296_ (_05972_, _05971_);
  or _14297_ (_05973_, _05972_, _05638_);
  or _14298_ (_05974_, _05973_, _05970_);
  and _14299_ (_05975_, _05974_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _14300_ (_05976_, _05975_, _05969_);
  or _14301_ (_05977_, _05976_, _05966_);
  and _14302_ (_05978_, _05977_, _05928_);
  and _14303_ (_05979_, _05978_, _05967_);
  nor _14304_ (_05980_, _05758_, _05381_);
  nor _14305_ (_05981_, _05768_, _05382_);
  or _14306_ (_05982_, _05981_, _05980_);
  and _14307_ (_05983_, _05982_, _05509_);
  not _14308_ (_05984_, _05937_);
  nand _14309_ (_05985_, _05984_, _05477_);
  and _14310_ (_05986_, _05985_, _05508_);
  nand _14311_ (_05987_, _05986_, _05759_);
  or _14312_ (_05988_, _05986_, _05759_);
  and _14313_ (_05989_, _05988_, _05481_);
  and _14314_ (_05990_, _05989_, _05987_);
  nor _14315_ (_05991_, _05990_, _05983_);
  nor _14316_ (_05992_, _05758_, _05370_);
  not _14317_ (_05993_, _05992_);
  and _14318_ (_05994_, _05775_, _05485_);
  not _14319_ (_05995_, _05994_);
  nor _14320_ (_05996_, _05774_, _05516_);
  not _14321_ (_05997_, _05996_);
  and _14322_ (_05998_, _05773_, _05501_);
  and _14323_ (_05999_, _05758_, _05504_);
  nor _14324_ (_06000_, _05999_, _05998_);
  and _14325_ (_06001_, _06000_, _05997_);
  and _14326_ (_06002_, _06001_, _05995_);
  and _14327_ (_06003_, _06002_, _05993_);
  nand _14328_ (_06004_, _06003_, _05991_);
  and _14329_ (_06005_, _06004_, _05927_);
  or _14330_ (_06006_, _06005_, _05979_);
  and _14331_ (_07277_, _06006_, _05141_);
  not _14332_ (_06007_, _05186_);
  and _14333_ (_06008_, _05650_, _06007_);
  and _14334_ (_06009_, _05280_, _05227_);
  and _14335_ (_06010_, _05647_, _05241_);
  nor _14336_ (_06011_, _05256_, _05172_);
  and _14337_ (_06012_, _06011_, _06010_);
  and _14338_ (_06013_, _06012_, _06009_);
  and _14339_ (_06014_, _06013_, _06008_);
  nand _14340_ (_06015_, _06014_, _05963_);
  nor _14341_ (_06016_, _05266_, _05256_);
  and _14342_ (_06017_, _06016_, _05648_);
  and _14343_ (_06018_, _05925_, _05172_);
  and _14344_ (_06019_, _06018_, _06008_);
  and _14345_ (_06020_, _06019_, _06017_);
  not _14346_ (_06021_, _06020_);
  or _14347_ (_06022_, _06014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _14348_ (_06023_, _06022_, _06021_);
  and _14349_ (_06024_, _06023_, _06015_);
  nor _14350_ (_06025_, _06021_, _05960_);
  or _14351_ (_06026_, _06025_, _06024_);
  and _14352_ (_07297_, _06026_, _05141_);
  and _14353_ (_06027_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand _14354_ (_06028_, _05633_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _14355_ (_06030_, _06028_, _05973_);
  and _14356_ (_06031_, _06030_, _06027_);
  and _14357_ (_06032_, _05650_, _05186_);
  and _14358_ (_06033_, _06032_, _05173_);
  and _14359_ (_06034_, _06033_, _05649_);
  and _14360_ (_06035_, _06034_, _05647_);
  or _14361_ (_06036_, _06035_, _06031_);
  and _14362_ (_06037_, _06036_, _05928_);
  nand _14363_ (_06038_, _06035_, _05963_);
  and _14364_ (_06039_, _06038_, _06037_);
  nor _14365_ (_06040_, _05795_, _05510_);
  nand _14366_ (_06041_, _05471_, _05381_);
  or _14367_ (_06042_, _05475_, _05381_);
  nand _14368_ (_06043_, _06042_, _06041_);
  nand _14369_ (_06044_, _06043_, _05404_);
  or _14370_ (_06045_, _06043_, _05404_);
  and _14371_ (_06046_, _06045_, _05481_);
  and _14372_ (_06047_, _06046_, _06044_);
  nor _14373_ (_06048_, _06047_, _06040_);
  nor _14374_ (_06049_, _05404_, _05370_);
  not _14375_ (_06050_, _06049_);
  and _14376_ (_06051_, _05798_, _05485_);
  not _14377_ (_06052_, _06051_);
  nor _14378_ (_06053_, _05797_, _05516_);
  not _14379_ (_06054_, _06053_);
  and _14380_ (_06055_, _05796_, _05501_);
  and _14381_ (_06056_, _05504_, _05404_);
  nor _14382_ (_06057_, _06056_, _06055_);
  and _14383_ (_06059_, _06057_, _06054_);
  and _14384_ (_06060_, _06059_, _06052_);
  and _14385_ (_06061_, _06060_, _06050_);
  and _14386_ (_06062_, _06061_, _06048_);
  nor _14387_ (_06063_, _06062_, _05928_);
  or _14388_ (_06064_, _06063_, _06039_);
  and _14389_ (_07616_, _06064_, _05141_);
  and _14390_ (_06065_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _14391_ (_06066_, _06065_);
  and _14392_ (_06067_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _05630_);
  and _14393_ (_06068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _14394_ (_06069_, _06068_, _06067_);
  and _14395_ (_06070_, _06069_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _14396_ (_06071_, _06070_, _05628_);
  and _14397_ (_06072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _14398_ (_06073_, _06072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _14399_ (_06074_, _06073_);
  and _14400_ (_06075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _14401_ (_06076_, _06075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _14402_ (_06077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _14403_ (_06078_, _06077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _14404_ (_06080_, _06078_, _06076_);
  and _14405_ (_06081_, _06080_, _06074_);
  not _14406_ (_06082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _14407_ (_06083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _14408_ (_06084_, _06083_, _06082_);
  nand _14409_ (_06085_, _06084_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _14410_ (_06086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _14411_ (_06087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _14412_ (_06088_, _06087_, _06086_);
  and _14413_ (_06089_, _06088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _14414_ (_06090_, _06089_);
  and _14415_ (_06091_, _06090_, _06085_);
  and _14416_ (_06092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _14417_ (_06093_, _06092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _14418_ (_06094_, _06093_);
  and _14419_ (_06095_, _06094_, _06091_);
  and _14420_ (_06096_, _06095_, _06081_);
  nor _14421_ (_06097_, _06096_, _06071_);
  and _14422_ (_06098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _05628_);
  not _14423_ (_06099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _14424_ (_06100_, _06084_, _06099_);
  not _14425_ (_06101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _14426_ (_06102_, _06088_, _06101_);
  nor _14427_ (_06103_, _06102_, _06100_);
  not _14428_ (_06104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _14429_ (_06105_, _06092_, _06104_);
  not _14430_ (_06106_, _06105_);
  not _14431_ (_06107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _14432_ (_06109_, _06072_, _06107_);
  not _14433_ (_06110_, _06109_);
  not _14434_ (_06111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _14435_ (_06112_, _06075_, _06111_);
  not _14436_ (_06113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _14437_ (_06114_, _06077_, _06113_);
  nor _14438_ (_06115_, _06114_, _06112_);
  and _14439_ (_06116_, _06115_, _06110_);
  and _14440_ (_06117_, _06116_, _06106_);
  nand _14441_ (_06118_, _06117_, _06103_);
  nand _14442_ (_06119_, _06118_, _06098_);
  not _14443_ (_06120_, _06119_);
  nor _14444_ (_06121_, _06120_, _06097_);
  and _14445_ (_06122_, _06121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not _14446_ (_06123_, _06097_);
  nor _14447_ (_06124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05630_);
  and _14448_ (_06125_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05630_);
  nor _14449_ (_06126_, _06125_, _06124_);
  nor _14450_ (_06127_, _06126_, _06123_);
  or _14451_ (_06128_, _06127_, _06122_);
  and _14452_ (_06129_, _06128_, _06066_);
  and _14453_ (_06130_, _06126_, _06065_);
  or _14454_ (_06131_, _06130_, _06129_);
  and _14455_ (_07816_, _06131_, _05141_);
  or _14456_ (_06132_, _06081_, _06071_);
  nor _14457_ (_06133_, _06119_, _06097_);
  not _14458_ (_06134_, _06133_);
  or _14459_ (_06135_, _06134_, _06116_);
  and _14460_ (_06136_, _06135_, _06132_);
  nor _14461_ (_06137_, _06065_, _05630_);
  not _14462_ (_06138_, _06137_);
  or _14463_ (_06139_, _06138_, _06136_);
  not _14464_ (_06140_, _06103_);
  and _14465_ (_06141_, _06140_, _06098_);
  and _14466_ (_06142_, _06105_, _06098_);
  or _14467_ (_06143_, _06142_, _06141_);
  or _14468_ (_06144_, _06143_, _06097_);
  not _14469_ (_06145_, _06095_);
  or _14470_ (_06146_, _06132_, _06145_);
  and _14471_ (_06147_, _06146_, _06137_);
  and _14472_ (_06148_, _06147_, _06144_);
  or _14473_ (_06150_, _06148_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _14474_ (_06151_, _06150_, _05141_);
  and _14475_ (_07981_, _06151_, _06139_);
  nor _14476_ (_06152_, _05277_, _05269_);
  and _14477_ (_06153_, _05292_, _06152_);
  or _14478_ (_06154_, _06153_, _05572_);
  and _14479_ (_06155_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nand _14480_ (_06156_, _05301_, _06152_);
  and _14481_ (_06157_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _14482_ (_06158_, _06157_, _06156_);
  nor _14483_ (_06159_, _05446_, _05370_);
  not _14484_ (_06160_, _06159_);
  or _14485_ (_06161_, _05446_, _05381_);
  and _14486_ (_06162_, _05538_, _06161_);
  or _14487_ (_06163_, _06162_, _05425_);
  nand _14488_ (_06164_, _06162_, _05425_);
  and _14489_ (_06165_, _06164_, _05481_);
  nand _14490_ (_06166_, _06165_, _06163_);
  or _14491_ (_06167_, _05810_, _05808_);
  or _14492_ (_06168_, _06167_, _05583_);
  or _14493_ (_06169_, _05808_, _05516_);
  nand _14494_ (_06170_, _05810_, _05501_);
  and _14495_ (_06171_, _05809_, _05509_);
  and _14496_ (_06172_, _05504_, _05446_);
  nor _14497_ (_06173_, _06172_, _06171_);
  and _14498_ (_06174_, _06173_, _06170_);
  and _14499_ (_06175_, _06174_, _06169_);
  and _14500_ (_06176_, _06175_, _06168_);
  and _14501_ (_06177_, _06176_, _06166_);
  and _14502_ (_06178_, _06177_, _06160_);
  not _14503_ (_06179_, _06178_);
  and _14504_ (_06180_, _05297_, _05291_);
  and _14505_ (_06181_, _06180_, _06179_);
  or _14506_ (_06182_, _06181_, _06158_);
  or _14507_ (_06183_, _06182_, _06155_);
  and _14508_ (_08821_, _06183_, _05141_);
  and _14509_ (_06184_, _05649_, _05289_);
  and _14510_ (_06185_, _06184_, _05647_);
  nand _14511_ (_06186_, _06185_, _05963_);
  not _14512_ (_06187_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _14513_ (_06188_, _05971_, _05638_);
  or _14514_ (_06189_, _06188_, _06028_);
  and _14515_ (_06190_, _06189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _14516_ (_06191_, _06190_, _06187_);
  or _14517_ (_06192_, _06191_, _06185_);
  and _14518_ (_06193_, _06192_, _05928_);
  and _14519_ (_06194_, _06193_, _06186_);
  nor _14520_ (_06195_, _06178_, _05928_);
  or _14521_ (_06197_, _06195_, _06194_);
  and _14522_ (_08859_, _06197_, _05141_);
  and _14523_ (_09119_, _05141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nand _14524_ (_06198_, _06119_, _05628_);
  or _14525_ (_06199_, _06198_, _06097_);
  nand _14526_ (_06200_, _06124_, _06065_);
  and _14527_ (_06201_, _06200_, _05141_);
  and _14528_ (_10115_, _06201_, _06199_);
  and _14529_ (_06202_, _05266_, _05227_);
  and _14530_ (_06203_, _05256_, _05173_);
  and _14531_ (_06204_, _06010_, _06203_);
  and _14532_ (_06205_, _06204_, _06202_);
  and _14533_ (_06206_, _05274_, _05197_);
  and _14534_ (_06207_, _06206_, _06007_);
  and _14535_ (_06208_, _05922_, _06207_);
  nor _14536_ (_06209_, _05186_, _05208_);
  nand _14537_ (_06210_, _05197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _14538_ (_06211_, _06210_, _06209_);
  or _14539_ (_06212_, _06211_, _06208_);
  and _14540_ (_06213_, _06212_, _06205_);
  nand _14541_ (_06214_, _06205_, _05197_);
  and _14542_ (_06215_, _06214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _14543_ (_06216_, _06215_, _05927_);
  or _14544_ (_06217_, _06216_, _06213_);
  nor _14545_ (_06218_, _05724_, _05382_);
  nor _14546_ (_06219_, _05715_, _05381_);
  or _14547_ (_06220_, _06219_, _06218_);
  and _14548_ (_06221_, _06220_, _05509_);
  or _14549_ (_06222_, _05941_, _05716_);
  nand _14550_ (_06223_, _06222_, _05943_);
  nand _14551_ (_06224_, _05758_, _05937_);
  and _14552_ (_06225_, _06224_, _05716_);
  or _14553_ (_06226_, _06225_, _05938_);
  nand _14554_ (_06227_, _06226_, _05381_);
  nand _14555_ (_06228_, _06227_, _06223_);
  and _14556_ (_06229_, _06228_, _05481_);
  nor _14557_ (_06230_, _06229_, _06221_);
  nor _14558_ (_06231_, _05715_, _05370_);
  not _14559_ (_06233_, _06231_);
  and _14560_ (_06234_, _05730_, _05485_);
  not _14561_ (_06235_, _06234_);
  nor _14562_ (_06236_, _05728_, _05516_);
  not _14563_ (_06237_, _06236_);
  and _14564_ (_06238_, _05727_, _05501_);
  and _14565_ (_06239_, _05715_, _05504_);
  nor _14566_ (_06240_, _06239_, _06238_);
  and _14567_ (_06241_, _06240_, _06237_);
  and _14568_ (_06242_, _06241_, _06235_);
  and _14569_ (_06243_, _06242_, _06233_);
  and _14570_ (_06244_, _06243_, _06230_);
  nand _14571_ (_06245_, _06244_, _05927_);
  and _14572_ (_06246_, _06245_, _05141_);
  and _14573_ (_10153_, _06246_, _06217_);
  nor _14574_ (_06247_, _06065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _14575_ (_06248_, _06247_);
  or _14576_ (_06249_, _06248_, _06136_);
  and _14577_ (_06250_, _06247_, _06146_);
  and _14578_ (_06251_, _06250_, _06144_);
  or _14579_ (_06253_, _06251_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _14580_ (_06254_, _06253_, _05141_);
  and _14581_ (_10191_, _06254_, _06249_);
  and _14582_ (_06255_, _06204_, _06009_);
  and _14583_ (_06256_, _06255_, _06008_);
  nand _14584_ (_06257_, _06256_, _05963_);
  or _14585_ (_06259_, _06256_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _14586_ (_06260_, _05280_, _05256_);
  and _14587_ (_06261_, _06260_, _05648_);
  and _14588_ (_06262_, _06261_, _05926_);
  not _14589_ (_06263_, _06262_);
  and _14590_ (_06264_, _06263_, _06259_);
  and _14591_ (_06265_, _06264_, _06257_);
  nor _14592_ (_06266_, _06263_, _05960_);
  or _14593_ (_06267_, _06266_, _06265_);
  and _14594_ (_10239_, _06267_, _05141_);
  or _14595_ (_06268_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _14596_ (_06269_, _06268_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor _14597_ (_06270_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and _14598_ (_06271_, _06270_, _05143_);
  and _14599_ (_06272_, _06271_, _06269_);
  and _14600_ (pc_log_change, _06272_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _14601_ (_06273_, _06004_, _05576_);
  not _14602_ (_06274_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _14603_ (_06275_, _05576_, _05297_);
  nor _14604_ (_06276_, _06275_, _06274_);
  or _14605_ (_06277_, _06276_, _06273_);
  or _14606_ (_06278_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _14607_ (_06279_, _06278_, _05141_);
  and _14608_ (_12316_, _06279_, _06277_);
  and _14609_ (_06280_, _05569_, _05297_);
  or _14610_ (_06281_, _06280_, _05574_);
  and _14611_ (_06282_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  not _14612_ (_06283_, _06244_);
  and _14613_ (_06284_, _06275_, _06283_);
  or _14614_ (_06285_, _06284_, _06282_);
  and _14615_ (_12641_, _06285_, _05141_);
  and _14616_ (_06286_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _14617_ (_06287_, _06275_, _05522_);
  or _14618_ (_06288_, _06287_, _06286_);
  and _14619_ (_12994_, _06288_, _05141_);
  and _14620_ (_06289_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  not _14621_ (_06290_, _06062_);
  and _14622_ (_06291_, _06275_, _06290_);
  or _14623_ (_06292_, _06291_, _06289_);
  and _14624_ (_00302_, _06292_, _05141_);
  and _14625_ (_06293_, _05141_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _14626_ (_06295_, _06293_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _14627_ (_06296_, _06271_, _05141_);
  and _14628_ (_06297_, _06269_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _14629_ (_06298_, _06297_, _06272_);
  not _14630_ (_06299_, _06298_);
  not _14631_ (_06300_, _06272_);
  not _14632_ (_06301_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  not _14633_ (_06302_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or _14634_ (_06303_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or _14635_ (_06304_, _06303_, _06302_);
  or _14636_ (_06305_, _06304_, _06301_);
  not _14637_ (_06306_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nand _14638_ (_06307_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or _14639_ (_06308_, _06307_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or _14640_ (_06309_, _06308_, _06306_);
  and _14641_ (_06310_, _06309_, _06305_);
  not _14642_ (_06311_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not _14643_ (_06312_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _14644_ (_06313_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _06302_);
  nand _14645_ (_06314_, _06313_, _06312_);
  or _14646_ (_06315_, _06314_, _06311_);
  and _14647_ (_06316_, _06315_, _06310_);
  not _14648_ (_06317_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _14649_ (_06318_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _14650_ (_06319_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], _06318_);
  nand _14651_ (_06320_, _06319_, _06302_);
  not _14652_ (_06321_, _06320_);
  nand _14653_ (_06322_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _14654_ (_06323_, _06322_, _06317_);
  not _14655_ (_06324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _14656_ (_06325_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or _14657_ (_06326_, _06325_, _06302_);
  or _14658_ (_06327_, _06326_, _06324_);
  and _14659_ (_06328_, _06325_, _06302_);
  nand _14660_ (_06329_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _14661_ (_06330_, _06329_, _06327_);
  and _14662_ (_06331_, _06330_, _06323_);
  nand _14663_ (_06332_, _06331_, _06316_);
  or _14664_ (_06333_, _06332_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14665_ (_06334_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14666_ (_06335_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _06334_);
  not _14667_ (_06336_, _06335_);
  and _14668_ (_06337_, _06336_, _06333_);
  or _14669_ (_06338_, _06337_, _06300_);
  nand _14670_ (_06339_, _06338_, _06299_);
  and _14671_ (_06340_, _06269_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _14672_ (_06341_, _06340_, _06272_);
  not _14673_ (_06342_, _06341_);
  not _14674_ (_06343_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _14675_ (_06344_, _06308_, _06343_);
  nand _14676_ (_06345_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _14677_ (_06346_, _06345_, _06344_);
  not _14678_ (_06347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _14679_ (_06348_, _06326_, _06347_);
  nand _14680_ (_06349_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _14681_ (_06350_, _06349_, _06348_);
  not _14682_ (_06351_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or _14683_ (_06352_, _06304_, _06351_);
  not _14684_ (_06353_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _14685_ (_06354_, _06314_, _06353_);
  and _14686_ (_06355_, _06354_, _06352_);
  and _14687_ (_06356_, _06355_, _06350_);
  nand _14688_ (_06357_, _06356_, _06346_);
  nand _14689_ (_06358_, _06357_, _06317_);
  nand _14690_ (_06360_, _06358_, _06334_);
  nor _14691_ (_06361_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _06334_);
  not _14692_ (_06362_, _06361_);
  and _14693_ (_06363_, _06362_, _06360_);
  or _14694_ (_06364_, _06363_, _06300_);
  nand _14695_ (_06365_, _06364_, _06342_);
  and _14696_ (_06366_, _06365_, _06339_);
  and _14697_ (_06367_, _06269_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _14698_ (_06368_, _06367_, _06272_);
  not _14699_ (_06369_, _06368_);
  not _14700_ (_06370_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _14701_ (_06371_, _06314_, _06370_);
  nand _14702_ (_06372_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _14703_ (_06373_, _06372_, _06371_);
  not _14704_ (_06374_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _14705_ (_06375_, _06308_, _06374_);
  not _14706_ (_06376_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or _14707_ (_06377_, _06304_, _06376_);
  and _14708_ (_06378_, _06377_, _06375_);
  not _14709_ (_06379_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _14710_ (_06380_, _06326_, _06379_);
  nand _14711_ (_06381_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _14712_ (_06382_, _06381_, _06380_);
  and _14713_ (_06383_, _06382_, _06378_);
  nand _14714_ (_06384_, _06383_, _06373_);
  nand _14715_ (_06385_, _06384_, _06317_);
  nand _14716_ (_06386_, _06385_, _06334_);
  nor _14717_ (_06387_, _06334_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  not _14718_ (_06388_, _06387_);
  and _14719_ (_06389_, _06388_, _06386_);
  or _14720_ (_06390_, _06389_, _06300_);
  and _14721_ (_06391_, _06390_, _06369_);
  and _14722_ (_06392_, _06269_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _14723_ (_06393_, _06392_, _06272_);
  not _14724_ (_06394_, _06393_);
  not _14725_ (_06395_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _14726_ (_06396_, _06308_, _06395_);
  nand _14727_ (_06397_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _14728_ (_06398_, _06397_, _06396_);
  not _14729_ (_06399_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _14730_ (_06400_, _06326_, _06399_);
  nand _14731_ (_06401_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _14732_ (_06402_, _06401_, _06400_);
  not _14733_ (_06403_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or _14734_ (_06404_, _06304_, _06403_);
  not _14735_ (_06406_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _14736_ (_06407_, _06314_, _06406_);
  and _14737_ (_06408_, _06407_, _06404_);
  and _14738_ (_06409_, _06408_, _06402_);
  and _14739_ (_06410_, _06409_, _06398_);
  or _14740_ (_06411_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _14741_ (_06412_, _06411_, _06410_);
  and _14742_ (_06413_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  not _14743_ (_06414_, _06413_);
  and _14744_ (_06415_, _06414_, _06412_);
  nand _14745_ (_06416_, _06415_, _06272_);
  and _14746_ (_06417_, _06416_, _06394_);
  not _14747_ (_06418_, _06417_);
  and _14748_ (_06419_, _06418_, _06391_);
  and _14749_ (_06420_, _06419_, _06366_);
  and _14750_ (_06421_, _06269_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _14751_ (_06422_, _06421_, _06272_);
  not _14752_ (_06423_, _06422_);
  not _14753_ (_06425_, _06326_);
  and _14754_ (_06426_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not _14755_ (_06427_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _14756_ (_06428_, _06304_, _06427_);
  not _14757_ (_06429_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _14758_ (_06430_, _06308_, _06429_);
  nand _14759_ (_06431_, _06430_, _06428_);
  nor _14760_ (_06432_, _06431_, _06426_);
  nand _14761_ (_06433_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not _14762_ (_06434_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _14763_ (_06436_, _06320_, _06434_);
  and _14764_ (_06437_, _06436_, _06433_);
  not _14765_ (_06438_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _14766_ (_06439_, _06314_, _06438_);
  and _14767_ (_06440_, _06439_, _06317_);
  and _14768_ (_06441_, _06440_, _06437_);
  nand _14769_ (_06442_, _06441_, _06432_);
  or _14770_ (_06444_, _06442_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14771_ (_06445_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _06334_);
  not _14772_ (_06446_, _06445_);
  and _14773_ (_06447_, _06446_, _06444_);
  or _14774_ (_06448_, _06447_, _06300_);
  and _14775_ (_06449_, _06448_, _06423_);
  not _14776_ (_06450_, _06449_);
  and _14777_ (_06451_, _06269_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _14778_ (_06452_, _06451_, _06272_);
  not _14779_ (_06453_, _06452_);
  nand _14780_ (_06454_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _14781_ (_06455_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _14782_ (_06456_, _06455_, _06454_);
  not _14783_ (_06457_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _14784_ (_06458_, _06326_, _06457_);
  not _14785_ (_06459_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or _14786_ (_06460_, _06304_, _06459_);
  and _14787_ (_06461_, _06460_, _06458_);
  not _14788_ (_06462_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _14789_ (_06463_, _06308_, _06462_);
  not _14790_ (_06464_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _14791_ (_06465_, _06314_, _06464_);
  and _14792_ (_06466_, _06465_, _06463_);
  and _14793_ (_06467_, _06466_, _06461_);
  and _14794_ (_06468_, _06467_, _06456_);
  or _14795_ (_06469_, _06468_, _06411_);
  and _14796_ (_06470_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  not _14797_ (_06471_, _06470_);
  and _14798_ (_06472_, _06471_, _06469_);
  nand _14799_ (_06473_, _06472_, _06272_);
  and _14800_ (_06474_, _06473_, _06453_);
  and _14801_ (_06475_, _06269_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _14802_ (_06476_, _06475_, _06272_);
  not _14803_ (_06477_, _06476_);
  nor _14804_ (_06478_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _14805_ (_06479_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand _14806_ (_06480_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _14807_ (_06481_, _06480_, _06479_);
  not _14808_ (_06482_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _14809_ (_06483_, _06326_, _06482_);
  not _14810_ (_06484_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _14811_ (_06485_, _06308_, _06484_);
  and _14812_ (_06486_, _06485_, _06483_);
  not _14813_ (_06487_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or _14814_ (_06488_, _06304_, _06487_);
  not _14815_ (_06489_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _14816_ (_06490_, _06314_, _06489_);
  and _14817_ (_06491_, _06490_, _06488_);
  and _14818_ (_06492_, _06491_, _06486_);
  nand _14819_ (_06493_, _06492_, _06481_);
  nand _14820_ (_06494_, _06493_, _06478_);
  and _14821_ (_06495_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not _14822_ (_06496_, _06495_);
  nand _14823_ (_06497_, _06496_, _06494_);
  or _14824_ (_06498_, _06497_, _06300_);
  and _14825_ (_06499_, _06498_, _06477_);
  and _14826_ (_06500_, _06269_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _14827_ (_06501_, _06500_, _06272_);
  not _14828_ (_06502_, _06501_);
  nand _14829_ (_06504_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _14830_ (_06505_, _06321_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _14831_ (_06506_, _06505_, _06504_);
  not _14832_ (_06508_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _14833_ (_06509_, _06326_, _06508_);
  not _14834_ (_06510_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _14835_ (_06511_, _06308_, _06510_);
  and _14836_ (_06512_, _06511_, _06509_);
  not _14837_ (_06514_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or _14838_ (_06515_, _06304_, _06514_);
  not _14839_ (_06516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _14840_ (_06517_, _06314_, _06516_);
  and _14841_ (_06518_, _06517_, _06515_);
  and _14842_ (_06519_, _06518_, _06512_);
  and _14843_ (_06520_, _06519_, _06506_);
  or _14844_ (_06521_, _06520_, _06411_);
  and _14845_ (_06522_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  not _14846_ (_06523_, _06522_);
  nand _14847_ (_06524_, _06523_, _06521_);
  or _14848_ (_06525_, _06524_, _06300_);
  and _14849_ (_06526_, _06525_, _06502_);
  and _14850_ (_06527_, _06526_, _06499_);
  and _14851_ (_06528_, _06527_, _06474_);
  and _14852_ (_06529_, _06528_, _06450_);
  and _14853_ (_06530_, _06529_, _06420_);
  and _14854_ (_06531_, _06364_, _06342_);
  and _14855_ (_06532_, _06338_, _06299_);
  nand _14856_ (_06533_, _06390_, _06369_);
  and _14857_ (_06534_, _06533_, _06532_);
  and _14858_ (_06535_, _06534_, _06418_);
  and _14859_ (_06536_, _06535_, _06531_);
  nand _14860_ (_06537_, _06498_, _06477_);
  nand _14861_ (_06538_, _06525_, _06502_);
  and _14862_ (_06539_, _06538_, _06537_);
  and _14863_ (_06540_, _06539_, _06474_);
  and _14864_ (_06541_, _06540_, _06536_);
  and _14865_ (_06542_, _06541_, _06450_);
  or _14866_ (_06543_, _06542_, _06530_);
  and _14867_ (_06544_, _06535_, _06365_);
  and _14868_ (_06545_, _06526_, _06537_);
  and _14869_ (_06546_, _06545_, _06474_);
  and _14870_ (_06547_, _06546_, _06450_);
  and _14871_ (_06548_, _06547_, _06544_);
  and _14872_ (_06549_, _06418_, _06533_);
  and _14873_ (_06550_, _06549_, _06366_);
  not _14874_ (_06551_, _06474_);
  and _14875_ (_06552_, _06539_, _06551_);
  and _14876_ (_06553_, _06552_, _06449_);
  and _14877_ (_06554_, _06553_, _06550_);
  and _14878_ (_06555_, _06538_, _06499_);
  and _14879_ (_06556_, _06555_, _06551_);
  and _14880_ (_06557_, _06556_, _06450_);
  and _14881_ (_06558_, _06557_, _06550_);
  or _14882_ (_06559_, _06558_, _06554_);
  and _14883_ (_06560_, _06547_, _06536_);
  or _14884_ (_06561_, _06560_, _06559_);
  or _14885_ (_06562_, _06561_, _06548_);
  and _14886_ (_06563_, _06545_, _06551_);
  and _14887_ (_06564_, _06563_, _06449_);
  and _14888_ (_06565_, _06563_, _06450_);
  and _14889_ (_06566_, _06556_, _06449_);
  or _14890_ (_06567_, _06566_, _06565_);
  or _14891_ (_06568_, _06567_, _06564_);
  and _14892_ (_06569_, _06568_, _06550_);
  and _14893_ (_06570_, _06546_, _06449_);
  and _14894_ (_06571_, _06570_, _06535_);
  and _14895_ (_06572_, _06540_, _06450_);
  and _14896_ (_06573_, _06550_, _06572_);
  and _14897_ (_06574_, _06527_, _06551_);
  and _14898_ (_06575_, _06574_, _06550_);
  or _14899_ (_06576_, _06575_, _06573_);
  or _14900_ (_06577_, _06576_, _06571_);
  or _14901_ (_06578_, _06577_, _06569_);
  or _14902_ (_06579_, _06578_, _06562_);
  or _14903_ (_06580_, _06579_, _06543_);
  and _14904_ (_06581_, _06580_, _06296_);
  or _14905_ (_00855_, _06581_, _06295_);
  nor _14906_ (_06582_, _05858_, _05856_);
  not _14907_ (_06583_, _06582_);
  nor _14908_ (_06584_, _05859_, _05845_);
  and _14909_ (_06585_, _06584_, _06583_);
  not _14910_ (_06586_, _06585_);
  nor _14911_ (_06587_, _05827_, _05821_);
  nor _14912_ (_06588_, _06587_, _05828_);
  nor _14913_ (_06589_, _06588_, _05657_);
  not _14914_ (_06590_, _06589_);
  not _14915_ (_06591_, _05883_);
  nor _14916_ (_06592_, _05887_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _14917_ (_06593_, _06592_, _05537_);
  nor _14918_ (_06594_, _06593_, _05469_);
  and _14919_ (_06595_, _05470_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _14920_ (_06596_, _06595_, _06594_);
  nor _14921_ (_06597_, _06596_, _06591_);
  not _14922_ (_06598_, _05355_);
  nor _14923_ (_06599_, _05469_, _06598_);
  and _14924_ (_06600_, _05354_, _05357_);
  and _14925_ (_06601_, _06600_, ABINPUT000000[3]);
  nor _14926_ (_06602_, _06601_, _06599_);
  not _14927_ (_06603_, _05363_);
  or _14928_ (_06604_, _05404_, _06603_);
  and _14929_ (_06605_, _05537_, _05367_);
  and _14930_ (_06606_, _05500_, _05349_);
  and _14931_ (_06607_, _06606_, ABINPUT000[3]);
  nor _14932_ (_06608_, _06607_, _06605_);
  and _14933_ (_06610_, _06608_, _06604_);
  and _14934_ (_06611_, _06610_, _06602_);
  and _14935_ (_06612_, _06611_, _05557_);
  not _14936_ (_06613_, _06612_);
  nor _14937_ (_06614_, _06613_, _06597_);
  and _14938_ (_06615_, _06614_, _05545_);
  and _14939_ (_06616_, _06615_, _06590_);
  and _14940_ (_06617_, _06616_, _06586_);
  and _14941_ (_06618_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05143_);
  and _14942_ (_06619_, _06618_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _14943_ (_06620_, _06206_, _05186_);
  and _14944_ (_06621_, _06018_, _05649_);
  and _14945_ (_06622_, _06621_, _06620_);
  nor _14946_ (_06623_, _06622_, _06619_);
  not _14947_ (_06624_, _06623_);
  nand _14948_ (_06625_, _06624_, _06617_);
  or _14949_ (_06626_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _14950_ (_06627_, _06626_, _05141_);
  and _14951_ (_01188_, _06627_, _06625_);
  nor _14952_ (_06628_, _05715_, _06598_);
  or _14953_ (_06629_, _05678_, _06603_);
  nand _14954_ (_06630_, _06230_, _06629_);
  not _14955_ (_06631_, _05367_);
  nor _14956_ (_06632_, _05758_, _06631_);
  or _14957_ (_06633_, _06236_, _06234_);
  or _14958_ (_06634_, _06633_, _06632_);
  or _14959_ (_06635_, _06634_, _06630_);
  not _14960_ (_06636_, _05885_);
  and _14961_ (_06637_, _05887_, _05883_);
  nor _14962_ (_06638_, _06637_, _05381_);
  and _14963_ (_06639_, _06638_, _06636_);
  not _14964_ (_06640_, _06639_);
  and _14965_ (_06641_, _06637_, _05373_);
  and _14966_ (_06642_, _06641_, _05759_);
  nor _14967_ (_06643_, _06642_, _05716_);
  nor _14968_ (_06644_, _06643_, _06640_);
  nor _14969_ (_06645_, _06641_, _05759_);
  nor _14970_ (_06646_, _06639_, _06645_);
  and _14971_ (_06647_, _06646_, _05716_);
  not _14972_ (_06648_, _05884_);
  nor _14973_ (_06649_, _06641_, _06648_);
  and _14974_ (_06650_, _06640_, _06649_);
  or _14975_ (_06651_, _06650_, _06647_);
  nor _14976_ (_06652_, _06651_, _06644_);
  nor _14977_ (_06653_, _06652_, _06591_);
  and _14978_ (_06654_, _06600_, ABINPUT000000[7]);
  nor _14979_ (_06655_, _06654_, _06653_);
  nand _14980_ (_06656_, _06655_, _06240_);
  and _14981_ (_06657_, _05876_, _05870_);
  not _14982_ (_06658_, _06657_);
  and _14983_ (_06659_, _05877_, _05844_);
  and _14984_ (_06660_, _06659_, _06658_);
  and _14985_ (_06661_, _05838_, _05782_);
  nor _14986_ (_06662_, _06661_, _05839_);
  nor _14987_ (_06663_, _06662_, _05657_);
  and _14988_ (_06664_, _06606_, ABINPUT000[7]);
  or _14989_ (_06665_, _06664_, _06663_);
  or _14990_ (_06666_, _06665_, _06660_);
  or _14991_ (_06667_, _06666_, _06656_);
  or _14992_ (_06668_, _06667_, _06635_);
  or _14993_ (_06669_, _06668_, _06628_);
  or _14994_ (_06670_, _06669_, _06623_);
  or _14995_ (_06671_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _14996_ (_06672_, _06671_, _05141_);
  and _14997_ (_01207_, _06672_, _06670_);
  or _14998_ (_06674_, _05572_, _05279_);
  and _14999_ (_06675_, _06674_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nand _15000_ (_06676_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _15001_ (_06677_, _06676_, _05278_);
  and _15002_ (_06678_, _05297_, _05269_);
  and _15003_ (_06679_, _06678_, _06179_);
  or _15004_ (_06680_, _06679_, _06677_);
  or _15005_ (_06681_, _06680_, _06675_);
  and _15006_ (_02780_, _06681_, _05141_);
  not _15007_ (_06682_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor _15008_ (_06683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nor _15009_ (_06684_, _06683_, _06682_);
  and _15010_ (_06685_, _06684_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _15011_ (_06686_, _06685_);
  and _15012_ (_06687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _15013_ (_06688_, _06687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor _15014_ (_06689_, _06688_, _06686_);
  not _15015_ (_06690_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not _15016_ (_06691_, _06683_);
  and _15017_ (_06692_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _15018_ (_06693_, _06692_, _06691_);
  nor _15019_ (_06694_, _06693_, _06685_);
  or _15020_ (_06695_, _06694_, _06690_);
  or _15021_ (_06696_, _06695_, _06689_);
  and _15022_ (_06697_, _06685_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _15023_ (_06698_, _06697_, _06687_);
  or _15024_ (_06699_, _06698_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _15025_ (_06700_, _06699_, _05141_);
  and _15026_ (_03603_, _06700_, _06696_);
  not _15027_ (_06701_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _15028_ (_06702_, _06678_, _06701_);
  not _15029_ (_06703_, _05604_);
  and _15030_ (_06705_, _06678_, _06703_);
  or _15031_ (_06706_, _06705_, _06702_);
  and _15032_ (_03622_, _06706_, _05141_);
  and _15033_ (_06707_, _05297_, _05273_);
  not _15034_ (_06708_, _06707_);
  or _15035_ (_06709_, _06708_, _06004_);
  or _15036_ (_06710_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _15037_ (_06711_, _06710_, _05141_);
  and _15038_ (_03936_, _06711_, _06709_);
  nor _15039_ (_06713_, rst, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _15040_ (_06714_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _15041_ (_06715_, _05141_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _15042_ (_06716_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _15043_ (_04037_, _06716_, _06714_);
  and _15044_ (_06718_, _05522_, _05277_);
  not _15045_ (_06719_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _15046_ (_06720_, _05277_, _06719_);
  or _15047_ (_06721_, _06720_, _05572_);
  or _15048_ (_06722_, _06721_, _06718_);
  or _15049_ (_06723_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _15050_ (_06724_, _06723_, _05141_);
  and _15051_ (_04141_, _06724_, _06722_);
  and _15052_ (_06725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _15053_ (_06726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _15054_ (_06727_, _06726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _15055_ (_06728_, _06727_, _06725_);
  or _15056_ (_06729_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  not _15057_ (_06730_, _06728_);
  or _15058_ (_06731_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _15059_ (_06732_, _06731_, _06729_);
  and _15060_ (_06733_, _05241_, _05228_);
  and _15061_ (_06734_, _06733_, _05267_);
  not _15062_ (_06735_, _05925_);
  nor _15063_ (_06736_, _06735_, _05172_);
  and _15064_ (_06737_, _06736_, _06620_);
  and _15065_ (_06738_, _06737_, _06734_);
  or _15066_ (_06739_, _06738_, _06732_);
  nand _15067_ (_06740_, _06738_, _06178_);
  and _15068_ (_06741_, _06740_, _06739_);
  and _15069_ (_06742_, _06033_, _05925_);
  and _15070_ (_06743_, _06742_, _06734_);
  or _15071_ (_06744_, _06743_, _06741_);
  not _15072_ (_06745_, _06743_);
  or _15073_ (_06746_, _06745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _15074_ (_06747_, _06746_, _05141_);
  and _15075_ (_05132_, _06747_, _06744_);
  or _15076_ (_06748_, _06708_, _05522_);
  or _15077_ (_06749_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _15078_ (_06750_, _06749_, _05141_);
  and _15079_ (_05139_, _06750_, _06748_);
  nand _15080_ (_06751_, _06678_, _05560_);
  or _15081_ (_06752_, _06678_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _15082_ (_06753_, _06752_, _05141_);
  and _15083_ (_05140_, _06753_, _06751_);
  and _15084_ (_06754_, _06293_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _15085_ (_06755_, _06419_, _06339_);
  and _15086_ (_06756_, _06755_, _06553_);
  and _15087_ (_06757_, _06552_, _06450_);
  and _15088_ (_06758_, _06757_, _06420_);
  and _15089_ (_06759_, _06531_, _06339_);
  and _15090_ (_06760_, _06759_, _06419_);
  or _15091_ (_06761_, _06757_, _06570_);
  and _15092_ (_06762_, _06761_, _06760_);
  or _15093_ (_06763_, _06762_, _06758_);
  or _15094_ (_06764_, _06763_, _06756_);
  and _15095_ (_06765_, _06540_, _06449_);
  and _15096_ (_06766_, _06555_, _06474_);
  and _15097_ (_06767_, _06766_, _06449_);
  or _15098_ (_06768_, _06767_, _06765_);
  and _15099_ (_06769_, _06768_, _06420_);
  and _15100_ (_06770_, _06391_, _06532_);
  and _15101_ (_06771_, _06770_, _06418_);
  and _15102_ (_06772_, _06771_, _06552_);
  or _15103_ (_06773_, _06770_, _06417_);
  and _15104_ (_06774_, _06773_, _06767_);
  or _15105_ (_06775_, _06774_, _06772_);
  or _15106_ (_06776_, _06775_, _06769_);
  and _15107_ (_06777_, _06761_, _06417_);
  and _15108_ (_06778_, _06449_, _06417_);
  and _15109_ (_06779_, _06778_, _06552_);
  or _15110_ (_06780_, _06779_, _06777_);
  and _15111_ (_06781_, _06550_, _06765_);
  and _15112_ (_06782_, _06766_, _06450_);
  and _15113_ (_06784_, _06782_, _06536_);
  or _15114_ (_06785_, _06784_, _06781_);
  or _15115_ (_06786_, _06785_, _06780_);
  or _15116_ (_06787_, _06786_, _06776_);
  or _15117_ (_06788_, _06787_, _06764_);
  and _15118_ (_06789_, _06788_, _06296_);
  or _15119_ (_05235_, _06789_, _06754_);
  not _15120_ (_06790_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _15121_ (_06791_, \oc8051_top_1.oc8051_decoder1.state [0], _05143_);
  and _15122_ (_06792_, _06791_, _06790_);
  and _15123_ (_06793_, _06782_, _06420_);
  and _15124_ (_06795_, _06572_, _06420_);
  nor _15125_ (_06796_, _06795_, _06793_);
  not _15126_ (_06797_, _06796_);
  and _15127_ (_06798_, _06797_, _06792_);
  and _15128_ (_06799_, _06760_, _06572_);
  and _15129_ (_06800_, _06799_, _06270_);
  or _15130_ (_06801_, _06800_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _15131_ (_06802_, _06801_, _06798_);
  or _15132_ (_06803_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05143_);
  and _15133_ (_06804_, _06803_, _05141_);
  and _15134_ (_05238_, _06804_, _06802_);
  not _15135_ (_06805_, _06541_);
  and _15136_ (_06806_, _06550_, _06529_);
  nor _15137_ (_06807_, _06449_, _06417_);
  and _15138_ (_06808_, _06807_, _06534_);
  and _15139_ (_06809_, _06808_, _06528_);
  nor _15140_ (_06810_, _06809_, _06806_);
  and _15141_ (_06811_, _06810_, _06805_);
  not _15142_ (_06812_, _06811_);
  and _15143_ (_06813_, _06812_, _06792_);
  or _15144_ (_06814_, _06813_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _15145_ (_06815_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _15146_ (_06816_, _06759_, _06549_);
  and _15147_ (_06818_, _06816_, _06449_);
  and _15148_ (_06819_, _06553_, _06544_);
  or _15149_ (_06820_, _06819_, _06818_);
  or _15150_ (_06821_, _06270_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _15151_ (_06822_, _06821_, _06542_);
  or _15152_ (_06823_, _06822_, _06820_);
  and _15153_ (_06824_, _06823_, _06815_);
  or _15154_ (_06825_, _06824_, _06814_);
  or _15155_ (_06826_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05143_);
  and _15156_ (_06827_, _06826_, _05141_);
  and _15157_ (_05251_, _06827_, _06825_);
  and _15158_ (_06828_, _06528_, _06449_);
  nand _15159_ (_06829_, _06828_, _06550_);
  and _15160_ (_06830_, _06829_, _06811_);
  not _15161_ (_06831_, _06296_);
  and _15162_ (_06832_, _06535_, _06528_);
  or _15163_ (_06833_, _06832_, _06831_);
  or _15164_ (_05304_, _06833_, _06830_);
  not _15165_ (_06834_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _15166_ (_06835_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05143_);
  and _15167_ (_06836_, _06835_, _06834_);
  not _15168_ (_06837_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _15169_ (_06838_, _06618_, _06837_);
  and _15170_ (_06839_, _06733_, _06260_);
  and _15171_ (_06840_, _06839_, _05272_);
  and _15172_ (_06841_, _06840_, _05925_);
  nor _15173_ (_06842_, _06841_, _06838_);
  not _15174_ (_06843_, _05691_);
  and _15175_ (_06844_, _05840_, _06843_);
  nor _15176_ (_06845_, _05840_, _06843_);
  nor _15177_ (_06846_, _06845_, _06844_);
  and _15178_ (_06847_, _06846_, _05656_);
  not _15179_ (_06848_, _06847_);
  nor _15180_ (_06849_, _05879_, _06843_);
  and _15181_ (_06850_, _05879_, _06843_);
  nor _15182_ (_06851_, _06850_, _06849_);
  and _15183_ (_06852_, _06851_, _05844_);
  nor _15184_ (_06853_, _06639_, _06649_);
  and _15185_ (_06854_, _06853_, _05678_);
  nor _15186_ (_06855_, _06853_, _05678_);
  or _15187_ (_06856_, _06855_, _06854_);
  and _15188_ (_06857_, _06856_, _05883_);
  nor _15189_ (_06858_, _05715_, _06631_);
  and _15190_ (_06859_, _05535_, _05909_);
  and _15191_ (_06860_, _05381_, _05907_);
  and _15192_ (_06861_, _06600_, ABINPUT000000[8]);
  or _15193_ (_06862_, _06861_, _06860_);
  or _15194_ (_06863_, _06862_, _06859_);
  nor _15195_ (_06864_, _06863_, _06858_);
  nor _15196_ (_06865_, _05678_, _06598_);
  and _15197_ (_06866_, _06606_, ABINPUT000[8]);
  nor _15198_ (_06867_, _06866_, _06865_);
  and _15199_ (_06868_, _06867_, _05956_);
  and _15200_ (_06869_, _06868_, _06864_);
  not _15201_ (_06870_, _06869_);
  nor _15202_ (_06871_, _06870_, _06857_);
  and _15203_ (_06872_, _06871_, _05949_);
  not _15204_ (_06873_, _06872_);
  nor _15205_ (_06874_, _06873_, _06852_);
  and _15206_ (_06875_, _06874_, _06848_);
  nor _15207_ (_06876_, _06875_, _06842_);
  and _15208_ (_06877_, _05241_, _05172_);
  and _15209_ (_06878_, _06877_, _05256_);
  nor _15210_ (_06879_, _05266_, _05227_);
  and _15211_ (_06880_, _06879_, _05647_);
  and _15212_ (_06881_, _06880_, _06878_);
  and _15213_ (_06882_, _06881_, _06008_);
  and _15214_ (_06883_, _06882_, _05963_);
  not _15215_ (_06884_, _06842_);
  nor _15216_ (_06885_, _06882_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _15217_ (_06886_, _06885_, _06884_);
  nor _15218_ (_06888_, _06886_, _06883_);
  nor _15219_ (_06889_, _06888_, _06876_);
  or _15220_ (_06890_, _06889_, _06836_);
  nor _15221_ (_06891_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _15222_ (_06892_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05663_);
  nor _15223_ (_06893_, _06892_, _06891_);
  nor _15224_ (_06894_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15225_ (_06895_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05699_);
  nor _15226_ (_06896_, _06895_, _06894_);
  not _15227_ (_06897_, _06896_);
  nor _15228_ (_06898_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _15229_ (_06899_, _05390_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _15230_ (_06900_, _06899_, _06898_);
  nand _15231_ (_06901_, _05880_, _05846_);
  nor _15232_ (_06902_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _15233_ (_06904_, _05411_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _15234_ (_06905_, _06904_, _06902_);
  and _15235_ (_06906_, _06905_, _06901_);
  nor _15236_ (_06907_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _15237_ (_06908_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05436_);
  nor _15238_ (_06909_, _06908_, _06907_);
  and _15239_ (_06910_, _06909_, _06906_);
  nor _15240_ (_06911_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _15241_ (_06912_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05455_);
  nor _15242_ (_06913_, _06912_, _06911_);
  and _15243_ (_06914_, _06913_, _06910_);
  and _15244_ (_06915_, _06914_, _06900_);
  nor _15245_ (_06916_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15246_ (_06917_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05739_);
  nor _15247_ (_06918_, _06917_, _06916_);
  nor _15248_ (_06919_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15249_ (_06920_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05317_);
  nor _15250_ (_06921_, _06920_, _06919_);
  and _15251_ (_06922_, _06921_, _06918_);
  nand _15252_ (_06923_, _06922_, _06915_);
  or _15253_ (_06924_, _06923_, _06897_);
  nor _15254_ (_06925_, _06924_, _06893_);
  and _15255_ (_06926_, _06924_, _06893_);
  or _15256_ (_06927_, _06926_, _06925_);
  and _15257_ (_06928_, _06927_, _05844_);
  and _15258_ (_06929_, _05768_, _05382_);
  not _15259_ (_06930_, _06929_);
  nand _15260_ (_06931_, _05495_, _05382_);
  nor _15261_ (_06932_, _05942_, _05678_);
  and _15262_ (_06933_, _06932_, _05584_);
  and _15263_ (_06934_, _06933_, _05809_);
  and _15264_ (_06935_, _06934_, _05799_);
  and _15265_ (_06936_, _06935_, _05830_);
  or _15266_ (_06937_, _06936_, _05381_);
  and _15267_ (_06938_, _06937_, _06931_);
  and _15268_ (_06939_, _06938_, _06930_);
  and _15269_ (_06940_, _05678_, _05581_);
  and _15270_ (_06941_, _06940_, _05938_);
  and _15271_ (_06942_, _06941_, _05807_);
  and _15272_ (_06943_, _06942_, _05532_);
  and _15273_ (_06944_, _06943_, _05795_);
  and _15274_ (_06945_, _06944_, _05495_);
  and _15275_ (_06946_, _06945_, _05768_);
  nor _15276_ (_06947_, _06946_, _05382_);
  not _15277_ (_06948_, _06947_);
  and _15278_ (_06949_, _06948_, _06939_);
  and _15279_ (_06950_, _05724_, _05382_);
  nor _15280_ (_06951_, _06950_, _06218_);
  and _15281_ (_06952_, _06951_, _06949_);
  or _15282_ (_06953_, _06952_, _05685_);
  nand _15283_ (_06954_, _06952_, _05685_);
  and _15284_ (_06955_, _06954_, _06953_);
  and _15285_ (_06956_, _06955_, _05481_);
  nor _15286_ (_06958_, _05678_, _05382_);
  nor _15287_ (_06959_, _05684_, _05381_);
  or _15288_ (_06961_, _06959_, _06958_);
  and _15289_ (_06963_, _06961_, _05509_);
  nor _15290_ (_06964_, _05404_, _05893_);
  nor _15291_ (_06965_, _05684_, _06598_);
  and _15292_ (_06967_, _06600_, ABINPUT000000[16]);
  and _15293_ (_06968_, _06606_, ABINPUT000[16]);
  or _15294_ (_06969_, _06968_, _06967_);
  or _15295_ (_06970_, _06969_, _06965_);
  or _15296_ (_06972_, _06970_, _06964_);
  or _15297_ (_06973_, _06972_, _06963_);
  or _15298_ (_06974_, _06973_, _06956_);
  or _15299_ (_06975_, _06974_, _06928_);
  nand _15300_ (_06976_, _06975_, _06836_);
  nand _15301_ (_06977_, _06976_, _06890_);
  and _15302_ (_05329_, _06977_, _05141_);
  and _15303_ (_06978_, _06293_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and _15304_ (_06979_, _06771_, _06546_);
  and _15305_ (_06980_, _06979_, _06450_);
  and _15306_ (_06981_, _06760_, _06570_);
  and _15307_ (_06982_, _06772_, _06449_);
  or _15308_ (_06983_, _06982_, _06981_);
  or _15309_ (_06985_, _06983_, _06980_);
  or _15310_ (_06986_, _06756_, _06571_);
  or _15311_ (_06987_, _06986_, _06784_);
  and _15312_ (_06988_, _06778_, _06546_);
  or _15313_ (_06989_, _06988_, _06779_);
  and _15314_ (_06990_, _06782_, _06544_);
  or _15315_ (_06992_, _06990_, _06989_);
  and _15316_ (_06993_, _06767_, _06544_);
  and _15317_ (_06994_, _06760_, _06547_);
  and _15318_ (_06995_, _06450_, _06417_);
  and _15319_ (_06996_, _06995_, _06545_);
  and _15320_ (_06997_, _06996_, _06474_);
  or _15321_ (_06998_, _06997_, _06994_);
  or _15322_ (_06999_, _06998_, _06993_);
  or _15323_ (_07000_, _06999_, _06992_);
  or _15324_ (_07001_, _07000_, _06987_);
  or _15325_ (_07002_, _07001_, _06985_);
  and _15326_ (_07003_, _07002_, _06296_);
  or _15327_ (_05340_, _07003_, _06978_);
  and _15328_ (_07004_, _06269_, _05143_);
  and _15329_ (_07005_, _07004_, _06815_);
  not _15330_ (_07006_, _06497_);
  nor _15331_ (_07007_, _06524_, _06472_);
  and _15332_ (_07008_, _07007_, _07006_);
  not _15333_ (_07009_, _06415_);
  nor _15334_ (_07010_, _07009_, _06389_);
  and _15335_ (_07011_, _07010_, _06337_);
  and _15336_ (_07012_, _07011_, _06363_);
  and _15337_ (_07013_, _07012_, _07008_);
  not _15338_ (_07014_, _06472_);
  nor _15339_ (_07015_, _06524_, _07014_);
  and _15340_ (_07016_, _07015_, _06497_);
  not _15341_ (_07017_, _06363_);
  and _15342_ (_07018_, _07011_, _07017_);
  and _15343_ (_07019_, _07018_, _07016_);
  nor _15344_ (_07020_, _07009_, _06337_);
  and _15345_ (_07021_, _07020_, _06389_);
  and _15346_ (_07022_, _07021_, _07017_);
  not _15347_ (_07023_, _06447_);
  and _15348_ (_07025_, _07007_, _07023_);
  and _15349_ (_07026_, _07025_, _07022_);
  or _15350_ (_07028_, _07026_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _15351_ (_07029_, _07028_, _07019_);
  or _15352_ (_07030_, _07029_, _07013_);
  and _15353_ (_07031_, _07030_, _07005_);
  nor _15354_ (_07032_, _07004_, _06815_);
  or _15355_ (_07033_, _07032_, rst);
  or _15356_ (_05369_, _07033_, _07031_);
  nor _15357_ (_07034_, _06993_, _06548_);
  and _15358_ (_07035_, _06760_, _06553_);
  or _15359_ (_07036_, _06981_, _07035_);
  and _15360_ (_07037_, _06565_, _06535_);
  nor _15361_ (_07039_, _07037_, _07036_);
  nand _15362_ (_07040_, _07039_, _07034_);
  and _15363_ (_07041_, _06527_, _06449_);
  and _15364_ (_07042_, _07041_, _06760_);
  or _15365_ (_07043_, _07042_, _06799_);
  and _15366_ (_07044_, _06550_, _06546_);
  or _15367_ (_07045_, _07044_, _07043_);
  or _15368_ (_07046_, _07045_, _06819_);
  and _15369_ (_07047_, _06544_, _06765_);
  or _15370_ (_07048_, _07047_, _06994_);
  nand _15371_ (_07049_, _06535_, _06365_);
  not _15372_ (_07050_, _06570_);
  or _15373_ (_07051_, _07050_, _07049_);
  nand _15374_ (_07052_, _06757_, _06760_);
  and _15375_ (_07053_, _06574_, _06450_);
  nand _15376_ (_07054_, _07053_, _06535_);
  and _15377_ (_07055_, _07054_, _07052_);
  nand _15378_ (_07056_, _07055_, _07051_);
  or _15379_ (_07057_, _07056_, _07048_);
  or _15380_ (_07058_, _07057_, _07046_);
  or _15381_ (_07059_, _07058_, _07040_);
  or _15382_ (_07060_, _06997_, _06979_);
  and _15383_ (_07062_, _06778_, _06527_);
  and _15384_ (_07063_, _06995_, _06766_);
  or _15385_ (_07064_, _07063_, _07062_);
  or _15386_ (_07065_, _07064_, _07060_);
  or _15387_ (_07066_, _07065_, _06780_);
  and _15388_ (_07067_, _06782_, _06771_);
  and _15389_ (_07068_, _06449_, _06418_);
  and _15390_ (_07069_, _07068_, _06770_);
  and _15391_ (_07070_, _07069_, _06527_);
  or _15392_ (_07071_, _07070_, _06772_);
  or _15393_ (_07072_, _07071_, _07067_);
  and _15394_ (_07073_, _06564_, _06535_);
  and _15395_ (_07074_, _06807_, _06770_);
  and _15396_ (_07076_, _07074_, _06540_);
  or _15397_ (_07077_, _07076_, _07073_);
  and _15398_ (_07078_, _06995_, _06540_);
  or _15399_ (_07079_, _07078_, _06818_);
  or _15400_ (_07080_, _07079_, _07077_);
  or _15401_ (_07081_, _07080_, _07072_);
  or _15402_ (_07083_, _07081_, _07066_);
  or _15403_ (_07084_, _07083_, _07059_);
  and _15404_ (_07085_, _07084_, _06271_);
  and _15405_ (_07086_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.wr );
  and _15406_ (_07087_, \oc8051_top_1.oc8051_decoder1.state [1], _05143_);
  and _15407_ (_07088_, _07087_, _06815_);
  and _15408_ (_07089_, _07088_, _06820_);
  or _15409_ (_07090_, _07089_, _06798_);
  and _15410_ (_07091_, _07088_, _06554_);
  or _15411_ (_07092_, _07091_, _07090_);
  or _15412_ (_07093_, _07092_, _07086_);
  or _15413_ (_07094_, _07093_, _07085_);
  and _15414_ (_05451_, _07094_, _05141_);
  not _15415_ (_07096_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor _15416_ (_07097_, _05291_, _07096_);
  and _15417_ (_07099_, _06004_, _05291_);
  or _15418_ (_07100_, _07099_, _05572_);
  or _15419_ (_07101_, _07100_, _07097_);
  or _15420_ (_07102_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _15421_ (_07103_, _07102_, _05141_);
  and _15422_ (_05468_, _07103_, _07101_);
  or _15423_ (_07104_, _06556_, _06765_);
  and _15424_ (_07105_, _06755_, _06556_);
  or _15425_ (_07106_, _07105_, _06773_);
  and _15426_ (_07107_, _07106_, _07104_);
  and _15427_ (_07108_, _06765_, _06420_);
  and _15428_ (_07109_, _06760_, _06765_);
  or _15429_ (_07110_, _07109_, _07108_);
  or _15430_ (_07111_, _07110_, _07107_);
  and _15431_ (_07112_, _07111_, _06271_);
  and _15432_ (_07113_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _15433_ (_07114_, _06796_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _15434_ (_07115_, _07114_, _07113_);
  or _15435_ (_07116_, _07115_, _07112_);
  and _15436_ (_05502_, _07116_, _05141_);
  not _15437_ (_07117_, _06270_);
  or _15438_ (_07118_, _06337_, _07117_);
  or _15439_ (_07119_, _06270_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _15440_ (_07120_, _07119_, _05141_);
  and _15441_ (_05558_, _07120_, _07118_);
  nor _15442_ (_05596_, _06472_, rst);
  nor _15443_ (_07121_, _06271_, _05660_);
  nor _15444_ (_07123_, _06308_, _06459_);
  nor _15445_ (_07124_, _06314_, _06462_);
  nor _15446_ (_07125_, _07124_, _07123_);
  and _15447_ (_07126_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _15448_ (_07127_, _06320_, _06464_);
  nor _15449_ (_07128_, _07127_, _07126_);
  and _15450_ (_07129_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _15451_ (_07130_, _06304_, _06457_);
  nor _15452_ (_07131_, _07130_, _07129_);
  and _15453_ (_07132_, _07131_, _07128_);
  and _15454_ (_07133_, _07132_, _07125_);
  and _15455_ (_07134_, _06271_, _06317_);
  not _15456_ (_07135_, _07134_);
  nor _15457_ (_07136_, _07135_, _07133_);
  nor _15458_ (_07137_, _07136_, _07121_);
  nor _15459_ (_05599_, _07137_, rst);
  not _15460_ (_07138_, _06619_);
  not _15461_ (_07139_, _06918_);
  nand _15462_ (_07140_, _06921_, _06915_);
  nand _15463_ (_07141_, _07140_, _07139_);
  or _15464_ (_07142_, _07140_, _07139_);
  and _15465_ (_07143_, _07142_, _05844_);
  and _15466_ (_07144_, _07143_, _07141_);
  nor _15467_ (_07145_, _06945_, _05382_);
  not _15468_ (_07146_, _07145_);
  and _15469_ (_07147_, _07146_, _06938_);
  and _15470_ (_07148_, _07147_, _05768_);
  nor _15471_ (_07149_, _07147_, _05768_);
  or _15472_ (_07150_, _07149_, _07148_);
  and _15473_ (_07151_, _07150_, _05481_);
  nand _15474_ (_07152_, _05758_, _05381_);
  nor _15475_ (_07153_, _06929_, _05510_);
  and _15476_ (_07154_, _07153_, _07152_);
  and _15477_ (_07155_, _05537_, _05892_);
  nor _15478_ (_07156_, _05768_, _06598_);
  and _15479_ (_07157_, _06600_, ABINPUT000000[14]);
  and _15480_ (_07158_, _06606_, ABINPUT000[14]);
  or _15481_ (_07159_, _07158_, _07157_);
  or _15482_ (_07161_, _07159_, _07156_);
  or _15483_ (_07162_, _07161_, _07155_);
  or _15484_ (_07163_, _07162_, _07154_);
  or _15485_ (_07164_, _07163_, _07151_);
  or _15486_ (_07166_, _07164_, _07144_);
  or _15487_ (_07167_, _07166_, _07138_);
  and _15488_ (_07168_, _06621_, _06032_);
  not _15489_ (_07169_, _07168_);
  nor _15490_ (_07170_, _05836_, _05786_);
  nor _15491_ (_07171_, _07170_, _05837_);
  nor _15492_ (_07172_, _07171_, _05657_);
  not _15493_ (_07173_, _07172_);
  and _15494_ (_07174_, _05869_, _05865_);
  not _15495_ (_07175_, _07174_);
  and _15496_ (_07176_, _05870_, _05844_);
  and _15497_ (_07177_, _07176_, _07175_);
  nor _15498_ (_07178_, _06642_, _06645_);
  nor _15499_ (_07179_, _07178_, _06640_);
  and _15500_ (_07180_, _07178_, _06640_);
  or _15501_ (_07181_, _07180_, _06591_);
  nor _15502_ (_07182_, _07181_, _07179_);
  nor _15503_ (_07183_, _06631_, _05346_);
  and _15504_ (_07184_, _06600_, ABINPUT000000[6]);
  and _15505_ (_07185_, _06606_, ABINPUT000[6]);
  nor _15506_ (_07186_, _07185_, _07184_);
  not _15507_ (_07187_, _07186_);
  nor _15508_ (_07188_, _07187_, _07183_);
  nor _15509_ (_07189_, _05758_, _06598_);
  not _15510_ (_07190_, _07189_);
  or _15511_ (_07191_, _05715_, _06603_);
  and _15512_ (_07192_, _07191_, _07190_);
  and _15513_ (_07193_, _07192_, _07188_);
  and _15514_ (_07194_, _07193_, _06002_);
  not _15515_ (_07195_, _07194_);
  nor _15516_ (_07196_, _07195_, _07182_);
  and _15517_ (_07197_, _07196_, _05991_);
  not _15518_ (_07198_, _07197_);
  nor _15519_ (_07199_, _07198_, _07177_);
  and _15520_ (_07200_, _07199_, _07173_);
  nor _15521_ (_07201_, _07200_, _07169_);
  and _15522_ (_07202_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _15523_ (_07203_, _07202_, _06619_);
  or _15524_ (_07204_, _07203_, _07201_);
  and _15525_ (_07205_, _07204_, _05141_);
  and _15526_ (_05687_, _07205_, _07167_);
  or _15527_ (_07207_, _06921_, _06915_);
  and _15528_ (_07208_, _07140_, _05844_);
  and _15529_ (_07209_, _07208_, _07207_);
  nor _15530_ (_07210_, _06944_, _05382_);
  not _15531_ (_07211_, _07210_);
  and _15532_ (_07212_, _07211_, _06937_);
  nand _15533_ (_07213_, _07212_, _05771_);
  or _15534_ (_07214_, _07212_, _05771_);
  and _15535_ (_07215_, _07214_, _07213_);
  and _15536_ (_07216_, _07215_, _05481_);
  nand _15537_ (_07217_, _05381_, _05346_);
  and _15538_ (_07218_, _06931_, _05509_);
  and _15539_ (_07219_, _07218_, _07217_);
  and _15540_ (_07220_, _05535_, _05892_);
  nor _15541_ (_07221_, _05495_, _06598_);
  and _15542_ (_07222_, _06600_, ABINPUT000000[13]);
  and _15543_ (_07223_, _06606_, ABINPUT000[13]);
  or _15544_ (_07224_, _07223_, _07222_);
  or _15545_ (_07225_, _07224_, _07221_);
  or _15546_ (_07226_, _07225_, _07220_);
  or _15547_ (_07227_, _07226_, _07219_);
  or _15548_ (_07228_, _07227_, _07216_);
  or _15549_ (_07229_, _07228_, _07209_);
  or _15550_ (_07230_, _07229_, _07138_);
  nor _15551_ (_07231_, _05835_, _05498_);
  and _15552_ (_07232_, _05835_, _05498_);
  nor _15553_ (_07233_, _07232_, _07231_);
  and _15554_ (_07234_, _07233_, _05656_);
  not _15555_ (_07235_, _07234_);
  nor _15556_ (_07236_, _05864_, _05498_);
  nor _15557_ (_07237_, _07236_, _05845_);
  and _15558_ (_07238_, _07237_, _05865_);
  nor _15559_ (_07239_, _05887_, _06591_);
  nor _15560_ (_07240_, _07239_, _05355_);
  nor _15561_ (_07241_, _07240_, _05346_);
  not _15562_ (_07242_, _07241_);
  and _15563_ (_07243_, _06637_, _05346_);
  or _15564_ (_07244_, _05758_, _06603_);
  nor _15565_ (_07245_, _05404_, _06631_);
  and _15566_ (_07246_, _06600_, ABINPUT000000[5]);
  and _15567_ (_07248_, _06606_, ABINPUT000[5]);
  nor _15568_ (_07249_, _07248_, _07246_);
  not _15569_ (_07250_, _07249_);
  nor _15570_ (_07251_, _07250_, _07245_);
  and _15571_ (_07252_, _07251_, _07244_);
  not _15572_ (_07253_, _07252_);
  nor _15573_ (_07254_, _07253_, _07243_);
  and _15574_ (_07255_, _07254_, _07242_);
  and _15575_ (_07256_, _07255_, _05521_);
  not _15576_ (_07257_, _07256_);
  nor _15577_ (_07258_, _07257_, _07238_);
  and _15578_ (_07259_, _07258_, _07235_);
  nor _15579_ (_07260_, _07259_, _07169_);
  and _15580_ (_07261_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _15581_ (_07262_, _07261_, _06619_);
  or _15582_ (_07263_, _07262_, _07260_);
  and _15583_ (_07264_, _07263_, _05141_);
  and _15584_ (_05690_, _07264_, _07230_);
  or _15585_ (_07265_, _06923_, _06896_);
  nand _15586_ (_07266_, _06923_, _06896_);
  nand _15587_ (_07267_, _07266_, _07265_);
  nand _15588_ (_07268_, _07267_, _05844_);
  and _15589_ (_07269_, _06949_, _05724_);
  nor _15590_ (_07270_, _06949_, _05724_);
  nor _15591_ (_07271_, _07270_, _07269_);
  nor _15592_ (_07272_, _07271_, _05597_);
  and _15593_ (_07273_, _06606_, ABINPUT000[15]);
  and _15594_ (_07274_, _05715_, _05381_);
  not _15595_ (_07275_, _07274_);
  nor _15596_ (_07276_, _06950_, _05510_);
  and _15597_ (_07278_, _07276_, _07275_);
  nor _15598_ (_07279_, _05469_, _05893_);
  nor _15599_ (_07280_, _05724_, _06598_);
  and _15600_ (_07281_, _06600_, ABINPUT000000[15]);
  or _15601_ (_07282_, _07281_, _07280_);
  or _15602_ (_07283_, _07282_, _07279_);
  or _15603_ (_07284_, _07283_, _07278_);
  nor _15604_ (_07285_, _07284_, _07273_);
  not _15605_ (_07286_, _07285_);
  nor _15606_ (_07287_, _07286_, _07272_);
  nand _15607_ (_07288_, _07287_, _07268_);
  or _15608_ (_07289_, _07288_, _07138_);
  and _15609_ (_07290_, _07168_, _06669_);
  and _15610_ (_07291_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _15611_ (_07292_, _07291_, _06619_);
  or _15612_ (_07293_, _07292_, _07290_);
  and _15613_ (_07294_, _07293_, _05141_);
  and _15614_ (_05698_, _07294_, _07289_);
  or _15615_ (_07295_, _06914_, _06900_);
  nor _15616_ (_07296_, _06915_, _05845_);
  nand _15617_ (_07298_, _07296_, _07295_);
  not _15618_ (_07299_, _05894_);
  or _15619_ (_07300_, _06935_, _05381_);
  nor _15620_ (_07301_, _06943_, _05382_);
  not _15621_ (_07302_, _07301_);
  and _15622_ (_07303_, _07302_, _07300_);
  nor _15623_ (_07304_, _07303_, _05830_);
  and _15624_ (_07305_, _07303_, _05830_);
  or _15625_ (_07306_, _07305_, _05597_);
  nor _15626_ (_07307_, _07306_, _07304_);
  nor _15627_ (_07308_, _05510_, _05404_);
  not _15628_ (_07309_, _07308_);
  nor _15629_ (_07310_, _05795_, _06598_);
  and _15630_ (_07311_, _06600_, ABINPUT000000[12]);
  and _15631_ (_07312_, _06606_, ABINPUT000[12]);
  nor _15632_ (_07313_, _07312_, _07311_);
  not _15633_ (_07314_, _07313_);
  nor _15634_ (_07315_, _07314_, _07310_);
  nand _15635_ (_07316_, _07315_, _07309_);
  nor _15636_ (_07317_, _07316_, _07307_);
  and _15637_ (_07318_, _07317_, _07299_);
  nand _15638_ (_07319_, _07318_, _07298_);
  or _15639_ (_07320_, _07319_, _07138_);
  nor _15640_ (_07321_, _05828_, _05819_);
  nor _15641_ (_07322_, _07321_, _05829_);
  nor _15642_ (_07323_, _07322_, _05657_);
  not _15643_ (_07324_, _07323_);
  nor _15644_ (_07325_, _05859_, _05854_);
  or _15645_ (_07326_, _07325_, _05845_);
  nor _15646_ (_07327_, _07326_, _05860_);
  not _15647_ (_07328_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _15648_ (_07329_, _05470_, _07328_);
  nor _15649_ (_07330_, _07329_, _05405_);
  not _15650_ (_07331_, _07330_);
  and _15651_ (_07332_, _07331_, _07239_);
  nor _15652_ (_07333_, _05404_, _06598_);
  and _15653_ (_07334_, _06600_, ABINPUT000000[4]);
  and _15654_ (_07335_, _06606_, ABINPUT000[4]);
  nor _15655_ (_07336_, _07335_, _07334_);
  not _15656_ (_07337_, _07336_);
  nor _15657_ (_07338_, _07337_, _07333_);
  or _15658_ (_07339_, _06603_, _05346_);
  nor _15659_ (_07340_, _05469_, _06631_);
  not _15660_ (_07341_, _07340_);
  and _15661_ (_07342_, _07341_, _07339_);
  and _15662_ (_07343_, _07342_, _07338_);
  not _15663_ (_07344_, _07343_);
  nor _15664_ (_07345_, _07344_, _07332_);
  and _15665_ (_07346_, _07345_, _06060_);
  and _15666_ (_07347_, _07346_, _06048_);
  not _15667_ (_07348_, _07347_);
  nor _15668_ (_07349_, _07348_, _07327_);
  and _15669_ (_07350_, _07349_, _07324_);
  nand _15670_ (_07351_, _07350_, _07168_);
  or _15671_ (_07352_, _07168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _15672_ (_07353_, _07352_, _07351_);
  or _15673_ (_07354_, _07353_, _06619_);
  and _15674_ (_07355_, _07354_, _05141_);
  and _15675_ (_05707_, _07355_, _07320_);
  or _15676_ (_07356_, _06913_, _06910_);
  nor _15677_ (_07357_, _06914_, _05845_);
  nand _15678_ (_07358_, _07357_, _07356_);
  or _15679_ (_07359_, _06934_, _05381_);
  nor _15680_ (_07360_, _06942_, _05382_);
  not _15681_ (_07361_, _07360_);
  and _15682_ (_07362_, _07361_, _07359_);
  and _15683_ (_07363_, _07362_, _05799_);
  nor _15684_ (_07364_, _07362_, _05799_);
  nor _15685_ (_07365_, _07364_, _07363_);
  and _15686_ (_07366_, _07365_, _05481_);
  nor _15687_ (_07367_, _05715_, _05893_);
  nor _15688_ (_07368_, _05532_, _06598_);
  and _15689_ (_07369_, _06600_, ABINPUT000000[11]);
  or _15690_ (_07370_, _07369_, _07368_);
  nor _15691_ (_07371_, _07370_, _07367_);
  nor _15692_ (_07372_, _05510_, _05469_);
  and _15693_ (_07373_, _06606_, ABINPUT000[11]);
  nor _15694_ (_07374_, _07373_, _07372_);
  and _15695_ (_07375_, _07374_, _07371_);
  not _15696_ (_07376_, _07375_);
  nor _15697_ (_07377_, _07376_, _07366_);
  nand _15698_ (_07378_, _07377_, _07358_);
  or _15699_ (_07379_, _07378_, _07138_);
  or _15700_ (_07380_, _07168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nand _15701_ (_07381_, _07168_, _06617_);
  and _15702_ (_07382_, _07381_, _07380_);
  or _15703_ (_07383_, _07382_, _06619_);
  and _15704_ (_07384_, _07383_, _05141_);
  and _15705_ (_05714_, _07384_, _07379_);
  or _15706_ (_07385_, _06909_, _06906_);
  nor _15707_ (_07386_, _06910_, _05845_);
  nand _15708_ (_07387_, _07386_, _07385_);
  nor _15709_ (_07388_, _06933_, _05381_);
  nor _15710_ (_07389_, _06941_, _05382_);
  nor _15711_ (_07390_, _07389_, _07388_);
  and _15712_ (_07391_, _07390_, _05807_);
  nor _15713_ (_07392_, _07390_, _05807_);
  or _15714_ (_07393_, _07392_, _07391_);
  and _15715_ (_07394_, _07393_, _05481_);
  nor _15716_ (_07395_, _05758_, _05893_);
  and _15717_ (_07396_, _05809_, _05355_);
  and _15718_ (_07397_, _06600_, ABINPUT000000[10]);
  or _15719_ (_07398_, _07397_, _07396_);
  nor _15720_ (_07399_, _07398_, _07395_);
  and _15721_ (_07400_, _05509_, _05537_);
  and _15722_ (_07401_, _06606_, ABINPUT000[10]);
  nor _15723_ (_07402_, _07401_, _07400_);
  and _15724_ (_07403_, _07402_, _07399_);
  not _15725_ (_07404_, _07403_);
  nor _15726_ (_07405_, _07404_, _07394_);
  nand _15727_ (_07406_, _07405_, _07387_);
  or _15728_ (_07407_, _07406_, _07138_);
  or _15729_ (_07408_, _07168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor _15730_ (_07409_, _05826_, _05824_);
  nor _15731_ (_07410_, _07409_, _05827_);
  nor _15732_ (_07411_, _07410_, _05657_);
  not _15733_ (_07412_, _07411_);
  or _15734_ (_07413_, _05469_, _06603_);
  and _15735_ (_07414_, _06600_, ABINPUT000000[2]);
  and _15736_ (_07415_, _06606_, ABINPUT000[2]);
  nor _15737_ (_07416_, _07415_, _07414_);
  and _15738_ (_07417_, _07416_, _07413_);
  and _15739_ (_07418_, _05535_, _05367_);
  and _15740_ (_07419_, _05537_, _05355_);
  nor _15741_ (_07420_, _07419_, _07418_);
  and _15742_ (_07421_, _07420_, _07417_);
  and _15743_ (_07422_, _07421_, _06177_);
  and _15744_ (_07423_, _06592_, _05537_);
  nor _15745_ (_07424_, _07423_, _06593_);
  nor _15746_ (_07425_, _07424_, _06591_);
  and _15747_ (_07426_, _06167_, _05590_);
  or _15748_ (_07427_, _07426_, _05848_);
  and _15749_ (_07428_, _07427_, _05855_);
  nor _15750_ (_07429_, _07427_, _05855_);
  or _15751_ (_07430_, _07429_, _07428_);
  and _15752_ (_07431_, _07430_, _05844_);
  nor _15753_ (_07432_, _07431_, _07425_);
  and _15754_ (_07433_, _07432_, _07422_);
  and _15755_ (_07434_, _07433_, _07412_);
  nand _15756_ (_07435_, _07434_, _07168_);
  and _15757_ (_07436_, _07435_, _07408_);
  or _15758_ (_07437_, _07436_, _06619_);
  and _15759_ (_07438_, _07437_, _05141_);
  and _15760_ (_05717_, _07438_, _07407_);
  or _15761_ (_07439_, _06905_, _06901_);
  nor _15762_ (_07440_, _06906_, _05845_);
  nand _15763_ (_07441_, _07440_, _07439_);
  nor _15764_ (_07442_, _05930_, _06958_);
  and _15765_ (_07444_, _07442_, _05944_);
  nor _15766_ (_07445_, _07444_, _05584_);
  and _15767_ (_07447_, _07444_, _05584_);
  nor _15768_ (_07448_, _07447_, _07445_);
  and _15769_ (_07450_, _07448_, _05481_);
  nor _15770_ (_07451_, _05893_, _05346_);
  nor _15771_ (_07452_, _05581_, _06598_);
  and _15772_ (_07453_, _06600_, ABINPUT000000[9]);
  or _15773_ (_07455_, _07453_, _07452_);
  nor _15774_ (_07456_, _07455_, _07451_);
  and _15775_ (_07458_, _05509_, _05535_);
  and _15776_ (_07459_, _06606_, ABINPUT000[9]);
  nor _15777_ (_07461_, _07459_, _07458_);
  and _15778_ (_07462_, _07461_, _07456_);
  not _15779_ (_07463_, _07462_);
  nor _15780_ (_07464_, _07463_, _07450_);
  nand _15781_ (_07466_, _07464_, _07441_);
  or _15782_ (_07467_, _07466_, _07138_);
  or _15783_ (_07468_, _07168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _15784_ (_07469_, _05883_, _05535_);
  and _15785_ (_07471_, _05936_, _05896_);
  nor _15786_ (_07472_, _07471_, _07469_);
  and _15787_ (_07473_, _05535_, _05355_);
  not _15788_ (_07474_, _07473_);
  and _15789_ (_07476_, _06606_, ABINPUT000[1]);
  and _15790_ (_07478_, _05381_, _05892_);
  and _15791_ (_07479_, _06600_, ABINPUT000000[1]);
  or _15792_ (_07480_, _07479_, _07478_);
  nor _15793_ (_07481_, _07480_, _07476_);
  and _15794_ (_07482_, _07481_, _07474_);
  and _15795_ (_07483_, _07482_, _07472_);
  and _15796_ (_07484_, _07483_, _05588_);
  nor _15797_ (_07485_, _05825_, _05381_);
  nor _15798_ (_07486_, _07485_, _05855_);
  not _15799_ (_07487_, _07486_);
  nor _15800_ (_07488_, _05844_, _05656_);
  nor _15801_ (_07489_, _07488_, _07487_);
  or _15802_ (_07490_, _05446_, _06603_);
  and _15803_ (_07491_, _07490_, _05600_);
  and _15804_ (_07492_, _07491_, _05594_);
  not _15805_ (_07494_, _07492_);
  nor _15806_ (_07495_, _07494_, _07489_);
  and _15807_ (_07496_, _07495_, _07484_);
  nand _15808_ (_07497_, _07496_, _07168_);
  and _15809_ (_07498_, _07497_, _07468_);
  or _15810_ (_07499_, _07498_, _06619_);
  and _15811_ (_07500_, _07499_, _05141_);
  and _15812_ (_05720_, _07500_, _07467_);
  and _15813_ (_05726_, _06363_, _05141_);
  and _15814_ (_05729_, _06337_, _05141_);
  and _15815_ (_05732_, _06389_, _05141_);
  nor _15816_ (_05735_, _06415_, rst);
  and _15817_ (_05738_, _06447_, _05141_);
  and _15818_ (_05741_, _06497_, _05141_);
  and _15819_ (_05744_, _06524_, _05141_);
  nor _15820_ (_07501_, _06271_, _05731_);
  nor _15821_ (_07502_, _06308_, _06487_);
  nor _15822_ (_07503_, _06314_, _06484_);
  nor _15823_ (_07504_, _07503_, _07502_);
  and _15824_ (_07505_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _15825_ (_07506_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _15826_ (_07507_, _07506_, _07505_);
  nor _15827_ (_07508_, _06304_, _06482_);
  nor _15828_ (_07509_, _06320_, _06489_);
  nor _15829_ (_07510_, _07509_, _07508_);
  and _15830_ (_07511_, _07510_, _07507_);
  and _15831_ (_07512_, _07511_, _07504_);
  nor _15832_ (_07513_, _07512_, _07135_);
  nor _15833_ (_07514_, _07513_, _07501_);
  nor _15834_ (_05756_, _07514_, rst);
  nor _15835_ (_07515_, _06271_, _05408_);
  not _15836_ (_07516_, _06271_);
  and _15837_ (_07517_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _15838_ (_07518_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor _15839_ (_07519_, _06320_, _06343_);
  nor _15840_ (_07520_, _07519_, _07518_);
  nor _15841_ (_07521_, _06308_, _06347_);
  and _15842_ (_07522_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _15843_ (_07523_, _07522_, _07521_);
  not _15844_ (_07524_, _06304_);
  and _15845_ (_07525_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _15846_ (_07526_, _06314_, _06351_);
  nor _15847_ (_07527_, _07526_, _07525_);
  and _15848_ (_07528_, _07527_, _07523_);
  and _15849_ (_07529_, _07528_, _07520_);
  nor _15850_ (_07530_, _07529_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15851_ (_07531_, _07530_, _07517_);
  nor _15852_ (_07532_, _07531_, _07516_);
  nor _15853_ (_07533_, _07532_, _07515_);
  nor _15854_ (_05760_, _07533_, rst);
  nor _15855_ (_07534_, _06271_, _05449_);
  and _15856_ (_07535_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15857_ (_07536_, _06308_, _06379_);
  nor _15858_ (_07537_, _06320_, _06374_);
  nor _15859_ (_07538_, _07537_, _07536_);
  and _15860_ (_07539_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor _15861_ (_07540_, _06314_, _06376_);
  nor _15862_ (_07541_, _07540_, _07539_);
  and _15863_ (_07542_, _07541_, _07538_);
  and _15864_ (_07543_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _15865_ (_07544_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _15866_ (_07545_, _07544_, _07543_);
  and _15867_ (_07546_, _07545_, _07542_);
  nor _15868_ (_07547_, _07546_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15869_ (_07548_, _07547_, _07535_);
  nor _15870_ (_07549_, _07548_, _07516_);
  nor _15871_ (_07550_, _07549_, _07534_);
  nor _15872_ (_05764_, _07550_, rst);
  and _15873_ (_07551_, _07516_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _15874_ (_07552_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _15875_ (_07554_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _15876_ (_07555_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _15877_ (_07556_, _07555_, _07554_);
  and _15878_ (_07557_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor _15879_ (_07559_, _06314_, _06403_);
  nor _15880_ (_07560_, _07559_, _07557_);
  nor _15881_ (_07561_, _06320_, _06395_);
  nor _15882_ (_07563_, _06308_, _06399_);
  nor _15883_ (_07564_, _07563_, _07561_);
  and _15884_ (_07566_, _07564_, _07560_);
  and _15885_ (_07567_, _07566_, _07556_);
  nor _15886_ (_07568_, _07567_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15887_ (_07570_, _07568_, _07552_);
  nor _15888_ (_07571_, _07570_, _07516_);
  nor _15889_ (_07572_, _07571_, _07551_);
  nor _15890_ (_05767_, _07572_, rst);
  nor _15891_ (_07574_, _06271_, _05307_);
  and _15892_ (_07576_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _15893_ (_07577_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor _15894_ (_07579_, _06320_, _06429_);
  nor _15895_ (_07580_, _07579_, _07577_);
  not _15896_ (_07581_, _06308_);
  and _15897_ (_07582_, _07581_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _15898_ (_07583_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _15899_ (_07584_, _07583_, _07582_);
  and _15900_ (_07585_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor _15901_ (_07586_, _06314_, _06427_);
  nor _15902_ (_07587_, _07586_, _07585_);
  and _15903_ (_07588_, _07587_, _07584_);
  and _15904_ (_07589_, _07588_, _07580_);
  nor _15905_ (_07590_, _07589_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15906_ (_07591_, _07590_, _07576_);
  nor _15907_ (_07592_, _07591_, _07516_);
  nor _15908_ (_07593_, _07592_, _07574_);
  nor _15909_ (_05770_, _07593_, rst);
  nand _15910_ (_07594_, _07200_, _06624_);
  or _15911_ (_07595_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _15912_ (_07596_, _07595_, _05141_);
  and _15913_ (_05780_, _07596_, _07594_);
  or _15914_ (_07597_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand _15915_ (_07598_, _07434_, _06624_);
  and _15916_ (_07599_, _07598_, _05141_);
  and _15917_ (_05783_, _07599_, _07597_);
  or _15918_ (_07600_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _15919_ (_07601_, _07496_, _06624_);
  and _15920_ (_07602_, _07601_, _05141_);
  and _15921_ (_05790_, _07602_, _07600_);
  nand _15922_ (_07603_, _07259_, _06624_);
  or _15923_ (_07604_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _15924_ (_07605_, _07604_, _05141_);
  and _15925_ (_05793_, _07605_, _07603_);
  and _15926_ (_07606_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _15927_ (_07607_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _15928_ (_07608_, pc_log_change, _07607_);
  or _15929_ (_07609_, _07608_, _07606_);
  and _15930_ (_05932_, _07609_, _05141_);
  nor _15931_ (_07610_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not _15932_ (_07611_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _15933_ (_07612_, _07611_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor _15934_ (_07613_, _07612_, _07610_);
  not _15935_ (_07614_, \oc8051_symbolic_cxrom1.regvalid [13]);
  not _15936_ (_07615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _15937_ (_07617_, _06307_, _06302_);
  nor _15938_ (_07618_, _07617_, _07516_);
  nor _15939_ (_07619_, _07618_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _15940_ (_07620_, _07619_, _07615_);
  nor _15941_ (_07621_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _15942_ (_07622_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _15943_ (_07623_, _07622_, _07621_);
  nor _15944_ (_07624_, _07623_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _15945_ (_07625_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _07611_);
  nor _15946_ (_07626_, _07625_, _07624_);
  and _15947_ (_07627_, _07626_, _07614_);
  nor _15948_ (_07628_, _07626_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _15949_ (_07629_, _07628_, _07627_);
  not _15950_ (_07630_, _07629_);
  nor _15951_ (_07631_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _15952_ (_07632_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _07611_);
  nor _15953_ (_07633_, _07632_, _07631_);
  not _15954_ (_07634_, _07633_);
  and _15955_ (_07635_, _07619_, _07615_);
  nor _15956_ (_07636_, _07635_, _07620_);
  nor _15957_ (_07637_, _07636_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _15958_ (_07638_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _07611_);
  nor _15959_ (_07639_, _07638_, _07637_);
  and _15960_ (_07640_, _07639_, _07634_);
  nand _15961_ (_07641_, _07640_, _07630_);
  and _15962_ (_07642_, _07641_, _07613_);
  nor _15963_ (_07643_, _07639_, _07634_);
  not _15964_ (_07644_, _07643_);
  not _15965_ (_07645_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _15966_ (_07646_, _07626_, _07645_);
  and _15967_ (_07647_, _07626_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _15968_ (_07648_, _07647_, _07646_);
  nor _15969_ (_07649_, _07648_, _07644_);
  and _15970_ (_07650_, _07639_, _07633_);
  not _15971_ (_07651_, _07650_);
  not _15972_ (_07652_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _15973_ (_07653_, _07626_, _07652_);
  and _15974_ (_07654_, _07626_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _15975_ (_07656_, _07654_, _07653_);
  nor _15976_ (_07657_, _07656_, _07651_);
  nor _15977_ (_07659_, _07657_, _07649_);
  not _15978_ (_07661_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _15979_ (_07662_, _07626_, _07661_);
  nor _15980_ (_07663_, _07626_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _15981_ (_07665_, _07663_);
  nor _15982_ (_07666_, _07639_, _07633_);
  nand _15983_ (_07668_, _07666_, _07665_);
  or _15984_ (_07669_, _07668_, _07662_);
  and _15985_ (_07671_, _07669_, _07659_);
  and _15986_ (_07673_, _07671_, _07642_);
  and _15987_ (_07674_, _07626_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _15988_ (_07675_, _07674_, _07643_);
  not _15989_ (_07676_, _07626_);
  and _15990_ (_07678_, _07643_, _07676_);
  and _15991_ (_07679_, _07678_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _15992_ (_07681_, _07679_, _07613_);
  or _15993_ (_07683_, _07681_, _07675_);
  not _15994_ (_07684_, _07666_);
  and _15995_ (_07685_, _07626_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not _15996_ (_07686_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _15997_ (_07688_, _07626_, _07686_);
  nor _15998_ (_07689_, _07688_, _07685_);
  nor _15999_ (_07690_, _07689_, _07684_);
  not _16000_ (_07691_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _16001_ (_07692_, _07626_, _07691_);
  nor _16002_ (_07693_, _07626_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _16003_ (_07694_, _07693_, _07692_);
  nor _16004_ (_07695_, _07694_, _07651_);
  not _16005_ (_07696_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _16006_ (_07697_, _07626_, _07696_);
  nor _16007_ (_07698_, _07626_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _16008_ (_07699_, _07698_, _07697_);
  not _16009_ (_07700_, _07699_);
  and _16010_ (_07701_, _07700_, _07640_);
  or _16011_ (_07702_, _07701_, _07695_);
  or _16012_ (_07703_, _07702_, _07690_);
  nor _16013_ (_07704_, _07703_, _07683_);
  nor _16014_ (_07705_, _07704_, _07673_);
  not _16015_ (_07706_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _16016_ (_07707_, _07613_, _07706_);
  or _16017_ (_07708_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _16018_ (_07709_, _07708_, _07707_);
  and _16019_ (_07710_, _07709_, _07650_);
  not _16020_ (_07711_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _16021_ (_07712_, _07613_, _07711_);
  or _16022_ (_07713_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _16023_ (_07714_, _07713_, _07712_);
  and _16024_ (_07715_, _07714_, _07643_);
  or _16025_ (_07716_, _07715_, _07710_);
  not _16026_ (_07717_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _16027_ (_07718_, _07613_, _07717_);
  or _16028_ (_07719_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _16029_ (_07720_, _07719_, _07718_);
  and _16030_ (_07721_, _07720_, _07640_);
  not _16031_ (_07722_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _16032_ (_07723_, _07613_, _07722_);
  or _16033_ (_07724_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _16034_ (_07725_, _07724_, _07723_);
  and _16035_ (_07726_, _07725_, _07666_);
  or _16036_ (_07727_, _07726_, _07721_);
  or _16037_ (_07728_, _07727_, _07716_);
  and _16038_ (_07729_, _07728_, _07626_);
  not _16039_ (_07730_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _16040_ (_07731_, _07613_, _07730_);
  or _16041_ (_07732_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _16042_ (_07733_, _07732_, _07731_);
  and _16043_ (_07734_, _07733_, _07643_);
  not _16044_ (_07735_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _16045_ (_07736_, _07613_, _07735_);
  or _16046_ (_07737_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _16047_ (_07738_, _07737_, _07736_);
  and _16048_ (_07739_, _07738_, _07650_);
  or _16049_ (_07740_, _07739_, _07734_);
  not _16050_ (_07741_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _16051_ (_07742_, _07613_, _07741_);
  or _16052_ (_07743_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _16053_ (_07744_, _07743_, _07742_);
  and _16054_ (_07745_, _07744_, _07640_);
  not _16055_ (_07746_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _16056_ (_07747_, _07613_, _07746_);
  or _16057_ (_07748_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _16058_ (_07750_, _07748_, _07747_);
  and _16059_ (_07751_, _07750_, _07666_);
  or _16060_ (_07752_, _07751_, _07745_);
  or _16061_ (_07753_, _07752_, _07740_);
  and _16062_ (_07754_, _07753_, _07676_);
  or _16063_ (_07756_, _07754_, _07729_);
  and _16064_ (_07757_, _07756_, _07705_);
  not _16065_ (_07758_, _07705_);
  and _16066_ (_07759_, _07758_, word_in[7]);
  or _16067_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _07759_, _07757_);
  nor _16068_ (_07761_, _07633_, _07613_);
  not _16069_ (_07763_, _07761_);
  and _16070_ (_07765_, _07633_, _07613_);
  and _16071_ (_07766_, _07765_, _07639_);
  nor _16072_ (_07768_, _07765_, _07639_);
  nor _16073_ (_07769_, _07768_, _07766_);
  not _16074_ (_07771_, _07769_);
  nor _16075_ (_07772_, _07771_, _07629_);
  not _16076_ (_07773_, _07766_);
  and _16077_ (_07774_, _07773_, _07626_);
  not _16078_ (_07776_, _07639_);
  nor _16079_ (_07777_, _07776_, _07626_);
  and _16080_ (_07779_, _07777_, _07765_);
  nor _16081_ (_07780_, _07779_, _07774_);
  and _16082_ (_07781_, _07780_, _07771_);
  and _16083_ (_07782_, _07781_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _16084_ (_07783_, _07780_, _07769_);
  and _16085_ (_07784_, _07783_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _16086_ (_07785_, _07784_, _07782_);
  nor _16087_ (_07786_, _07785_, _07772_);
  nor _16088_ (_07787_, _07786_, _07763_);
  and _16089_ (_07788_, _07634_, _07613_);
  not _16090_ (_07789_, _07788_);
  nor _16091_ (_07790_, _07771_, _07694_);
  and _16092_ (_07791_, _07781_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _16093_ (_07792_, _07783_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _16094_ (_07793_, _07792_, _07791_);
  nor _16095_ (_07794_, _07793_, _07790_);
  nor _16096_ (_07795_, _07794_, _07789_);
  nor _16097_ (_07796_, _07795_, _07787_);
  not _16098_ (_07797_, _07613_);
  and _16099_ (_07798_, _07633_, _07797_);
  not _16100_ (_07799_, _07798_);
  nor _16101_ (_07800_, _07771_, _07656_);
  and _16102_ (_07801_, _07781_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _16103_ (_07802_, _07783_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _16104_ (_07803_, _07802_, _07801_);
  nor _16105_ (_07804_, _07803_, _07800_);
  nor _16106_ (_07805_, _07804_, _07799_);
  not _16107_ (_07806_, _07765_);
  and _16108_ (_07807_, _07769_, _07676_);
  and _16109_ (_07808_, _07807_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _16110_ (_07809_, _07783_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16111_ (_07810_, _07781_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _16112_ (_07811_, _07769_, _07626_);
  and _16113_ (_07812_, _07811_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _16114_ (_07813_, _07812_, _07810_);
  or _16115_ (_07814_, _07813_, _07809_);
  nor _16116_ (_07815_, _07814_, _07808_);
  nor _16117_ (_07817_, _07815_, _07806_);
  nor _16118_ (_07818_, _07817_, _07805_);
  and _16119_ (_07819_, _07818_, _07796_);
  or _16120_ (_07820_, _07761_, _07765_);
  not _16121_ (_07821_, _07820_);
  not _16122_ (_07822_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _16123_ (_07823_, _07613_, _07822_);
  or _16124_ (_07824_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _16125_ (_07825_, _07824_, _07823_);
  and _16126_ (_07826_, _07825_, _07821_);
  not _16127_ (_07827_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _16128_ (_07828_, _07613_, _07827_);
  or _16129_ (_07829_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _16130_ (_07830_, _07829_, _07828_);
  and _16131_ (_07831_, _07830_, _07820_);
  or _16132_ (_07832_, _07831_, _07826_);
  and _16133_ (_07833_, _07832_, _07783_);
  not _16134_ (_07834_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _16135_ (_07835_, _07613_, _07834_);
  or _16136_ (_07836_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _16137_ (_07837_, _07836_, _07835_);
  and _16138_ (_07838_, _07837_, _07821_);
  not _16139_ (_07839_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _16140_ (_07840_, _07613_, _07839_);
  or _16141_ (_07841_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _16142_ (_07842_, _07841_, _07840_);
  and _16143_ (_07843_, _07842_, _07820_);
  or _16144_ (_07844_, _07843_, _07838_);
  and _16145_ (_07845_, _07844_, _07781_);
  not _16146_ (_07846_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _16147_ (_07847_, _07613_, _07846_);
  or _16148_ (_07848_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _16149_ (_07849_, _07848_, _07847_);
  and _16150_ (_07850_, _07849_, _07821_);
  not _16151_ (_07851_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _16152_ (_07852_, _07613_, _07851_);
  or _16153_ (_07853_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _16154_ (_07854_, _07853_, _07852_);
  and _16155_ (_07855_, _07854_, _07820_);
  or _16156_ (_07856_, _07855_, _07850_);
  and _16157_ (_07857_, _07856_, _07807_);
  not _16158_ (_07858_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _16159_ (_07859_, _07613_, _07858_);
  or _16160_ (_07860_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _16161_ (_07861_, _07860_, _07859_);
  and _16162_ (_07862_, _07861_, _07821_);
  not _16163_ (_07864_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _16164_ (_07865_, _07613_, _07864_);
  or _16165_ (_07867_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _16166_ (_07868_, _07867_, _07865_);
  and _16167_ (_07870_, _07868_, _07820_);
  or _16168_ (_07871_, _07870_, _07862_);
  and _16169_ (_07872_, _07871_, _07811_);
  or _16170_ (_07874_, _07872_, _07857_);
  or _16171_ (_07875_, _07874_, _07845_);
  nor _16172_ (_07877_, _07875_, _07833_);
  nor _16173_ (_07878_, _07877_, _07819_);
  and _16174_ (_07880_, _07819_, word_in[15]);
  or _16175_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _07880_, _07878_);
  nor _16176_ (_07882_, _07666_, _07650_);
  not _16177_ (_07883_, _07882_);
  nor _16178_ (_07884_, _07883_, _07629_);
  nor _16179_ (_07886_, _07650_, _07626_);
  and _16180_ (_07887_, _07650_, _07626_);
  nor _16181_ (_07888_, _07887_, _07886_);
  and _16182_ (_07889_, _07888_, _07883_);
  and _16183_ (_07890_, _07889_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _16184_ (_07891_, _07888_, _07882_);
  and _16185_ (_07892_, _07891_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16186_ (_07893_, _07892_, _07890_);
  nor _16187_ (_07894_, _07893_, _07884_);
  nor _16188_ (_07895_, _07894_, _07806_);
  and _16189_ (_07896_, _07891_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _16190_ (_07897_, _07896_);
  nor _16191_ (_07898_, _07883_, _07656_);
  and _16192_ (_07899_, _07889_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16193_ (_07900_, _07899_, _07898_);
  and _16194_ (_07901_, _07900_, _07897_);
  nor _16195_ (_07902_, _07901_, _07789_);
  nor _16196_ (_07903_, _07902_, _07895_);
  nor _16197_ (_07904_, _07883_, _07694_);
  and _16198_ (_07905_, _07889_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16199_ (_07906_, _07891_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16200_ (_07907_, _07906_, _07905_);
  nor _16201_ (_07908_, _07907_, _07904_);
  nor _16202_ (_07909_, _07908_, _07763_);
  nor _16203_ (_07910_, _07883_, _07699_);
  and _16204_ (_07911_, _07889_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16205_ (_07912_, _07891_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _16206_ (_07913_, _07912_, _07911_);
  nor _16207_ (_07914_, _07913_, _07910_);
  nor _16208_ (_07915_, _07914_, _07799_);
  nor _16209_ (_07916_, _07915_, _07909_);
  and _16210_ (_07917_, _07916_, _07903_);
  and _16211_ (_07918_, _07917_, word_in[23]);
  and _16212_ (_07919_, _07744_, _07643_);
  and _16213_ (_07920_, _07733_, _07666_);
  or _16214_ (_07921_, _07920_, _07919_);
  and _16215_ (_07922_, _07738_, _07640_);
  and _16216_ (_07923_, _07750_, _07650_);
  or _16217_ (_07924_, _07923_, _07922_);
  or _16218_ (_07925_, _07924_, _07921_);
  or _16219_ (_07926_, _07925_, _07888_);
  not _16220_ (_07927_, _07888_);
  and _16221_ (_07928_, _07720_, _07643_);
  and _16222_ (_07929_, _07714_, _07666_);
  or _16223_ (_07930_, _07929_, _07928_);
  and _16224_ (_07931_, _07709_, _07640_);
  and _16225_ (_07932_, _07725_, _07650_);
  or _16226_ (_07933_, _07932_, _07931_);
  or _16227_ (_07934_, _07933_, _07930_);
  or _16228_ (_07935_, _07934_, _07927_);
  nand _16229_ (_07936_, _07935_, _07926_);
  nor _16230_ (_07937_, _07936_, _07917_);
  or _16231_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _07937_, _07918_);
  nor _16232_ (_07938_, _07763_, _07639_);
  not _16233_ (_07939_, _07938_);
  nand _16234_ (_07940_, _07763_, _07639_);
  and _16235_ (_07941_, _07940_, _07939_);
  not _16236_ (_07942_, _07941_);
  nor _16237_ (_07943_, _07699_, _07942_);
  nor _16238_ (_07944_, _07940_, _07626_);
  and _16239_ (_07945_, _07940_, _07626_);
  nor _16240_ (_07946_, _07945_, _07944_);
  and _16241_ (_07947_, _07946_, _07942_);
  and _16242_ (_07948_, _07947_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16243_ (_07949_, _07946_, _07941_);
  and _16244_ (_07950_, _07949_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _16245_ (_07951_, _07950_, _07948_);
  nor _16246_ (_07952_, _07951_, _07943_);
  nor _16247_ (_07954_, _07952_, _07789_);
  and _16248_ (_07955_, _07938_, _07646_);
  nor _16249_ (_07956_, _07942_, _07656_);
  and _16250_ (_07958_, _07949_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _16251_ (_07959_, _07958_, _07956_);
  and _16252_ (_07960_, _07959_, _07761_);
  nor _16253_ (_07962_, _07960_, _07955_);
  not _16254_ (_07963_, _07962_);
  nor _16255_ (_07964_, _07963_, _07954_);
  nor _16256_ (_07966_, _07694_, _07942_);
  and _16257_ (_07967_, _07949_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16258_ (_07968_, _07947_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16259_ (_07970_, _07968_, _07967_);
  nor _16260_ (_07972_, _07970_, _07966_);
  nor _16261_ (_07973_, _07972_, _07806_);
  nor _16262_ (_07975_, _07942_, _07629_);
  and _16263_ (_07977_, _07949_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16264_ (_07978_, _07947_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16265_ (_07979_, _07978_, _07977_);
  nor _16266_ (_07980_, _07979_, _07975_);
  nor _16267_ (_07982_, _07980_, _07799_);
  nor _16268_ (_07983_, _07982_, _07973_);
  and _16269_ (_07984_, _07983_, _07964_);
  and _16270_ (_07985_, _07842_, _07821_);
  and _16271_ (_07986_, _07837_, _07820_);
  or _16272_ (_07987_, _07986_, _07985_);
  and _16273_ (_07988_, _07987_, _07947_);
  and _16274_ (_07989_, _07830_, _07821_);
  and _16275_ (_07990_, _07825_, _07820_);
  or _16276_ (_07991_, _07990_, _07989_);
  and _16277_ (_07992_, _07991_, _07949_);
  and _16278_ (_07993_, _07941_, _07676_);
  and _16279_ (_07994_, _07854_, _07821_);
  and _16280_ (_07995_, _07849_, _07820_);
  or _16281_ (_07996_, _07995_, _07994_);
  and _16282_ (_07997_, _07996_, _07993_);
  and _16283_ (_07998_, _07868_, _07821_);
  and _16284_ (_07999_, _07861_, _07820_);
  or _16285_ (_08000_, _07999_, _07998_);
  and _16286_ (_08001_, _07945_, _07939_);
  and _16287_ (_08002_, _08001_, _08000_);
  or _16288_ (_08003_, _08002_, _07997_);
  or _16289_ (_08004_, _08003_, _07992_);
  nor _16290_ (_08005_, _08004_, _07988_);
  nor _16291_ (_08006_, _08005_, _07984_);
  and _16292_ (_08007_, _07984_, word_in[31]);
  or _16293_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08007_, _08006_);
  and _16294_ (_08008_, _07639_, _07626_);
  or _16295_ (_08009_, _08008_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _16296_ (_06029_, _08009_, _05141_);
  and _16297_ (_08010_, _07984_, _05141_);
  and _16298_ (_08011_, _08010_, word_in[31]);
  and _16299_ (_08012_, _08008_, _07761_);
  and _16300_ (_08013_, _08010_, _08012_);
  and _16301_ (_08014_, _08013_, _08011_);
  not _16302_ (_08015_, _08013_);
  and _16303_ (_08016_, _07917_, _05141_);
  and _16304_ (_08017_, _08016_, _07882_);
  and _16305_ (_08018_, _08017_, _07888_);
  and _16306_ (_08019_, _08018_, _07788_);
  not _16307_ (_08020_, _08019_);
  and _16308_ (_08021_, _07819_, _05141_);
  and _16309_ (_08022_, _08021_, _07798_);
  and _16310_ (_08023_, _08022_, _07811_);
  and _16311_ (_08024_, _07673_, _05141_);
  and _16312_ (_08025_, _08024_, _07633_);
  nor _16313_ (_08026_, _07705_, rst);
  and _16314_ (_08027_, _08026_, _08008_);
  and _16315_ (_08028_, _08027_, _08025_);
  and _16316_ (_08029_, _08026_, word_in[7]);
  and _16317_ (_08030_, _08029_, _08028_);
  nor _16318_ (_08031_, _08028_, _07706_);
  nor _16319_ (_08032_, _08031_, _08030_);
  nor _16320_ (_08033_, _08032_, _08023_);
  and _16321_ (_08034_, _08023_, word_in[15]);
  or _16322_ (_08035_, _08034_, _08033_);
  and _16323_ (_08036_, _08035_, _08020_);
  and _16324_ (_08037_, _08016_, word_in[23]);
  and _16325_ (_08038_, _08037_, _08019_);
  or _16326_ (_08039_, _08038_, _08036_);
  and _16327_ (_08040_, _08039_, _08015_);
  or _16328_ (_06058_, _08040_, _08014_);
  or _16329_ (_08041_, _07947_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _16330_ (_06079_, _08041_, _05141_);
  and _16331_ (_08043_, _07798_, _07947_);
  and _16332_ (_08044_, _07766_, _07626_);
  and _16333_ (_08046_, _07666_, _07676_);
  or _16334_ (_08047_, _08046_, _08044_);
  or _16335_ (_08049_, _08047_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16336_ (_08050_, _08049_, _08043_);
  and _16337_ (_06108_, _08050_, _05141_);
  and _16338_ (_08052_, _07993_, _07798_);
  or _16339_ (_08054_, _08052_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16340_ (_08055_, _08054_, _08047_);
  and _16341_ (_06149_, _08055_, _05141_);
  or _16342_ (_08057_, _07639_, _07626_);
  nand _16343_ (_08059_, _08057_, _07645_);
  and _16344_ (_06196_, _08059_, _05141_);
  or _16345_ (_08061_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand _16346_ (_08062_, _07619_, _06347_);
  and _16347_ (_08063_, _08062_, _05141_);
  and _16348_ (_06232_, _08063_, _08061_);
  and _16349_ (_08064_, _07993_, _07765_);
  and _16350_ (_08065_, _07777_, _07761_);
  or _16351_ (_08066_, _08065_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _16352_ (_08067_, _08066_, _08057_);
  nor _16353_ (_08068_, _08067_, _08064_);
  nor _16354_ (_08069_, _08068_, _07781_);
  and _16355_ (_08070_, _07821_, _07993_);
  and _16356_ (_08071_, _07938_, _07676_);
  or _16357_ (_08072_, _08071_, _08044_);
  and _16358_ (_08073_, _08072_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _16359_ (_08074_, _08073_, _08070_);
  or _16360_ (_08075_, _08074_, _08069_);
  and _16361_ (_06252_, _08075_, _05141_);
  not _16362_ (_08076_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _16363_ (_08077_, _05622_, _08076_);
  not _16364_ (_08078_, _05622_);
  nor _16365_ (_08079_, _06062_, _08078_);
  or _16366_ (_08080_, _08079_, _08077_);
  and _16367_ (_06258_, _08080_, _05141_);
  not _16368_ (_08081_, _08057_);
  nor _16369_ (_08082_, _08081_, _08044_);
  not _16370_ (_08083_, _07886_);
  or _16371_ (_08084_, _08065_, _08064_);
  or _16372_ (_08085_, _08084_, _08083_);
  and _16373_ (_08086_, _08085_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _16374_ (_08087_, _07788_, _07777_);
  and _16375_ (_08088_, _08046_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _16376_ (_08089_, _08052_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16377_ (_08090_, _08089_, _08088_);
  or _16378_ (_08091_, _08090_, _08087_);
  or _16379_ (_08092_, _08091_, _08086_);
  or _16380_ (_08093_, _07774_, _07944_);
  and _16381_ (_08094_, _08093_, _08092_);
  and _16382_ (_08095_, _07993_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16383_ (_08096_, _08095_, _08065_);
  or _16384_ (_08097_, _08096_, _08094_);
  and _16385_ (_08098_, _08097_, _08082_);
  and _16386_ (_08099_, _08092_, _08044_);
  and _16387_ (_08100_, _08071_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _16388_ (_08101_, _07788_, _07993_);
  and _16389_ (_08102_, _08101_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16390_ (_08103_, _08102_, _08052_);
  or _16391_ (_08104_, _08103_, _08100_);
  or _16392_ (_08105_, _08104_, _08064_);
  or _16393_ (_08106_, _08105_, _08099_);
  or _16394_ (_08107_, _08106_, _08098_);
  and _16395_ (_06294_, _08107_, _05141_);
  nand _16396_ (_08108_, _07639_, _07613_);
  nand _16397_ (_08109_, _07886_, _08108_);
  and _16398_ (_08110_, _07798_, _07777_);
  or _16399_ (_08111_, _08110_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _16400_ (_08112_, _08111_, _08109_);
  and _16401_ (_08113_, _08112_, _08083_);
  and _16402_ (_08114_, _08084_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _16403_ (_08115_, _08114_, _08087_);
  or _16404_ (_08116_, _08115_, _08113_);
  and _16405_ (_08117_, _08116_, _08093_);
  and _16406_ (_08118_, _08111_, _08044_);
  and _16407_ (_08119_, _08052_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _16408_ (_08121_, _08046_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _16409_ (_08122_, _08121_, _08064_);
  or _16410_ (_08124_, _08122_, _08119_);
  or _16411_ (_08125_, _08124_, _08065_);
  or _16412_ (_08126_, _08125_, _08118_);
  or _16413_ (_08127_, _08126_, _08117_);
  and _16414_ (_06359_, _08127_, _05141_);
  and _16415_ (_08128_, _05622_, _05522_);
  not _16416_ (_08129_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor _16417_ (_08130_, _05622_, _08129_);
  or _16418_ (_08131_, _08130_, _08128_);
  and _16419_ (_06405_, _08131_, _05141_);
  not _16420_ (_08132_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _16421_ (_08133_, _05622_, _08132_);
  nor _16422_ (_08134_, _08078_, _05560_);
  or _16423_ (_08135_, _08134_, _08133_);
  and _16424_ (_06424_, _08135_, _05141_);
  and _16425_ (_08136_, _07821_, _07777_);
  and _16426_ (_08137_, _07941_, _07653_);
  and _16427_ (_08138_, _07938_, _07653_);
  or _16428_ (_08139_, _08138_, _08065_);
  or _16429_ (_08140_, _08139_, _08137_);
  or _16430_ (_08142_, _07766_, _07626_);
  and _16431_ (_08143_, _07653_, _07776_);
  or _16432_ (_08144_, _08110_, _07626_);
  and _16433_ (_08145_, _08144_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _16434_ (_08146_, _07633_, _07652_);
  and _16435_ (_08147_, _08146_, _07777_);
  or _16436_ (_08148_, _08147_, _07779_);
  or _16437_ (_08149_, _08148_, _08145_);
  or _16438_ (_08150_, _08149_, _08143_);
  and _16439_ (_08151_, _08150_, _08142_);
  or _16440_ (_08152_, _08151_, _08140_);
  or _16441_ (_08153_, _08152_, _08136_);
  and _16442_ (_06435_, _08153_, _05141_);
  and _16443_ (_08154_, _06179_, _05622_);
  not _16444_ (_08155_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor _16445_ (_08156_, _05622_, _08155_);
  or _16446_ (_08157_, _08156_, _08154_);
  and _16447_ (_06443_, _08157_, _05141_);
  not _16448_ (_08158_, _06836_);
  nor _16449_ (_08159_, _06207_, _05708_);
  or _16450_ (_08160_, _08159_, _06208_);
  or _16451_ (_08161_, _06838_, _06836_);
  nor _16452_ (_08162_, _08161_, _06841_);
  and _16453_ (_08163_, _08162_, _06881_);
  nand _16454_ (_08164_, _08163_, _08160_);
  and _16455_ (_08165_, _06884_, _06669_);
  and _16456_ (_08166_, _05256_, _05172_);
  and _16457_ (_08167_, _08166_, _06879_);
  and _16458_ (_08168_, _08167_, _05241_);
  and _16459_ (_08169_, _08168_, _05647_);
  not _16460_ (_08170_, _08169_);
  and _16461_ (_08171_, _08170_, _08162_);
  and _16462_ (_08172_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _16463_ (_08173_, _08172_, _08165_);
  nand _16464_ (_08174_, _08173_, _08164_);
  nand _16465_ (_08175_, _08174_, _08158_);
  nand _16466_ (_08176_, _07288_, _06836_);
  nand _16467_ (_08177_, _08176_, _08175_);
  and _16468_ (_06503_, _08177_, _05141_);
  and _16469_ (_08178_, _05922_, _05288_);
  nor _16470_ (_08179_, _05288_, _05441_);
  or _16471_ (_08180_, _08179_, _08178_);
  nand _16472_ (_08181_, _08180_, _08163_);
  and _16473_ (_08182_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _16474_ (_08183_, _07434_, _06842_);
  nor _16475_ (_08184_, _08183_, _08182_);
  and _16476_ (_08185_, _08184_, _08158_);
  nand _16477_ (_08186_, _08185_, _08181_);
  or _16478_ (_08187_, _07406_, _08158_);
  and _16479_ (_08188_, _08187_, _08186_);
  and _16480_ (_06507_, _08188_, _05141_);
  and _16481_ (_08189_, _07938_, _07626_);
  or _16482_ (_08190_, _08189_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16483_ (_08191_, _08190_, _07626_);
  not _16484_ (_08192_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _16485_ (_08193_, _08057_, _08192_);
  and _16486_ (_08194_, _08065_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _16487_ (_08195_, _08087_, _07779_);
  or _16488_ (_08196_, _08195_, _08194_);
  or _16489_ (_08197_, _08196_, _08193_);
  or _16490_ (_08198_, _08197_, _08191_);
  or _16491_ (_08199_, _08198_, _08110_);
  and _16492_ (_06513_, _08199_, _05141_);
  and _16493_ (_08200_, _07886_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16494_ (_08201_, _07939_, _07626_);
  and _16495_ (_08202_, _08201_, _07773_);
  and _16496_ (_08203_, _08001_, _07788_);
  nor _16497_ (_08204_, _07886_, _07661_);
  or _16498_ (_08205_, _08204_, _08203_);
  and _16499_ (_08206_, _08205_, _08202_);
  and _16500_ (_08207_, _07650_, _07676_);
  and _16501_ (_08208_, _08207_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _16502_ (_08209_, _08208_, _08189_);
  or _16503_ (_08211_, _08209_, _08206_);
  and _16504_ (_08212_, _08211_, _07774_);
  and _16505_ (_08213_, _08205_, _08044_);
  or _16506_ (_08214_, _08213_, _08207_);
  or _16507_ (_08215_, _08214_, _08212_);
  or _16508_ (_08216_, _08215_, _08200_);
  and _16509_ (_06609_, _08216_, _05141_);
  and _16510_ (_08217_, _07798_, _07945_);
  not _16511_ (_08218_, _07768_);
  and _16512_ (_08220_, _08218_, _07674_);
  or _16513_ (_08221_, _08220_, _08217_);
  and _16514_ (_08222_, _08046_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16515_ (_08223_, _07882_, _07676_);
  and _16516_ (_08225_, _08223_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16517_ (_08226_, _08110_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _16518_ (_08227_, _08226_, _07779_);
  or _16519_ (_08228_, _08227_, _08225_);
  or _16520_ (_08230_, _08228_, _08222_);
  or _16521_ (_08231_, _08230_, _08203_);
  or _16522_ (_08232_, _08231_, _08189_);
  or _16523_ (_08233_, _08232_, _08221_);
  and _16524_ (_06704_, _08233_, _05141_);
  and _16525_ (_08235_, _06004_, _05622_);
  not _16526_ (_08237_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _16527_ (_08238_, _05622_, _08237_);
  or _16528_ (_08239_, _08238_, _08235_);
  and _16529_ (_06712_, _08239_, _05141_);
  and _16530_ (_08241_, _05648_, _05281_);
  and _16531_ (_08242_, _06736_, _05288_);
  and _16532_ (_08243_, _08242_, _08241_);
  and _16533_ (_08245_, _06691_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _16534_ (_08246_, _08245_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or _16535_ (_08247_, _08246_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _16536_ (_08248_, _08246_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _16537_ (_08249_, _08248_, rst);
  nand _16538_ (_08250_, _08249_, _08247_);
  nor _16539_ (_06717_, _08250_, _08243_);
  and _16540_ (_08251_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and _16541_ (_08252_, _06275_, _05561_);
  or _16542_ (_08253_, _08252_, _08251_);
  and _16543_ (_06783_, _08253_, _05141_);
  and _16544_ (_08254_, _07945_, _07765_);
  and _16545_ (_08255_, _08008_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _16546_ (_08256_, _08255_, _08254_);
  not _16547_ (_08257_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16548_ (_08258_, _07626_, _08257_);
  or _16549_ (_08259_, _08189_, _08217_);
  or _16550_ (_08260_, _08259_, _08258_);
  or _16551_ (_08261_, _08260_, _08203_);
  or _16552_ (_08262_, _08261_, _08256_);
  and _16553_ (_06794_, _08262_, _05141_);
  and _16554_ (_08263_, _08248_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _16555_ (_08264_, _08263_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _16556_ (_08265_, _08263_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _16557_ (_08266_, _08265_, _08264_);
  nand _16558_ (_08267_, _08266_, _05141_);
  nor _16559_ (_06817_, _08267_, _08243_);
  and _16560_ (_08268_, _08008_, _07763_);
  and _16561_ (_08269_, _08268_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _16562_ (_08270_, _07678_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _16563_ (_08271_, _08189_, _08046_);
  or _16564_ (_08272_, _08271_, _07777_);
  and _16565_ (_08273_, _08272_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _16566_ (_08274_, _08273_, _08001_);
  or _16567_ (_08275_, _08274_, _08270_);
  or _16568_ (_08276_, _08275_, _08269_);
  and _16569_ (_06887_, _08276_, _05141_);
  or _16570_ (_08277_, _08248_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _16571_ (_08278_, _08263_, rst);
  nand _16572_ (_08279_, _08278_, _08277_);
  nor _16573_ (_06903_, _08279_, _08243_);
  and _16574_ (_08280_, _06012_, _06202_);
  and _16575_ (_08281_, _05922_, _06032_);
  or _16576_ (_08282_, _05650_, _06007_);
  not _16577_ (_08283_, _08282_);
  and _16578_ (_08284_, _08283_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _16579_ (_08285_, _08284_, _08281_);
  and _16580_ (_08286_, _08285_, _08280_);
  nand _16581_ (_08287_, _08280_, _05186_);
  and _16582_ (_08288_, _08287_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _16583_ (_08289_, _08241_, _05926_);
  or _16584_ (_08290_, _08289_, _08288_);
  or _16585_ (_08291_, _08290_, _08286_);
  nand _16586_ (_08292_, _08289_, _06062_);
  and _16587_ (_08293_, _08292_, _05141_);
  and _16588_ (_06957_, _08293_, _08291_);
  not _16589_ (_08294_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _16590_ (_08295_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _16591_ (_08296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _08295_);
  nand _16592_ (_08297_, _08296_, _08294_);
  or _16593_ (_08298_, _08296_, rxd_i);
  and _16594_ (_08299_, _08298_, _08297_);
  nor _16595_ (_08300_, _06683_, _06690_);
  and _16596_ (_08301_, _08300_, _06686_);
  and _16597_ (_08302_, _08301_, _08299_);
  nor _16598_ (_08303_, _08301_, _08294_);
  or _16599_ (_08304_, _08303_, rst);
  or _16600_ (_06960_, _08304_, _08302_);
  and _16601_ (_08305_, _06621_, _06008_);
  not _16602_ (_08306_, _08305_);
  or _16603_ (_08307_, _08306_, _06004_);
  or _16604_ (_08308_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _16605_ (_08309_, _08308_, _05141_);
  and _16606_ (_06962_, _08309_, _08307_);
  nand _16607_ (_08311_, _08305_, _05604_);
  or _16608_ (_08313_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _16609_ (_08315_, _08313_, _05141_);
  and _16610_ (_06966_, _08315_, _08311_);
  nor _16611_ (_08316_, _07634_, _07626_);
  or _16612_ (_08318_, _08316_, _07887_);
  and _16613_ (_08319_, _08318_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _16614_ (_08320_, _07643_, _07626_);
  or _16615_ (_08322_, _08012_, _08320_);
  nor _16616_ (_08323_, _08008_, _07614_);
  or _16617_ (_08324_, _08323_, _08268_);
  and _16618_ (_08326_, _08324_, _07634_);
  or _16619_ (_08327_, _08326_, _08322_);
  or _16620_ (_08328_, _08327_, _08319_);
  and _16621_ (_06971_, _08328_, _05141_);
  not _16622_ (_08330_, _06821_);
  and _16623_ (_08332_, _06765_, _06536_);
  and _16624_ (_08333_, _06574_, _06449_);
  and _16625_ (_08334_, _08333_, _06536_);
  or _16626_ (_08336_, _08334_, _06784_);
  nor _16627_ (_08337_, _08336_, _08332_);
  or _16628_ (_08338_, _08337_, _08330_);
  nor _16629_ (_08339_, _06538_, _06474_);
  and _16630_ (_08340_, _08339_, _06550_);
  and _16631_ (_08341_, _08340_, _07088_);
  not _16632_ (_08342_, _08341_);
  and _16633_ (_08343_, _08342_, _06796_);
  nand _16634_ (_08344_, _08343_, _08338_);
  and _16635_ (_06984_, _08344_, _05141_);
  not _16636_ (_08345_, _06738_);
  nor _16637_ (_08346_, _08345_, _06244_);
  and _16638_ (_08347_, _06736_, _06032_);
  and _16639_ (_08348_, _08347_, _06734_);
  and _16640_ (_08349_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _16641_ (_08350_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _16642_ (_08351_, _08350_, _08349_);
  nor _16643_ (_08352_, _08351_, _06738_);
  or _16644_ (_08353_, _08352_, _08348_);
  or _16645_ (_08354_, _08353_, _08346_);
  not _16646_ (_08355_, _08348_);
  or _16647_ (_08356_, _08355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _16648_ (_08357_, _08356_, _05141_);
  and _16649_ (_06991_, _08357_, _08354_);
  and _16650_ (_08358_, _08280_, _06207_);
  nand _16651_ (_08359_, _08358_, _05963_);
  not _16652_ (_08360_, _08289_);
  or _16653_ (_08361_, _08358_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _16654_ (_08362_, _08361_, _08360_);
  and _16655_ (_08363_, _08362_, _08359_);
  nor _16656_ (_08364_, _08360_, _06244_);
  or _16657_ (_08365_, _08364_, _08363_);
  and _16658_ (_07024_, _08365_, _05141_);
  not _16659_ (_08366_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _16660_ (_08367_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _08366_);
  or _16661_ (_08368_, _08367_, _06683_);
  nor _16662_ (_08369_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _16663_ (_08370_, _08369_, _08368_);
  or _16664_ (_08371_, _08370_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _16665_ (_08372_, _08371_, _08280_);
  and _16666_ (_08373_, _05922_, _05210_);
  not _16667_ (_08374_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _16668_ (_08375_, _05210_, _08374_);
  nand _16669_ (_08376_, _08375_, _08280_);
  or _16670_ (_08377_, _08376_, _08373_);
  and _16671_ (_08378_, _08377_, _08372_);
  or _16672_ (_08379_, _08378_, _08289_);
  nand _16673_ (_08380_, _08289_, _05604_);
  and _16674_ (_08381_, _08380_, _05141_);
  and _16675_ (_07027_, _08381_, _08379_);
  and _16676_ (_08382_, _08243_, _06683_);
  and _16677_ (_08383_, _08382_, _05561_);
  and _16678_ (_08384_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _16679_ (_08385_, _08384_, _06683_);
  nor _16680_ (_08386_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _16681_ (_08387_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _16682_ (_08388_, _08387_, _08386_);
  and _16683_ (_08389_, _08388_, _08246_);
  nor _16684_ (_08390_, _08389_, _08385_);
  not _16685_ (_08391_, _08390_);
  and _16686_ (_08392_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _16687_ (_08393_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _16688_ (_08394_, _08393_, _08392_);
  nor _16689_ (_08395_, _08394_, _08243_);
  and _16690_ (_08396_, _08243_, _06691_);
  and _16691_ (_08397_, _08396_, _06179_);
  or _16692_ (_08398_, _08397_, _08395_);
  or _16693_ (_08399_, _08398_, _08383_);
  and _16694_ (_07038_, _08399_, _05141_);
  and _16695_ (_08401_, _07319_, _06836_);
  and _16696_ (_08402_, _06881_, _06032_);
  nand _16697_ (_08404_, _08402_, _05963_);
  not _16698_ (_08405_, _08162_);
  nor _16699_ (_08406_, _08402_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _16700_ (_08408_, _08406_, _08405_);
  and _16701_ (_08409_, _08408_, _08404_);
  nor _16702_ (_08411_, _07350_, _06842_);
  or _16703_ (_08412_, _08411_, _08409_);
  and _16704_ (_08414_, _08412_, _08158_);
  or _16705_ (_08415_, _08414_, _08401_);
  and _16706_ (_07061_, _08415_, _05141_);
  nor _16707_ (_08417_, _06738_, _06730_);
  or _16708_ (_08418_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  not _16709_ (_08420_, _08417_);
  or _16710_ (_08422_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _16711_ (_08423_, _08422_, _08418_);
  and _16712_ (_08424_, _08423_, _08355_);
  nor _16713_ (_08425_, _08355_, _06062_);
  or _16714_ (_08426_, _08425_, _08424_);
  and _16715_ (_07075_, _08426_, _05141_);
  or _16716_ (_08427_, _07811_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _16717_ (_07082_, _08427_, _05141_);
  nand _16718_ (_08428_, _06743_, _06244_);
  or _16719_ (_08429_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _16720_ (_08430_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _16721_ (_08431_, _08430_, _08429_);
  or _16722_ (_08432_, _08431_, _06743_);
  and _16723_ (_08433_, _08432_, _05141_);
  and _16724_ (_07095_, _08433_, _08428_);
  and _16725_ (_08434_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not _16726_ (_08435_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _16727_ (_08436_, \oc8051_top_1.oc8051_sfr1.pres_ow , _08435_);
  nor _16728_ (_08437_, _08436_, _08434_);
  not _16729_ (_08438_, _08437_);
  and _16730_ (_08439_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _16731_ (_08440_, _08439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  not _16732_ (_08441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor _16733_ (_08442_, _06727_, _08441_);
  and _16734_ (_08443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _16735_ (_08444_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _16736_ (_08445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _16737_ (_08446_, _08445_, _08444_);
  and _16738_ (_08447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _16739_ (_08448_, _08447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _16740_ (_08449_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _16741_ (_08450_, _08449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _16742_ (_08451_, _08450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _16743_ (_08452_, _08451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _16744_ (_08453_, _08452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _16745_ (_08454_, _08453_, _08446_);
  and _16746_ (_08455_, _08454_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _16747_ (_08456_, _08455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _16748_ (_08457_, _08456_, _08443_);
  nand _16749_ (_08458_, _08457_, _08442_);
  nand _16750_ (_08459_, _08458_, _08440_);
  not _16751_ (_08460_, _06726_);
  not _16752_ (_08461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _16753_ (_08462_, _06725_, _08461_);
  nor _16754_ (_08463_, _08462_, _08460_);
  not _16755_ (_08464_, _08463_);
  or _16756_ (_08465_, _08439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _16757_ (_08466_, _08465_, _08464_);
  and _16758_ (_08467_, _08466_, _08459_);
  and _16759_ (_08468_, _08463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _16760_ (_08469_, _05209_, _06007_);
  and _16761_ (_08470_, _06736_, _08469_);
  and _16762_ (_08471_, _08470_, _06734_);
  or _16763_ (_08472_, _08471_, _08468_);
  or _16764_ (_08474_, _08472_, _08467_);
  nand _16765_ (_08475_, _08471_, _05604_);
  and _16766_ (_08476_, _05964_, _05925_);
  and _16767_ (_08478_, _08476_, _06734_);
  not _16768_ (_08479_, _08478_);
  and _16769_ (_08480_, _08479_, _08475_);
  and _16770_ (_08481_, _08480_, _08474_);
  and _16771_ (_08482_, _08478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _16772_ (_08483_, _08482_, _08481_);
  and _16773_ (_07098_, _08483_, _05141_);
  not _16774_ (_08484_, _05277_);
  nor _16775_ (_08485_, _06062_, _08484_);
  not _16776_ (_08487_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _16777_ (_08488_, _05277_, _08487_);
  or _16778_ (_08489_, _08488_, _05572_);
  or _16779_ (_08491_, _08489_, _08485_);
  or _16780_ (_08492_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _16781_ (_08494_, _08492_, _05141_);
  and _16782_ (_07122_, _08494_, _08491_);
  nand _16783_ (_08496_, _07466_, _06836_);
  nor _16784_ (_08497_, _05210_, _05420_);
  or _16785_ (_08499_, _08497_, _08373_);
  nand _16786_ (_08500_, _08499_, _08163_);
  nor _16787_ (_08501_, _06881_, _05420_);
  nor _16788_ (_08503_, _08501_, _06884_);
  and _16789_ (_08504_, _08503_, _08500_);
  nor _16790_ (_08505_, _07496_, _06836_);
  nor _16791_ (_08507_, _08505_, _08162_);
  or _16792_ (_08508_, _08507_, _08504_);
  nand _16793_ (_08509_, _08508_, _08496_);
  and _16794_ (_07160_, _08509_, _05141_);
  and _16795_ (_08511_, _08396_, _06703_);
  and _16796_ (_08512_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _16797_ (_08513_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _16798_ (_08514_, _08513_, _08512_);
  nor _16799_ (_08515_, _08514_, _08243_);
  and _16800_ (_08516_, _08382_, _06179_);
  or _16801_ (_08518_, _08516_, _08515_);
  or _16802_ (_08519_, _08518_, _08511_);
  and _16803_ (_07165_, _08519_, _05141_);
  and _16804_ (_08520_, _05299_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _16805_ (_08521_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _16806_ (_08522_, _08521_, _05303_);
  and _16807_ (_08523_, _06179_, _05523_);
  or _16808_ (_08524_, _08523_, _08522_);
  or _16809_ (_08525_, _08524_, _08520_);
  and _16810_ (_07247_, _08525_, _05141_);
  and _16811_ (_08526_, _08016_, _08043_);
  not _16812_ (_08527_, _08526_);
  and _16813_ (_08528_, _08021_, _08044_);
  not _16814_ (_08529_, _08528_);
  and _16815_ (_08530_, _08026_, _07633_);
  nor _16816_ (_08531_, _08530_, _08024_);
  and _16817_ (_08532_, _08026_, _08081_);
  and _16818_ (_08533_, _08532_, _08531_);
  and _16819_ (_08534_, _08533_, word_in[0]);
  not _16820_ (_08535_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _16821_ (_08536_, _08533_, _08535_);
  or _16822_ (_08537_, _08536_, _08534_);
  and _16823_ (_08538_, _08537_, _08529_);
  and _16824_ (_08539_, _08528_, word_in[8]);
  or _16825_ (_08540_, _08539_, _08538_);
  and _16826_ (_08541_, _08540_, _08527_);
  and _16827_ (_08542_, _07788_, _08008_);
  and _16828_ (_08543_, _08010_, _08542_);
  and _16829_ (_08544_, _08016_, word_in[16]);
  and _16830_ (_08545_, _08544_, _08043_);
  or _16831_ (_08546_, _08545_, _08543_);
  or _16832_ (_08547_, _08546_, _08541_);
  not _16833_ (_08548_, _08543_);
  or _16834_ (_08549_, _08548_, word_in[24]);
  and _16835_ (_07443_, _08549_, _08547_);
  or _16836_ (_08550_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not _16837_ (_08551_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _16838_ (_08552_, pc_log_change, _08551_);
  and _16839_ (_08553_, _08552_, _05141_);
  and _16840_ (_07446_, _08553_, _08550_);
  not _16841_ (_08554_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _16842_ (_08555_, _08533_, _08554_);
  and _16843_ (_08556_, _08026_, word_in[1]);
  and _16844_ (_08557_, _08556_, _08533_);
  or _16845_ (_08558_, _08557_, _08555_);
  or _16846_ (_08559_, _08558_, _08528_);
  or _16847_ (_08560_, _08529_, word_in[9]);
  and _16848_ (_08561_, _08560_, _08559_);
  or _16849_ (_08562_, _08561_, _08526_);
  nor _16850_ (_08563_, _08527_, word_in[17]);
  nor _16851_ (_08564_, _08563_, _08543_);
  and _16852_ (_08565_, _08564_, _08562_);
  and _16853_ (_08566_, _08010_, word_in[25]);
  and _16854_ (_08567_, _08566_, _08543_);
  or _16855_ (_07449_, _08567_, _08565_);
  and _16856_ (_08568_, _08010_, word_in[26]);
  and _16857_ (_08569_, _08568_, _08543_);
  not _16858_ (_08570_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _16859_ (_08571_, _08533_, _08570_);
  and _16860_ (_08572_, _08026_, word_in[2]);
  and _16861_ (_08573_, _08572_, _08533_);
  or _16862_ (_08574_, _08573_, _08571_);
  or _16863_ (_08575_, _08574_, _08528_);
  or _16864_ (_08576_, _08529_, word_in[10]);
  and _16865_ (_08577_, _08576_, _08575_);
  or _16866_ (_08578_, _08577_, _08526_);
  nor _16867_ (_08579_, _08527_, word_in[18]);
  nor _16868_ (_08580_, _08579_, _08543_);
  and _16869_ (_08581_, _08580_, _08578_);
  or _16870_ (_07454_, _08581_, _08569_);
  nor _16871_ (_07457_, _05625_, rst);
  and _16872_ (_08582_, _08010_, word_in[27]);
  and _16873_ (_08583_, _08582_, _08543_);
  not _16874_ (_08584_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _16875_ (_08585_, _08533_, _08584_);
  and _16876_ (_08586_, _08026_, word_in[3]);
  and _16877_ (_08587_, _08586_, _08533_);
  or _16878_ (_08588_, _08587_, _08585_);
  and _16879_ (_08589_, _08588_, _08529_);
  and _16880_ (_08590_, _08528_, word_in[11]);
  or _16881_ (_08591_, _08590_, _08589_);
  or _16882_ (_08592_, _08591_, _08526_);
  nor _16883_ (_08593_, _08527_, word_in[19]);
  nor _16884_ (_08594_, _08593_, _08543_);
  and _16885_ (_08595_, _08594_, _08592_);
  or _16886_ (_07460_, _08595_, _08583_);
  not _16887_ (_08596_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _16888_ (_08597_, _08533_, _08596_);
  and _16889_ (_08598_, _08026_, word_in[4]);
  and _16890_ (_08599_, _08598_, _08533_);
  or _16891_ (_08600_, _08599_, _08597_);
  or _16892_ (_08601_, _08600_, _08528_);
  or _16893_ (_08602_, _08529_, word_in[12]);
  and _16894_ (_08603_, _08602_, _08601_);
  or _16895_ (_08604_, _08603_, _08526_);
  nor _16896_ (_08605_, _08527_, word_in[20]);
  nor _16897_ (_08606_, _08605_, _08543_);
  and _16898_ (_08607_, _08606_, _08604_);
  and _16899_ (_08608_, _08010_, word_in[28]);
  and _16900_ (_08609_, _08608_, _08543_);
  or _16901_ (_07465_, _08609_, _08607_);
  not _16902_ (_08610_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _16903_ (_08611_, _08533_, _08610_);
  and _16904_ (_08612_, _08026_, word_in[5]);
  and _16905_ (_08613_, _08612_, _08533_);
  or _16906_ (_08614_, _08613_, _08611_);
  or _16907_ (_08615_, _08614_, _08528_);
  or _16908_ (_08616_, _08529_, word_in[13]);
  and _16909_ (_08617_, _08616_, _08615_);
  or _16910_ (_08618_, _08617_, _08526_);
  nor _16911_ (_08619_, _08527_, word_in[21]);
  nor _16912_ (_08620_, _08619_, _08543_);
  and _16913_ (_08621_, _08620_, _08618_);
  and _16914_ (_08622_, _08010_, word_in[29]);
  and _16915_ (_08623_, _08622_, _08543_);
  or _16916_ (_07470_, _08623_, _08621_);
  and _16917_ (_08624_, _08010_, word_in[30]);
  and _16918_ (_08625_, _08624_, _08543_);
  not _16919_ (_08626_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _16920_ (_08627_, _08533_, _08626_);
  and _16921_ (_08628_, _08026_, word_in[6]);
  and _16922_ (_08629_, _08628_, _08533_);
  or _16923_ (_08630_, _08629_, _08627_);
  or _16924_ (_08631_, _08630_, _08528_);
  or _16925_ (_08632_, _08529_, word_in[14]);
  and _16926_ (_08633_, _08632_, _08631_);
  or _16927_ (_08634_, _08633_, _08526_);
  nor _16928_ (_08635_, _08527_, word_in[22]);
  nor _16929_ (_08636_, _08635_, _08543_);
  and _16930_ (_08637_, _08636_, _08634_);
  or _16931_ (_07475_, _08637_, _08625_);
  nor _16932_ (_08638_, _08533_, _07839_);
  and _16933_ (_08639_, _08533_, _08029_);
  or _16934_ (_08640_, _08639_, _08638_);
  or _16935_ (_08641_, _08640_, _08528_);
  not _16936_ (_08642_, word_in[15]);
  nand _16937_ (_08643_, _08528_, _08642_);
  and _16938_ (_08644_, _08643_, _08641_);
  or _16939_ (_08645_, _08644_, _08526_);
  or _16940_ (_08646_, _08527_, word_in[23]);
  and _16941_ (_08647_, _08646_, _08548_);
  and _16942_ (_08648_, _08647_, _08645_);
  and _16943_ (_08649_, _08543_, word_in[31]);
  or _16944_ (_07477_, _08649_, _08648_);
  and _16945_ (_08650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _16946_ (_08651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _16947_ (_08652_, _05626_, _08651_);
  not _16948_ (_08653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _16949_ (_08654_, _08653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _16950_ (_08655_, _08654_, _08652_);
  nor _16951_ (_08656_, _08655_, _08650_);
  or _16952_ (_08657_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _16953_ (_08658_, _08657_, _05141_);
  nor _16954_ (_07493_, _08658_, _08656_);
  and _16955_ (_08659_, _08010_, _08043_);
  not _16956_ (_08660_, _08659_);
  and _16957_ (_08661_, _08016_, _07765_);
  and _16958_ (_08662_, _08661_, _07891_);
  not _16959_ (_08663_, _08662_);
  and _16960_ (_08664_, _08021_, _07761_);
  and _16961_ (_08665_, _08664_, _07781_);
  and _16962_ (_08666_, _08026_, word_in[0]);
  and _16963_ (_08667_, _08026_, _08057_);
  and _16964_ (_08668_, _08024_, _07634_);
  not _16965_ (_08669_, _08668_);
  nor _16966_ (_08670_, _08669_, _08667_);
  and _16967_ (_08671_, _08670_, _08666_);
  not _16968_ (_08672_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _16969_ (_08673_, _08670_, _08672_);
  nor _16970_ (_08674_, _08673_, _08671_);
  nor _16971_ (_08675_, _08674_, _08665_);
  and _16972_ (_08676_, _08665_, word_in[8]);
  or _16973_ (_08677_, _08676_, _08675_);
  and _16974_ (_08678_, _08677_, _08663_);
  and _16975_ (_08680_, _08662_, _08544_);
  or _16976_ (_08681_, _08680_, _08678_);
  and _16977_ (_08683_, _08681_, _08660_);
  and _16978_ (_08684_, _08659_, word_in[24]);
  or _16979_ (_07553_, _08684_, _08683_);
  not _16980_ (_08685_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _16981_ (_08686_, _08670_, _08685_);
  and _16982_ (_08687_, _08670_, _08556_);
  nor _16983_ (_08688_, _08687_, _08686_);
  nor _16984_ (_08689_, _08688_, _08665_);
  and _16985_ (_08690_, _08665_, word_in[9]);
  or _16986_ (_08692_, _08690_, _08689_);
  and _16987_ (_08693_, _08692_, _08663_);
  and _16988_ (_08694_, _08016_, word_in[17]);
  and _16989_ (_08695_, _08662_, _08694_);
  or _16990_ (_08696_, _08695_, _08693_);
  and _16991_ (_08697_, _08696_, _08660_);
  and _16992_ (_08698_, _08659_, word_in[25]);
  or _16993_ (_07558_, _08698_, _08697_);
  and _16994_ (_08699_, _08670_, _08572_);
  not _16995_ (_08700_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _16996_ (_08701_, _08670_, _08700_);
  nor _16997_ (_08702_, _08701_, _08699_);
  nor _16998_ (_08703_, _08702_, _08665_);
  and _16999_ (_08704_, _08665_, word_in[10]);
  or _17000_ (_08705_, _08704_, _08703_);
  and _17001_ (_08706_, _08705_, _08663_);
  and _17002_ (_08707_, _08016_, word_in[18]);
  and _17003_ (_08708_, _08662_, _08707_);
  or _17004_ (_08709_, _08708_, _08706_);
  and _17005_ (_08710_, _08709_, _08660_);
  and _17006_ (_08711_, _08659_, word_in[26]);
  or _17007_ (_07562_, _08711_, _08710_);
  and _17008_ (_08712_, _08016_, word_in[19]);
  and _17009_ (_08713_, _08662_, _08712_);
  not _17010_ (_08714_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _17011_ (_08715_, _08670_, _08714_);
  and _17012_ (_08716_, _08670_, _08586_);
  nor _17013_ (_08717_, _08716_, _08715_);
  nor _17014_ (_08718_, _08717_, _08665_);
  and _17015_ (_08719_, _08665_, word_in[11]);
  or _17016_ (_08720_, _08719_, _08718_);
  and _17017_ (_08721_, _08720_, _08663_);
  or _17018_ (_08722_, _08721_, _08713_);
  and _17019_ (_08723_, _08722_, _08660_);
  and _17020_ (_08724_, _08659_, word_in[27]);
  or _17021_ (_07565_, _08724_, _08723_);
  and _17022_ (_08725_, _08670_, _08598_);
  not _17023_ (_08726_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _17024_ (_08727_, _08670_, _08726_);
  nor _17025_ (_08728_, _08727_, _08725_);
  nor _17026_ (_08729_, _08728_, _08665_);
  and _17027_ (_08730_, _08665_, word_in[12]);
  or _17028_ (_08731_, _08730_, _08729_);
  and _17029_ (_08732_, _08731_, _08663_);
  and _17030_ (_08733_, _08016_, word_in[20]);
  and _17031_ (_08734_, _08662_, _08733_);
  or _17032_ (_08735_, _08734_, _08732_);
  and _17033_ (_08736_, _08735_, _08660_);
  and _17034_ (_08737_, _08659_, word_in[28]);
  or _17035_ (_07569_, _08737_, _08736_);
  and _17036_ (_08738_, _08670_, _08612_);
  not _17037_ (_08739_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _17038_ (_08740_, _08670_, _08739_);
  nor _17039_ (_08741_, _08740_, _08738_);
  nor _17040_ (_08742_, _08741_, _08665_);
  and _17041_ (_08743_, _08665_, word_in[13]);
  or _17042_ (_08744_, _08743_, _08742_);
  and _17043_ (_08745_, _08744_, _08663_);
  and _17044_ (_08746_, _08016_, word_in[21]);
  and _17045_ (_08747_, _08662_, _08746_);
  or _17046_ (_08748_, _08747_, _08745_);
  and _17047_ (_08749_, _08748_, _08660_);
  and _17048_ (_08750_, _08659_, word_in[29]);
  or _17049_ (_07573_, _08750_, _08749_);
  and _17050_ (_08751_, _08670_, _08628_);
  not _17051_ (_08752_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _17052_ (_08753_, _08670_, _08752_);
  nor _17053_ (_08754_, _08753_, _08751_);
  nor _17054_ (_08755_, _08754_, _08665_);
  and _17055_ (_08756_, _08665_, word_in[14]);
  or _17056_ (_08757_, _08756_, _08755_);
  and _17057_ (_08758_, _08757_, _08663_);
  and _17058_ (_08759_, _08016_, word_in[22]);
  and _17059_ (_08760_, _08662_, _08759_);
  or _17060_ (_08761_, _08760_, _08758_);
  and _17061_ (_08762_, _08761_, _08660_);
  and _17062_ (_08763_, _08659_, word_in[30]);
  or _17063_ (_07575_, _08763_, _08762_);
  nor _17064_ (_08764_, _08670_, _07746_);
  and _17065_ (_08765_, _08670_, _08029_);
  or _17066_ (_08766_, _08765_, _08764_);
  or _17067_ (_08767_, _08766_, _08665_);
  nand _17068_ (_08768_, _08665_, _08642_);
  and _17069_ (_08769_, _08768_, _08767_);
  or _17070_ (_08771_, _08769_, _08662_);
  or _17071_ (_08772_, _08663_, _08037_);
  and _17072_ (_08773_, _08772_, _08660_);
  and _17073_ (_08774_, _08773_, _08771_);
  and _17074_ (_08776_, _08659_, word_in[31]);
  or _17075_ (_07578_, _08776_, _08774_);
  and _17076_ (_08778_, _08016_, _07761_);
  and _17077_ (_08779_, _08778_, _07891_);
  not _17078_ (_08780_, _08779_);
  and _17079_ (_08782_, _08021_, _07788_);
  and _17080_ (_08783_, _08782_, _07781_);
  not _17081_ (_08784_, _08024_);
  and _17082_ (_08786_, _08530_, _08784_);
  and _17083_ (_08787_, _08786_, _08081_);
  and _17084_ (_08789_, _08787_, _08666_);
  not _17085_ (_08790_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _17086_ (_08791_, _08787_, _08790_);
  nor _17087_ (_08793_, _08791_, _08789_);
  nor _17088_ (_08794_, _08793_, _08783_);
  and _17089_ (_08795_, _08783_, word_in[8]);
  or _17090_ (_08797_, _08795_, _08794_);
  and _17091_ (_08798_, _08797_, _08780_);
  and _17092_ (_08799_, _08010_, _07765_);
  and _17093_ (_08800_, _08799_, _07947_);
  and _17094_ (_08801_, _08779_, _08544_);
  or _17095_ (_08802_, _08801_, _08800_);
  or _17096_ (_08803_, _08802_, _08798_);
  not _17097_ (_08804_, _08800_);
  or _17098_ (_08805_, _08804_, word_in[24]);
  and _17099_ (_07655_, _08805_, _08803_);
  and _17100_ (_08806_, _05563_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _17101_ (_08807_, _06004_, _05523_);
  or _17102_ (_08808_, _08807_, _08806_);
  and _17103_ (_07658_, _08808_, _05141_);
  and _17104_ (_08809_, _08787_, _08556_);
  not _17105_ (_08810_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _17106_ (_08811_, _08787_, _08810_);
  nor _17107_ (_08812_, _08811_, _08809_);
  nor _17108_ (_08813_, _08812_, _08783_);
  and _17109_ (_08814_, _08783_, word_in[9]);
  or _17110_ (_08815_, _08814_, _08813_);
  and _17111_ (_08816_, _08815_, _08780_);
  and _17112_ (_08817_, _08779_, _08694_);
  or _17113_ (_08818_, _08817_, _08800_);
  or _17114_ (_08819_, _08818_, _08816_);
  or _17115_ (_08820_, _08804_, word_in[25]);
  and _17116_ (_07660_, _08820_, _08819_);
  and _17117_ (_08822_, _08787_, _08572_);
  not _17118_ (_08823_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _17119_ (_08824_, _08787_, _08823_);
  nor _17120_ (_08825_, _08824_, _08822_);
  nor _17121_ (_08826_, _08825_, _08783_);
  and _17122_ (_08827_, _08783_, word_in[10]);
  or _17123_ (_08828_, _08827_, _08826_);
  and _17124_ (_08829_, _08828_, _08780_);
  and _17125_ (_08830_, _08779_, word_in[18]);
  or _17126_ (_08831_, _08830_, _08800_);
  or _17127_ (_08832_, _08831_, _08829_);
  or _17128_ (_08833_, _08804_, word_in[26]);
  and _17129_ (_07664_, _08833_, _08832_);
  and _17130_ (_08834_, _08779_, word_in[19]);
  and _17131_ (_08835_, _08787_, _08586_);
  not _17132_ (_08836_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _17133_ (_08837_, _08787_, _08836_);
  nor _17134_ (_08838_, _08837_, _08835_);
  nor _17135_ (_08839_, _08838_, _08783_);
  and _17136_ (_08840_, _08783_, word_in[11]);
  or _17137_ (_08841_, _08840_, _08839_);
  and _17138_ (_08842_, _08841_, _08780_);
  or _17139_ (_08843_, _08842_, _08834_);
  and _17140_ (_08844_, _08843_, _08804_);
  and _17141_ (_08845_, _08800_, word_in[27]);
  or _17142_ (_07667_, _08845_, _08844_);
  and _17143_ (_08846_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _17144_ (_08847_, _06004_, _05617_);
  or _17145_ (_08848_, _08847_, _08846_);
  and _17146_ (_07670_, _08848_, _05141_);
  and _17147_ (_08849_, _08787_, _08598_);
  not _17148_ (_08850_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _17149_ (_08851_, _08787_, _08850_);
  nor _17150_ (_08852_, _08851_, _08849_);
  nor _17151_ (_08853_, _08852_, _08783_);
  and _17152_ (_08854_, _08783_, word_in[12]);
  or _17153_ (_08855_, _08854_, _08853_);
  and _17154_ (_08856_, _08855_, _08780_);
  and _17155_ (_08857_, _08779_, word_in[20]);
  or _17156_ (_08858_, _08857_, _08800_);
  or _17157_ (_08860_, _08858_, _08856_);
  or _17158_ (_08861_, _08804_, word_in[28]);
  and _17159_ (_07672_, _08861_, _08860_);
  not _17160_ (_08862_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _17161_ (_08863_, _08787_, _08862_);
  and _17162_ (_08864_, _08787_, _08612_);
  or _17163_ (_08865_, _08864_, _08863_);
  or _17164_ (_08866_, _08865_, _08783_);
  not _17165_ (_08868_, _08783_);
  or _17166_ (_08869_, _08868_, word_in[13]);
  and _17167_ (_08871_, _08869_, _08866_);
  or _17168_ (_08872_, _08871_, _08779_);
  or _17169_ (_08874_, _08780_, word_in[21]);
  and _17170_ (_08875_, _08874_, _08804_);
  and _17171_ (_08876_, _08875_, _08872_);
  and _17172_ (_08878_, _08800_, word_in[29]);
  or _17173_ (_07677_, _08878_, _08876_);
  and _17174_ (_08880_, _05614_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand _17175_ (_08881_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor _17176_ (_08883_, _08881_, _05609_);
  and _17177_ (_08884_, _05605_, _05283_);
  or _17178_ (_08885_, _08884_, _08883_);
  or _17179_ (_08886_, _08885_, _08880_);
  and _17180_ (_07680_, _08886_, _05141_);
  and _17181_ (_08888_, _08787_, _08628_);
  not _17182_ (_08890_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _17183_ (_08891_, _08787_, _08890_);
  nor _17184_ (_08892_, _08891_, _08888_);
  nor _17185_ (_08893_, _08892_, _08783_);
  and _17186_ (_08894_, _08783_, word_in[14]);
  or _17187_ (_08895_, _08894_, _08893_);
  and _17188_ (_08896_, _08895_, _08780_);
  and _17189_ (_08897_, _08779_, _08759_);
  or _17190_ (_08898_, _08897_, _08800_);
  or _17191_ (_08899_, _08898_, _08896_);
  or _17192_ (_08900_, _08804_, word_in[30]);
  and _17193_ (_07682_, _08900_, _08899_);
  and _17194_ (_08901_, _08787_, _08029_);
  nor _17195_ (_08902_, _08787_, _07834_);
  or _17196_ (_08903_, _08902_, _08901_);
  or _17197_ (_08904_, _08903_, _08783_);
  nand _17198_ (_08905_, _08783_, _08642_);
  and _17199_ (_08906_, _08905_, _08780_);
  and _17200_ (_08907_, _08906_, _08904_);
  and _17201_ (_08908_, _08779_, _08037_);
  or _17202_ (_08909_, _08908_, _08800_);
  or _17203_ (_08910_, _08909_, _08907_);
  or _17204_ (_08911_, _08804_, word_in[31]);
  and _17205_ (_07687_, _08911_, _08910_);
  or _17206_ (_08912_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand _17207_ (_08913_, _07619_, _06399_);
  and _17208_ (_08914_, _08913_, _05141_);
  and _17209_ (_07749_, _08914_, _08912_);
  and _17210_ (_08915_, _08010_, _08071_);
  not _17211_ (_08916_, _08915_);
  and _17212_ (_08917_, _08016_, _07788_);
  and _17213_ (_08918_, _08917_, _07891_);
  not _17214_ (_08919_, _08918_);
  and _17215_ (_08920_, _08022_, _07781_);
  not _17216_ (_08921_, _08025_);
  nor _17217_ (_08922_, _08667_, _08921_);
  and _17218_ (_08923_, _08922_, _08666_);
  not _17219_ (_08924_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _17220_ (_08925_, _08922_, _08924_);
  nor _17221_ (_08926_, _08925_, _08923_);
  nor _17222_ (_08927_, _08926_, _08920_);
  and _17223_ (_08928_, _08920_, word_in[8]);
  or _17224_ (_08929_, _08928_, _08927_);
  and _17225_ (_08930_, _08929_, _08919_);
  and _17226_ (_08931_, _08918_, word_in[16]);
  or _17227_ (_08932_, _08931_, _08930_);
  and _17228_ (_08933_, _08932_, _08916_);
  and _17229_ (_08934_, _08915_, word_in[24]);
  or _17230_ (_07755_, _08934_, _08933_);
  and _17231_ (_08935_, _08918_, word_in[17]);
  and _17232_ (_08936_, _08922_, _08556_);
  not _17233_ (_08937_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _17234_ (_08938_, _08922_, _08937_);
  nor _17235_ (_08939_, _08938_, _08936_);
  nor _17236_ (_08940_, _08939_, _08920_);
  and _17237_ (_08941_, _08920_, word_in[9]);
  or _17238_ (_08942_, _08941_, _08940_);
  and _17239_ (_08943_, _08942_, _08919_);
  or _17240_ (_08944_, _08943_, _08935_);
  and _17241_ (_08945_, _08944_, _08916_);
  and _17242_ (_08946_, _08915_, word_in[25]);
  or _17243_ (_07760_, _08946_, _08945_);
  and _17244_ (_08947_, _08915_, word_in[26]);
  and _17245_ (_08948_, _08922_, _08572_);
  not _17246_ (_08949_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _17247_ (_08950_, _08922_, _08949_);
  nor _17248_ (_08951_, _08950_, _08948_);
  nor _17249_ (_08952_, _08951_, _08920_);
  and _17250_ (_08953_, _08920_, word_in[10]);
  or _17251_ (_08954_, _08953_, _08952_);
  or _17252_ (_08955_, _08954_, _08918_);
  or _17253_ (_08956_, _08919_, _08707_);
  and _17254_ (_08957_, _08956_, _08916_);
  and _17255_ (_08958_, _08957_, _08955_);
  or _17256_ (_07762_, _08958_, _08947_);
  and _17257_ (_08959_, _08922_, _08586_);
  not _17258_ (_08960_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _17259_ (_08961_, _08922_, _08960_);
  nor _17260_ (_08962_, _08961_, _08959_);
  nor _17261_ (_08963_, _08962_, _08920_);
  and _17262_ (_08964_, _08920_, word_in[11]);
  or _17263_ (_08965_, _08964_, _08963_);
  and _17264_ (_08966_, _08965_, _08919_);
  and _17265_ (_08967_, _08918_, word_in[19]);
  or _17266_ (_08968_, _08967_, _08915_);
  or _17267_ (_08969_, _08968_, _08966_);
  or _17268_ (_08970_, _08916_, word_in[27]);
  and _17269_ (_07764_, _08970_, _08969_);
  and _17270_ (_08971_, _08922_, _08598_);
  not _17271_ (_08972_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _17272_ (_08973_, _08922_, _08972_);
  nor _17273_ (_08974_, _08973_, _08971_);
  nor _17274_ (_08975_, _08974_, _08920_);
  and _17275_ (_08976_, _08920_, word_in[12]);
  or _17276_ (_08977_, _08976_, _08975_);
  and _17277_ (_08978_, _08977_, _08919_);
  and _17278_ (_08979_, _08918_, word_in[20]);
  or _17279_ (_08980_, _08979_, _08915_);
  or _17280_ (_08981_, _08980_, _08978_);
  or _17281_ (_08982_, _08916_, word_in[28]);
  and _17282_ (_07767_, _08982_, _08981_);
  and _17283_ (_08983_, _08922_, _08612_);
  not _17284_ (_08984_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _17285_ (_08985_, _08922_, _08984_);
  nor _17286_ (_08986_, _08985_, _08983_);
  nor _17287_ (_08987_, _08986_, _08920_);
  and _17288_ (_08988_, _08920_, word_in[13]);
  or _17289_ (_08989_, _08988_, _08987_);
  and _17290_ (_08990_, _08989_, _08919_);
  and _17291_ (_08992_, _08918_, _08746_);
  or _17292_ (_08993_, _08992_, _08915_);
  or _17293_ (_08994_, _08993_, _08990_);
  or _17294_ (_08995_, _08916_, word_in[29]);
  and _17295_ (_07770_, _08995_, _08994_);
  and _17296_ (_08996_, _08915_, word_in[30]);
  and _17297_ (_08997_, _08922_, _08628_);
  not _17298_ (_08998_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _17299_ (_08999_, _08922_, _08998_);
  nor _17300_ (_09000_, _08999_, _08997_);
  nor _17301_ (_09001_, _09000_, _08920_);
  and _17302_ (_09002_, _08920_, word_in[14]);
  or _17303_ (_09003_, _09002_, _09001_);
  or _17304_ (_09004_, _09003_, _08918_);
  or _17305_ (_09005_, _08919_, _08759_);
  and _17306_ (_09006_, _09005_, _08916_);
  and _17307_ (_09007_, _09006_, _09004_);
  or _17308_ (_07775_, _09007_, _08996_);
  nor _17309_ (_09008_, _08922_, _07730_);
  and _17310_ (_09009_, _08922_, _08029_);
  or _17311_ (_09010_, _09009_, _09008_);
  or _17312_ (_09011_, _09010_, _08920_);
  nand _17313_ (_09012_, _08920_, _08642_);
  and _17314_ (_09013_, _09012_, _09011_);
  or _17315_ (_09014_, _09013_, _08918_);
  or _17316_ (_09015_, _08919_, _08037_);
  and _17317_ (_09016_, _09015_, _08916_);
  and _17318_ (_09017_, _09016_, _09014_);
  and _17319_ (_09018_, _08915_, word_in[31]);
  or _17320_ (_07778_, _09018_, _09017_);
  and _17321_ (_09019_, _08017_, _07927_);
  and _17322_ (_09020_, _09019_, _07798_);
  not _17323_ (_09021_, _09020_);
  and _17324_ (_09022_, _08021_, _08064_);
  not _17325_ (_09023_, _09022_);
  or _17326_ (_09024_, _09023_, word_in[8]);
  not _17327_ (_09025_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _17328_ (_09026_, _08026_, _07777_);
  and _17329_ (_09027_, _09026_, _08531_);
  nor _17330_ (_09028_, _09027_, _09025_);
  and _17331_ (_09029_, _09027_, word_in[0]);
  or _17332_ (_09030_, _09029_, _09028_);
  or _17333_ (_09031_, _09030_, _09022_);
  and _17334_ (_09032_, _09031_, _09024_);
  and _17335_ (_09033_, _09032_, _09021_);
  and _17336_ (_09034_, _08010_, _07941_);
  and _17337_ (_09035_, _09034_, _07946_);
  and _17338_ (_09036_, _09035_, _07788_);
  and _17339_ (_09037_, _09020_, _08544_);
  or _17340_ (_09038_, _09037_, _09036_);
  or _17341_ (_09039_, _09038_, _09033_);
  and _17342_ (_09040_, _08010_, word_in[24]);
  not _17343_ (_09041_, _09036_);
  or _17344_ (_09042_, _09041_, _09040_);
  and _17345_ (_07863_, _09042_, _09039_);
  not _17346_ (_09043_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _17347_ (_09044_, _09027_, _09043_);
  and _17348_ (_09045_, _09027_, word_in[1]);
  or _17349_ (_09046_, _09045_, _09044_);
  and _17350_ (_09047_, _09046_, _09023_);
  and _17351_ (_09048_, _09022_, word_in[9]);
  or _17352_ (_09049_, _09048_, _09047_);
  and _17353_ (_09050_, _09049_, _09021_);
  and _17354_ (_09051_, _09020_, _08694_);
  or _17355_ (_09052_, _09051_, _09036_);
  or _17356_ (_09053_, _09052_, _09050_);
  or _17357_ (_09054_, _09041_, _08566_);
  and _17358_ (_07866_, _09054_, _09053_);
  not _17359_ (_09055_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _17360_ (_09056_, _09027_, _09055_);
  and _17361_ (_09057_, _09027_, word_in[2]);
  or _17362_ (_09058_, _09057_, _09056_);
  or _17363_ (_09059_, _09058_, _09022_);
  or _17364_ (_09060_, _09023_, word_in[10]);
  and _17365_ (_09061_, _09060_, _09059_);
  and _17366_ (_09062_, _09061_, _09021_);
  and _17367_ (_09063_, _09020_, _08707_);
  or _17368_ (_09064_, _09063_, _09036_);
  or _17369_ (_09065_, _09064_, _09062_);
  or _17370_ (_09066_, _09041_, _08568_);
  and _17371_ (_07869_, _09066_, _09065_);
  not _17372_ (_09067_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _17373_ (_09068_, _09027_, _09067_);
  and _17374_ (_09069_, _09027_, word_in[3]);
  or _17375_ (_09070_, _09069_, _09068_);
  and _17376_ (_09071_, _09070_, _09023_);
  and _17377_ (_09072_, _09022_, word_in[11]);
  or _17378_ (_09073_, _09072_, _09071_);
  and _17379_ (_09074_, _09073_, _09021_);
  and _17380_ (_09075_, _09020_, _08712_);
  or _17381_ (_09076_, _09075_, _09036_);
  or _17382_ (_09077_, _09076_, _09074_);
  or _17383_ (_09078_, _09041_, _08582_);
  and _17384_ (_07873_, _09078_, _09077_);
  not _17385_ (_09079_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _17386_ (_09080_, _09027_, _09079_);
  and _17387_ (_09081_, _09027_, word_in[4]);
  or _17388_ (_09082_, _09081_, _09080_);
  or _17389_ (_09083_, _09082_, _09022_);
  or _17390_ (_09084_, _09023_, word_in[12]);
  and _17391_ (_09085_, _09084_, _09083_);
  and _17392_ (_09086_, _09085_, _09021_);
  and _17393_ (_09087_, _09020_, _08733_);
  or _17394_ (_09088_, _09087_, _09036_);
  or _17395_ (_09089_, _09088_, _09086_);
  or _17396_ (_09090_, _09041_, _08608_);
  and _17397_ (_07876_, _09090_, _09089_);
  not _17398_ (_09091_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _17399_ (_09092_, _09027_, _09091_);
  and _17400_ (_09093_, _09027_, word_in[5]);
  or _17401_ (_09094_, _09093_, _09092_);
  and _17402_ (_09095_, _09094_, _09023_);
  and _17403_ (_09096_, _09022_, word_in[13]);
  or _17404_ (_09097_, _09096_, _09095_);
  and _17405_ (_09098_, _09097_, _09021_);
  and _17406_ (_09099_, _09020_, _08746_);
  or _17407_ (_09100_, _09099_, _09036_);
  or _17408_ (_09101_, _09100_, _09098_);
  or _17409_ (_09102_, _09041_, _08622_);
  and _17410_ (_07879_, _09102_, _09101_);
  not _17411_ (_09103_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _17412_ (_09104_, _09027_, _09103_);
  and _17413_ (_09105_, _09027_, word_in[6]);
  or _17414_ (_09106_, _09105_, _09104_);
  and _17415_ (_09107_, _09106_, _09023_);
  and _17416_ (_09108_, _09022_, word_in[14]);
  or _17417_ (_09110_, _09108_, _09107_);
  and _17418_ (_09111_, _09110_, _09021_);
  and _17419_ (_09112_, _09020_, _08759_);
  or _17420_ (_09113_, _09112_, _09036_);
  or _17421_ (_09114_, _09113_, _09111_);
  or _17422_ (_09115_, _09041_, _08624_);
  and _17423_ (_07881_, _09115_, _09114_);
  nor _17424_ (_09116_, _09027_, _07851_);
  and _17425_ (_09117_, _09027_, word_in[7]);
  or _17426_ (_09118_, _09117_, _09116_);
  and _17427_ (_09120_, _09118_, _09023_);
  and _17428_ (_09121_, _09022_, word_in[15]);
  or _17429_ (_09122_, _09121_, _09120_);
  and _17430_ (_09123_, _09122_, _09021_);
  and _17431_ (_09124_, _09020_, _08037_);
  or _17432_ (_09125_, _09124_, _09036_);
  or _17433_ (_09126_, _09125_, _09123_);
  or _17434_ (_09127_, _09041_, _08011_);
  and _17435_ (_07885_, _09127_, _09126_);
  and _17436_ (_09128_, _08664_, _07807_);
  not _17437_ (_09129_, _09128_);
  or _17438_ (_09130_, _09129_, word_in[8]);
  and _17439_ (_09131_, _09019_, _07765_);
  not _17440_ (_09132_, _09131_);
  not _17441_ (_09133_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _17442_ (_09134_, _09026_, _08668_);
  nor _17443_ (_09135_, _09134_, _09133_);
  and _17444_ (_09136_, _09134_, word_in[0]);
  or _17445_ (_09137_, _09136_, _09135_);
  or _17446_ (_09138_, _09137_, _09128_);
  and _17447_ (_09139_, _09138_, _09132_);
  and _17448_ (_09140_, _09139_, _09130_);
  and _17449_ (_09141_, _09035_, _07798_);
  and _17450_ (_09142_, _09131_, _08544_);
  or _17451_ (_09144_, _09142_, _09141_);
  or _17452_ (_09145_, _09144_, _09140_);
  not _17453_ (_09146_, _09141_);
  or _17454_ (_09147_, _09146_, word_in[24]);
  and _17455_ (_07953_, _09147_, _09145_);
  and _17456_ (_09148_, _09131_, _08694_);
  and _17457_ (_09149_, _09134_, word_in[1]);
  not _17458_ (_09150_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _17459_ (_09151_, _09134_, _09150_);
  nor _17460_ (_09152_, _09151_, _09149_);
  nor _17461_ (_09153_, _09152_, _09128_);
  and _17462_ (_09154_, _09128_, word_in[9]);
  or _17463_ (_09155_, _09154_, _09153_);
  and _17464_ (_09156_, _09155_, _09132_);
  or _17465_ (_09157_, _09156_, _09148_);
  and _17466_ (_09158_, _09157_, _09146_);
  and _17467_ (_09159_, _09141_, word_in[25]);
  or _17468_ (_07957_, _09159_, _09158_);
  or _17469_ (_09160_, _09132_, _08707_);
  not _17470_ (_09161_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _17471_ (_09162_, _09134_, _09161_);
  and _17472_ (_09163_, _09134_, word_in[2]);
  or _17473_ (_09164_, _09163_, _09162_);
  or _17474_ (_09165_, _09164_, _09128_);
  or _17475_ (_09166_, _09129_, word_in[10]);
  and _17476_ (_09167_, _09166_, _09165_);
  or _17477_ (_09168_, _09167_, _09131_);
  and _17478_ (_09169_, _09168_, _09160_);
  and _17479_ (_09171_, _09169_, _09146_);
  and _17480_ (_09172_, _09141_, word_in[26]);
  or _17481_ (_07961_, _09172_, _09171_);
  or _17482_ (_09174_, _09132_, _08712_);
  not _17483_ (_09175_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _17484_ (_09176_, _09134_, _09175_);
  and _17485_ (_09177_, _09134_, word_in[3]);
  or _17486_ (_09178_, _09177_, _09176_);
  or _17487_ (_09179_, _09178_, _09128_);
  or _17488_ (_09180_, _09129_, word_in[11]);
  and _17489_ (_09181_, _09180_, _09179_);
  or _17490_ (_09182_, _09181_, _09131_);
  and _17491_ (_09183_, _09182_, _09174_);
  or _17492_ (_09184_, _09183_, _09141_);
  or _17493_ (_09185_, _09146_, word_in[27]);
  and _17494_ (_07965_, _09185_, _09184_);
  not _17495_ (_09186_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _17496_ (_09187_, _09134_, _09186_);
  and _17497_ (_09188_, _09134_, word_in[4]);
  nor _17498_ (_09189_, _09188_, _09187_);
  nor _17499_ (_09190_, _09189_, _09128_);
  and _17500_ (_09191_, _09128_, word_in[12]);
  or _17501_ (_09192_, _09191_, _09190_);
  and _17502_ (_09193_, _09192_, _09132_);
  and _17503_ (_09194_, _09131_, _08733_);
  or _17504_ (_09195_, _09194_, _09141_);
  or _17505_ (_09196_, _09195_, _09193_);
  or _17506_ (_09197_, _09146_, word_in[28]);
  and _17507_ (_07969_, _09197_, _09196_);
  not _17508_ (_09198_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _17509_ (_09199_, _09134_, _09198_);
  and _17510_ (_09200_, _09134_, word_in[5]);
  nor _17511_ (_09201_, _09200_, _09199_);
  nor _17512_ (_09202_, _09201_, _09128_);
  and _17513_ (_09203_, _09128_, word_in[13]);
  or _17514_ (_09204_, _09203_, _09202_);
  and _17515_ (_09205_, _09204_, _09132_);
  and _17516_ (_09206_, _09131_, _08746_);
  or _17517_ (_09207_, _09206_, _09141_);
  or _17518_ (_09208_, _09207_, _09205_);
  or _17519_ (_09209_, _09146_, word_in[29]);
  and _17520_ (_07971_, _09209_, _09208_);
  or _17521_ (_09210_, _09132_, _08759_);
  not _17522_ (_09211_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _17523_ (_09212_, _09134_, _09211_);
  and _17524_ (_09213_, _09134_, word_in[6]);
  or _17525_ (_09214_, _09213_, _09212_);
  or _17526_ (_09215_, _09214_, _09128_);
  or _17527_ (_09216_, _09129_, word_in[14]);
  and _17528_ (_09217_, _09216_, _09215_);
  or _17529_ (_09218_, _09217_, _09131_);
  and _17530_ (_09219_, _09218_, _09210_);
  and _17531_ (_09220_, _09219_, _09146_);
  and _17532_ (_09221_, _09141_, word_in[30]);
  or _17533_ (_07974_, _09221_, _09220_);
  or _17534_ (_09222_, _09132_, _08037_);
  nor _17535_ (_09223_, _09134_, _07741_);
  and _17536_ (_09224_, _09134_, word_in[7]);
  or _17537_ (_09225_, _09224_, _09223_);
  or _17538_ (_09226_, _09225_, _09128_);
  nand _17539_ (_09227_, _09128_, _08642_);
  and _17540_ (_09228_, _09227_, _09226_);
  or _17541_ (_09229_, _09228_, _09131_);
  and _17542_ (_09230_, _09229_, _09222_);
  and _17543_ (_09231_, _09230_, _09146_);
  and _17544_ (_09232_, _09141_, word_in[31]);
  or _17545_ (_07976_, _09232_, _09231_);
  and _17546_ (_09233_, _09035_, _07765_);
  and _17547_ (_09234_, _09019_, _07761_);
  and _17548_ (_09235_, _08782_, _07807_);
  not _17549_ (_09236_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _17550_ (_09237_, _08786_, _07777_);
  nor _17551_ (_09238_, _09237_, _09236_);
  and _17552_ (_09239_, _09237_, _08666_);
  or _17553_ (_09240_, _09239_, _09238_);
  or _17554_ (_09241_, _09240_, _09235_);
  not _17555_ (_09242_, _09235_);
  or _17556_ (_09243_, _09242_, word_in[8]);
  and _17557_ (_09244_, _09243_, _09241_);
  or _17558_ (_09245_, _09244_, _09234_);
  not _17559_ (_09246_, _09234_);
  or _17560_ (_09247_, _09246_, _08544_);
  and _17561_ (_09248_, _09247_, _09245_);
  or _17562_ (_09249_, _09248_, _09233_);
  not _17563_ (_09250_, _09233_);
  or _17564_ (_09251_, _09250_, word_in[24]);
  and _17565_ (_08042_, _09251_, _09249_);
  and _17566_ (_09252_, _09237_, _08556_);
  not _17567_ (_09253_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _17568_ (_09254_, _09237_, _09253_);
  nor _17569_ (_09255_, _09254_, _09252_);
  nor _17570_ (_09256_, _09255_, _09235_);
  and _17571_ (_09257_, _09235_, word_in[9]);
  or _17572_ (_09258_, _09257_, _09256_);
  and _17573_ (_09259_, _09258_, _09246_);
  and _17574_ (_09260_, _09234_, _08694_);
  or _17575_ (_09261_, _09260_, _09233_);
  or _17576_ (_09262_, _09261_, _09259_);
  or _17577_ (_09263_, _09250_, word_in[25]);
  and _17578_ (_08045_, _09263_, _09262_);
  not _17579_ (_09264_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _17580_ (_09265_, _09237_, _09264_);
  and _17581_ (_09266_, _09237_, _08572_);
  or _17582_ (_09267_, _09266_, _09265_);
  or _17583_ (_09268_, _09267_, _09235_);
  or _17584_ (_09269_, _09242_, word_in[10]);
  and _17585_ (_09270_, _09269_, _09268_);
  or _17586_ (_09271_, _09270_, _09234_);
  or _17587_ (_09272_, _09246_, _08707_);
  and _17588_ (_09273_, _09272_, _09271_);
  and _17589_ (_09274_, _09273_, _09250_);
  and _17590_ (_09275_, _09233_, word_in[26]);
  or _17591_ (_08048_, _09275_, _09274_);
  not _17592_ (_09276_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _17593_ (_09277_, _09237_, _09276_);
  and _17594_ (_09278_, _09237_, _08586_);
  or _17595_ (_09279_, _09278_, _09277_);
  or _17596_ (_09280_, _09279_, _09235_);
  or _17597_ (_09281_, _09242_, word_in[11]);
  and _17598_ (_09282_, _09281_, _09280_);
  or _17599_ (_09283_, _09282_, _09234_);
  or _17600_ (_09284_, _09246_, _08712_);
  and _17601_ (_09285_, _09284_, _09283_);
  or _17602_ (_09286_, _09285_, _09233_);
  or _17603_ (_09287_, _09250_, word_in[27]);
  and _17604_ (_08051_, _09287_, _09286_);
  or _17605_ (_09288_, _09246_, _08733_);
  not _17606_ (_09289_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _17607_ (_09290_, _09237_, _09289_);
  and _17608_ (_09291_, _09237_, _08598_);
  or _17609_ (_09292_, _09291_, _09290_);
  or _17610_ (_09293_, _09292_, _09235_);
  or _17611_ (_09294_, _09242_, word_in[12]);
  and _17612_ (_09295_, _09294_, _09293_);
  or _17613_ (_09296_, _09295_, _09234_);
  and _17614_ (_09297_, _09296_, _09288_);
  or _17615_ (_09298_, _09297_, _09233_);
  or _17616_ (_09299_, _09250_, word_in[28]);
  and _17617_ (_08053_, _09299_, _09298_);
  and _17618_ (_09300_, _09237_, _08612_);
  not _17619_ (_09301_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _17620_ (_09302_, _09237_, _09301_);
  nor _17621_ (_09303_, _09302_, _09300_);
  nor _17622_ (_09304_, _09303_, _09235_);
  and _17623_ (_09305_, _09235_, word_in[13]);
  or _17624_ (_09306_, _09305_, _09304_);
  and _17625_ (_09307_, _09306_, _09246_);
  and _17626_ (_09308_, _09234_, _08746_);
  or _17627_ (_09309_, _09308_, _09307_);
  and _17628_ (_09310_, _09309_, _09250_);
  and _17629_ (_09311_, _09233_, word_in[29]);
  or _17630_ (_08056_, _09311_, _09310_);
  and _17631_ (_09312_, _09237_, _08628_);
  not _17632_ (_09313_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _17633_ (_09314_, _09237_, _09313_);
  nor _17634_ (_09315_, _09314_, _09312_);
  nor _17635_ (_09316_, _09315_, _09235_);
  and _17636_ (_09317_, _09235_, word_in[14]);
  or _17637_ (_09318_, _09317_, _09316_);
  and _17638_ (_09319_, _09318_, _09246_);
  and _17639_ (_09320_, _09234_, _08759_);
  or _17640_ (_09321_, _09320_, _09233_);
  or _17641_ (_09322_, _09321_, _09319_);
  or _17642_ (_09323_, _09250_, word_in[30]);
  and _17643_ (_08058_, _09323_, _09322_);
  nor _17644_ (_09324_, _09237_, _07846_);
  and _17645_ (_09325_, _09237_, _08029_);
  or _17646_ (_09326_, _09325_, _09324_);
  or _17647_ (_09327_, _09326_, _09235_);
  nand _17648_ (_09328_, _09235_, _08642_);
  and _17649_ (_09329_, _09328_, _09327_);
  or _17650_ (_09330_, _09329_, _09234_);
  or _17651_ (_09331_, _09246_, _08037_);
  and _17652_ (_09332_, _09331_, _09330_);
  or _17653_ (_09333_, _09332_, _09233_);
  or _17654_ (_09334_, _09250_, word_in[31]);
  and _17655_ (_08060_, _09334_, _09333_);
  and _17656_ (_09335_, _08010_, _08065_);
  and _17657_ (_09336_, _09335_, _09040_);
  not _17658_ (_09337_, _09335_);
  and _17659_ (_09338_, _09019_, _07788_);
  not _17660_ (_09339_, _09338_);
  and _17661_ (_09340_, _08022_, _07807_);
  and _17662_ (_09341_, _09026_, _08025_);
  and _17663_ (_09342_, _09341_, word_in[0]);
  not _17664_ (_09343_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _17665_ (_09344_, _09341_, _09343_);
  nor _17666_ (_09345_, _09344_, _09342_);
  nor _17667_ (_09346_, _09345_, _09340_);
  and _17668_ (_09347_, _09340_, word_in[8]);
  or _17669_ (_09348_, _09347_, _09346_);
  and _17670_ (_09349_, _09348_, _09339_);
  and _17671_ (_09350_, _09338_, _08544_);
  or _17672_ (_09351_, _09350_, _09349_);
  and _17673_ (_09352_, _09351_, _09337_);
  or _17674_ (_08120_, _09352_, _09336_);
  and _17675_ (_09353_, _09338_, _08694_);
  not _17676_ (_09354_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _17677_ (_09355_, _09341_, _09354_);
  and _17678_ (_09356_, _09341_, word_in[1]);
  nor _17679_ (_09357_, _09356_, _09355_);
  nor _17680_ (_09358_, _09357_, _09340_);
  and _17681_ (_09359_, _09340_, word_in[9]);
  or _17682_ (_09360_, _09359_, _09358_);
  and _17683_ (_09361_, _09360_, _09339_);
  or _17684_ (_09362_, _09361_, _09353_);
  and _17685_ (_09363_, _09362_, _09337_);
  and _17686_ (_09364_, _09335_, word_in[25]);
  or _17687_ (_08123_, _09364_, _09363_);
  and _17688_ (_09365_, _09338_, _08707_);
  not _17689_ (_09366_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _17690_ (_09367_, _09341_, _09366_);
  and _17691_ (_09368_, _09341_, word_in[2]);
  nor _17692_ (_09369_, _09368_, _09367_);
  nor _17693_ (_09370_, _09369_, _09340_);
  and _17694_ (_09371_, _09340_, word_in[10]);
  or _17695_ (_09372_, _09371_, _09370_);
  and _17696_ (_09373_, _09372_, _09339_);
  or _17697_ (_09374_, _09373_, _09365_);
  and _17698_ (_09375_, _09374_, _09337_);
  and _17699_ (_09376_, _09335_, word_in[26]);
  or _17700_ (_13490_, _09376_, _09375_);
  and _17701_ (_09377_, _09338_, _08712_);
  not _17702_ (_09378_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _17703_ (_09379_, _09341_, _09378_);
  and _17704_ (_09380_, _09341_, word_in[3]);
  nor _17705_ (_09381_, _09380_, _09379_);
  nor _17706_ (_09382_, _09381_, _09340_);
  and _17707_ (_09383_, _09340_, word_in[11]);
  or _17708_ (_09384_, _09383_, _09382_);
  and _17709_ (_09385_, _09384_, _09339_);
  or _17710_ (_09386_, _09385_, _09377_);
  and _17711_ (_09387_, _09386_, _09337_);
  and _17712_ (_09388_, _09335_, word_in[27]);
  or _17713_ (_13491_, _09388_, _09387_);
  and _17714_ (_09389_, _09338_, _08733_);
  not _17715_ (_09390_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _17716_ (_09391_, _09341_, _09390_);
  and _17717_ (_09392_, _09341_, word_in[4]);
  nor _17718_ (_09393_, _09392_, _09391_);
  nor _17719_ (_09394_, _09393_, _09340_);
  and _17720_ (_09395_, _09340_, word_in[12]);
  or _17721_ (_09396_, _09395_, _09394_);
  and _17722_ (_09397_, _09396_, _09339_);
  or _17723_ (_09398_, _09397_, _09389_);
  and _17724_ (_09399_, _09398_, _09337_);
  and _17725_ (_09400_, _09335_, word_in[28]);
  or _17726_ (_13492_, _09400_, _09399_);
  and _17727_ (_09401_, _09338_, _08746_);
  not _17728_ (_09402_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _17729_ (_09403_, _09341_, _09402_);
  and _17730_ (_09404_, _09341_, word_in[5]);
  nor _17731_ (_09405_, _09404_, _09403_);
  nor _17732_ (_09406_, _09405_, _09340_);
  and _17733_ (_09407_, _09340_, word_in[13]);
  or _17734_ (_09408_, _09407_, _09406_);
  and _17735_ (_09409_, _09408_, _09339_);
  or _17736_ (_09410_, _09409_, _09401_);
  and _17737_ (_09411_, _09410_, _09337_);
  and _17738_ (_09412_, _09335_, word_in[29]);
  or _17739_ (_13493_, _09412_, _09411_);
  not _17740_ (_09413_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _17741_ (_09414_, _09341_, _09413_);
  and _17742_ (_09415_, _09341_, word_in[6]);
  or _17743_ (_09416_, _09415_, _09414_);
  or _17744_ (_09417_, _09416_, _09340_);
  not _17745_ (_09418_, word_in[14]);
  nand _17746_ (_09419_, _09340_, _09418_);
  and _17747_ (_09420_, _09419_, _09417_);
  or _17748_ (_09421_, _09420_, _09338_);
  or _17749_ (_09422_, _09339_, _08759_);
  and _17750_ (_09423_, _09422_, _09337_);
  and _17751_ (_09424_, _09423_, _09421_);
  and _17752_ (_09425_, _09335_, word_in[30]);
  or _17753_ (_13494_, _09425_, _09424_);
  nor _17754_ (_09426_, _09341_, _07735_);
  and _17755_ (_09427_, _09341_, word_in[7]);
  or _17756_ (_09428_, _09427_, _09426_);
  or _17757_ (_09429_, _09428_, _09340_);
  nand _17758_ (_09430_, _09340_, _08642_);
  and _17759_ (_09431_, _09430_, _09429_);
  or _17760_ (_09432_, _09431_, _09338_);
  or _17761_ (_09433_, _09339_, _08037_);
  and _17762_ (_09434_, _09433_, _09432_);
  or _17763_ (_09435_, _09434_, _09335_);
  or _17764_ (_09436_, _09337_, word_in[31]);
  and _17765_ (_08141_, _09436_, _09435_);
  not _17766_ (_09437_, _08385_);
  not _17767_ (_09438_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _17768_ (_09439_, _08389_, _09438_);
  and _17769_ (_09440_, _08389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _17770_ (_09441_, _09440_, _09439_);
  and _17771_ (_09442_, _09441_, _09437_);
  nor _17772_ (_09443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor _17773_ (_09444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _17774_ (_09445_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _17775_ (_09446_, _09445_, _09444_);
  nor _17776_ (_09447_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _17777_ (_09448_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _17778_ (_09449_, _09448_, _09447_);
  and _17779_ (_09450_, _09449_, _09446_);
  and _17780_ (_09451_, _09450_, _09443_);
  and _17781_ (_09452_, _09451_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _17782_ (_09453_, _09452_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _17783_ (_09454_, _09453_, _08385_);
  nor _17784_ (_09455_, _09454_, _09442_);
  nor _17785_ (_09456_, _09455_, _08243_);
  nor _17786_ (_09457_, _06691_, _05604_);
  and _17787_ (_09458_, _09457_, _08243_);
  or _17788_ (_09459_, _09458_, _09456_);
  and _17789_ (_08210_, _09459_, _05141_);
  and _17790_ (_09460_, _08010_, _07949_);
  and _17791_ (_09461_, _09460_, _07788_);
  not _17792_ (_09462_, _09461_);
  and _17793_ (_09463_, _08016_, _08110_);
  and _17794_ (_09464_, _09463_, word_in[16]);
  not _17795_ (_09465_, _09463_);
  and _17796_ (_09466_, _08021_, _07779_);
  not _17797_ (_09467_, _09466_);
  not _17798_ (_09468_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _17799_ (_09469_, _07776_, _07626_);
  and _17800_ (_09470_, _08026_, _09469_);
  and _17801_ (_09471_, _09470_, _08531_);
  nor _17802_ (_09472_, _09471_, _09468_);
  and _17803_ (_09473_, _09471_, word_in[0]);
  or _17804_ (_09474_, _09473_, _09472_);
  and _17805_ (_09475_, _09474_, _09467_);
  and _17806_ (_09476_, _09466_, word_in[8]);
  or _17807_ (_09477_, _09476_, _09475_);
  and _17808_ (_09478_, _09477_, _09465_);
  or _17809_ (_09479_, _09478_, _09464_);
  and _17810_ (_09480_, _09479_, _09462_);
  and _17811_ (_09481_, _09461_, word_in[24]);
  or _17812_ (_13495_, _09481_, _09480_);
  and _17813_ (_09482_, _09463_, word_in[17]);
  not _17814_ (_09483_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _17815_ (_09484_, _09471_, _09483_);
  and _17816_ (_09485_, _09471_, word_in[1]);
  or _17817_ (_09486_, _09485_, _09484_);
  and _17818_ (_09487_, _09486_, _09467_);
  and _17819_ (_09488_, _09466_, word_in[9]);
  or _17820_ (_09489_, _09488_, _09487_);
  and _17821_ (_09490_, _09489_, _09465_);
  or _17822_ (_09491_, _09490_, _09482_);
  and _17823_ (_09492_, _09491_, _09462_);
  and _17824_ (_09493_, _09461_, word_in[25]);
  or _17825_ (_08219_, _09493_, _09492_);
  and _17826_ (_09494_, _09463_, word_in[18]);
  not _17827_ (_09495_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _17828_ (_09496_, _09471_, _09495_);
  and _17829_ (_09497_, _09471_, word_in[2]);
  or _17830_ (_09498_, _09497_, _09496_);
  and _17831_ (_09499_, _09498_, _09467_);
  and _17832_ (_09500_, _09466_, word_in[10]);
  or _17833_ (_09501_, _09500_, _09499_);
  and _17834_ (_09502_, _09501_, _09465_);
  or _17835_ (_09503_, _09502_, _09494_);
  and _17836_ (_09504_, _09503_, _09462_);
  and _17837_ (_09505_, _09461_, word_in[26]);
  or _17838_ (_08224_, _09505_, _09504_);
  and _17839_ (_09506_, _09463_, word_in[19]);
  not _17840_ (_09507_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _17841_ (_09508_, _09471_, _09507_);
  and _17842_ (_09509_, _09471_, word_in[3]);
  or _17843_ (_09510_, _09509_, _09508_);
  and _17844_ (_09511_, _09510_, _09467_);
  and _17845_ (_09512_, _09466_, word_in[11]);
  or _17846_ (_09513_, _09512_, _09511_);
  and _17847_ (_09514_, _09513_, _09465_);
  or _17848_ (_09515_, _09514_, _09506_);
  and _17849_ (_09516_, _09515_, _09462_);
  and _17850_ (_09517_, _09461_, word_in[27]);
  or _17851_ (_08229_, _09517_, _09516_);
  and _17852_ (_09518_, _09463_, word_in[20]);
  not _17853_ (_09519_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _17854_ (_09520_, _09471_, _09519_);
  and _17855_ (_09521_, _09471_, word_in[4]);
  or _17856_ (_09522_, _09521_, _09520_);
  and _17857_ (_09523_, _09522_, _09467_);
  and _17858_ (_09524_, _09466_, word_in[12]);
  or _17859_ (_09525_, _09524_, _09523_);
  and _17860_ (_09526_, _09525_, _09465_);
  or _17861_ (_09527_, _09526_, _09518_);
  and _17862_ (_09528_, _09527_, _09462_);
  and _17863_ (_09529_, _09461_, word_in[28]);
  or _17864_ (_08234_, _09529_, _09528_);
  and _17865_ (_09530_, _09463_, word_in[21]);
  not _17866_ (_09531_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _17867_ (_09532_, _09471_, _09531_);
  and _17868_ (_09533_, _09471_, word_in[5]);
  or _17869_ (_09534_, _09533_, _09532_);
  and _17870_ (_09535_, _09534_, _09467_);
  and _17871_ (_09536_, _09466_, word_in[13]);
  or _17872_ (_09537_, _09536_, _09535_);
  and _17873_ (_09538_, _09537_, _09465_);
  or _17874_ (_09539_, _09538_, _09530_);
  and _17875_ (_09540_, _09539_, _09462_);
  and _17876_ (_09541_, _09461_, word_in[29]);
  or _17877_ (_08236_, _09541_, _09540_);
  and _17878_ (_09542_, _09463_, word_in[22]);
  not _17879_ (_09543_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _17880_ (_09544_, _09471_, _09543_);
  and _17881_ (_09545_, _09471_, word_in[6]);
  or _17882_ (_09546_, _09545_, _09544_);
  and _17883_ (_09547_, _09546_, _09467_);
  and _17884_ (_09548_, _09466_, word_in[14]);
  or _17885_ (_09549_, _09548_, _09547_);
  and _17886_ (_09550_, _09549_, _09465_);
  or _17887_ (_09551_, _09550_, _09542_);
  and _17888_ (_09552_, _09551_, _09462_);
  and _17889_ (_09553_, _09461_, word_in[30]);
  or _17890_ (_08240_, _09553_, _09552_);
  and _17891_ (_09554_, _09463_, word_in[23]);
  nor _17892_ (_09555_, _09471_, _07827_);
  and _17893_ (_09556_, _09471_, word_in[7]);
  or _17894_ (_09557_, _09556_, _09555_);
  and _17895_ (_09558_, _09557_, _09467_);
  and _17896_ (_09559_, _09466_, word_in[15]);
  or _17897_ (_09560_, _09559_, _09558_);
  and _17898_ (_09561_, _09560_, _09465_);
  or _17899_ (_09562_, _09561_, _09554_);
  and _17900_ (_09563_, _09562_, _09462_);
  and _17901_ (_09565_, _09461_, word_in[31]);
  or _17902_ (_08244_, _09565_, _09563_);
  and _17903_ (_09566_, _08010_, _08110_);
  not _17904_ (_09567_, _09566_);
  and _17905_ (_09568_, _08661_, _07889_);
  and _17906_ (_09570_, _09568_, _08544_);
  not _17907_ (_09571_, _09568_);
  and _17908_ (_09573_, _08664_, _07783_);
  and _17909_ (_09574_, _09470_, _08668_);
  and _17910_ (_09575_, _09574_, _08666_);
  not _17911_ (_09576_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _17912_ (_09577_, _09574_, _09576_);
  nor _17913_ (_09578_, _09577_, _09575_);
  nor _17914_ (_09579_, _09578_, _09573_);
  and _17915_ (_09580_, _09573_, word_in[8]);
  or _17916_ (_09581_, _09580_, _09579_);
  and _17917_ (_09582_, _09581_, _09571_);
  or _17918_ (_09583_, _09582_, _09570_);
  and _17919_ (_09584_, _09583_, _09567_);
  and _17920_ (_09585_, _09566_, word_in[24]);
  or _17921_ (_08310_, _09585_, _09584_);
  and _17922_ (_09586_, _06695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _17923_ (_09587_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _17924_ (_09588_, _09587_, _06687_);
  and _17925_ (_09589_, _09588_, _06697_);
  or _17926_ (_09590_, _09589_, _09586_);
  and _17927_ (_08312_, _09590_, _05141_);
  and _17928_ (_09591_, _09574_, _08556_);
  not _17929_ (_09592_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _17930_ (_09593_, _09574_, _09592_);
  nor _17931_ (_09594_, _09593_, _09591_);
  nor _17932_ (_09595_, _09594_, _09573_);
  and _17933_ (_09596_, _09573_, word_in[9]);
  or _17934_ (_09597_, _09596_, _09595_);
  or _17935_ (_09598_, _09597_, _09568_);
  or _17936_ (_09599_, _09571_, _08694_);
  and _17937_ (_09600_, _09599_, _09567_);
  and _17938_ (_09601_, _09600_, _09598_);
  and _17939_ (_09602_, _09566_, word_in[25]);
  or _17940_ (_08314_, _09602_, _09601_);
  or _17941_ (_09603_, _09571_, _08707_);
  not _17942_ (_09604_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _17943_ (_09605_, _09574_, _09604_);
  and _17944_ (_09606_, _09574_, _08572_);
  or _17945_ (_09607_, _09606_, _09605_);
  or _17946_ (_09608_, _09607_, _09573_);
  not _17947_ (_09609_, _09573_);
  or _17948_ (_09610_, _09609_, word_in[10]);
  and _17949_ (_09611_, _09610_, _09608_);
  or _17950_ (_09612_, _09611_, _09568_);
  and _17951_ (_09613_, _09612_, _09603_);
  or _17952_ (_09614_, _09613_, _09566_);
  or _17953_ (_09615_, _09567_, word_in[26]);
  and _17954_ (_08317_, _09615_, _09614_);
  and _17955_ (_09616_, _09574_, _08586_);
  not _17956_ (_09617_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _17957_ (_09618_, _09574_, _09617_);
  nor _17958_ (_09619_, _09618_, _09616_);
  nor _17959_ (_09620_, _09619_, _09573_);
  and _17960_ (_09621_, _09573_, word_in[11]);
  or _17961_ (_09622_, _09621_, _09620_);
  and _17962_ (_09623_, _09622_, _09571_);
  and _17963_ (_09624_, _09568_, _08712_);
  or _17964_ (_09625_, _09624_, _09566_);
  or _17965_ (_09626_, _09625_, _09623_);
  or _17966_ (_09627_, _09567_, word_in[27]);
  and _17967_ (_08321_, _09627_, _09626_);
  not _17968_ (_09628_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _17969_ (_09629_, _09574_, _09628_);
  and _17970_ (_09630_, _09574_, _08598_);
  or _17971_ (_09631_, _09630_, _09629_);
  or _17972_ (_09632_, _09631_, _09573_);
  or _17973_ (_09633_, _09609_, word_in[12]);
  and _17974_ (_09634_, _09633_, _09632_);
  or _17975_ (_09635_, _09634_, _09568_);
  or _17976_ (_09636_, _09571_, _08733_);
  and _17977_ (_09637_, _09636_, _09567_);
  and _17978_ (_09638_, _09637_, _09635_);
  and _17979_ (_09639_, _09566_, word_in[28]);
  or _17980_ (_08325_, _09639_, _09638_);
  not _17981_ (_09640_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _17982_ (_09641_, _09574_, _09640_);
  and _17983_ (_09642_, _09574_, _08612_);
  or _17984_ (_09643_, _09642_, _09641_);
  or _17985_ (_09644_, _09643_, _09573_);
  or _17986_ (_09645_, _09609_, word_in[13]);
  and _17987_ (_09646_, _09645_, _09644_);
  or _17988_ (_09647_, _09646_, _09568_);
  or _17989_ (_09648_, _09571_, _08746_);
  and _17990_ (_09649_, _09648_, _09567_);
  and _17991_ (_09650_, _09649_, _09647_);
  and _17992_ (_09651_, _09566_, word_in[29]);
  or _17993_ (_08329_, _09651_, _09650_);
  not _17994_ (_09652_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _17995_ (_09653_, _09574_, _09652_);
  and _17996_ (_09654_, _09574_, _08628_);
  or _17997_ (_09655_, _09654_, _09653_);
  or _17998_ (_09656_, _09655_, _09573_);
  nand _17999_ (_09657_, _09573_, _09418_);
  and _18000_ (_09658_, _09657_, _09656_);
  or _18001_ (_09659_, _09658_, _09568_);
  or _18002_ (_09660_, _09571_, _08759_);
  and _18003_ (_09661_, _09660_, _09659_);
  or _18004_ (_09662_, _09661_, _09566_);
  or _18005_ (_09663_, _09567_, word_in[30]);
  and _18006_ (_08331_, _09663_, _09662_);
  or _18007_ (_09664_, _09571_, _08037_);
  nor _18008_ (_09665_, _09574_, _07722_);
  and _18009_ (_09666_, _09574_, _08029_);
  or _18010_ (_09667_, _09666_, _09665_);
  or _18011_ (_09668_, _09667_, _09573_);
  nand _18012_ (_09669_, _09573_, _08642_);
  and _18013_ (_09670_, _09669_, _09668_);
  or _18014_ (_09671_, _09670_, _09568_);
  and _18015_ (_09672_, _09671_, _09664_);
  or _18016_ (_09673_, _09672_, _09566_);
  or _18017_ (_09674_, _09567_, word_in[31]);
  and _18018_ (_08335_, _09674_, _09673_);
  and _18019_ (_09675_, _09460_, _07765_);
  and _18020_ (_09676_, _08778_, _07889_);
  not _18021_ (_09677_, _09676_);
  or _18022_ (_09678_, _09677_, _08544_);
  and _18023_ (_09679_, _08782_, _07783_);
  not _18024_ (_09680_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _18025_ (_09681_, _09470_, _08786_);
  nor _18026_ (_09682_, _09681_, _09680_);
  and _18027_ (_09683_, _09681_, _08666_);
  or _18028_ (_09684_, _09683_, _09682_);
  or _18029_ (_09685_, _09684_, _09679_);
  not _18030_ (_09686_, _09679_);
  or _18031_ (_09687_, _09686_, word_in[8]);
  and _18032_ (_09688_, _09687_, _09685_);
  or _18033_ (_09690_, _09688_, _09676_);
  and _18034_ (_09691_, _09690_, _09678_);
  or _18035_ (_09692_, _09691_, _09675_);
  not _18036_ (_09693_, _09675_);
  or _18037_ (_09694_, _09693_, word_in[24]);
  and _18038_ (_08400_, _09694_, _09692_);
  not _18039_ (_09695_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _18040_ (_09696_, _09681_, _09695_);
  and _18041_ (_09697_, _09681_, _08556_);
  or _18042_ (_09698_, _09697_, _09696_);
  or _18043_ (_09699_, _09698_, _09679_);
  or _18044_ (_09700_, _09686_, word_in[9]);
  and _18045_ (_09701_, _09700_, _09699_);
  or _18046_ (_09702_, _09701_, _09676_);
  or _18047_ (_09703_, _09677_, _08694_);
  and _18048_ (_09704_, _09703_, _09693_);
  and _18049_ (_09705_, _09704_, _09702_);
  and _18050_ (_09706_, _09675_, word_in[25]);
  or _18051_ (_08403_, _09706_, _09705_);
  or _18052_ (_09707_, _09677_, _08707_);
  not _18053_ (_09708_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _18054_ (_09709_, _09681_, _09708_);
  and _18055_ (_09710_, _09681_, _08572_);
  or _18056_ (_09711_, _09710_, _09709_);
  or _18057_ (_09712_, _09711_, _09679_);
  or _18058_ (_09713_, _09686_, word_in[10]);
  and _18059_ (_09714_, _09713_, _09712_);
  or _18060_ (_09715_, _09714_, _09676_);
  and _18061_ (_09716_, _09715_, _09707_);
  or _18062_ (_09717_, _09716_, _09675_);
  or _18063_ (_09718_, _09693_, word_in[26]);
  and _18064_ (_08407_, _09718_, _09717_);
  or _18065_ (_09719_, _09677_, _08712_);
  not _18066_ (_09720_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _18067_ (_09721_, _09681_, _09720_);
  and _18068_ (_09722_, _09681_, _08586_);
  or _18069_ (_09723_, _09722_, _09721_);
  or _18070_ (_09724_, _09723_, _09679_);
  or _18071_ (_09725_, _09686_, word_in[11]);
  and _18072_ (_09726_, _09725_, _09724_);
  or _18073_ (_09727_, _09726_, _09676_);
  and _18074_ (_09728_, _09727_, _09719_);
  or _18075_ (_09729_, _09728_, _09675_);
  or _18076_ (_09730_, _09693_, word_in[27]);
  and _18077_ (_08410_, _09730_, _09729_);
  not _18078_ (_09731_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _18079_ (_09732_, _09681_, _09731_);
  and _18080_ (_09733_, _09681_, _08598_);
  or _18081_ (_09734_, _09733_, _09732_);
  or _18082_ (_09735_, _09734_, _09679_);
  or _18083_ (_09736_, _09686_, word_in[12]);
  and _18084_ (_09737_, _09736_, _09735_);
  or _18085_ (_09738_, _09737_, _09676_);
  or _18086_ (_09739_, _09677_, _08733_);
  and _18087_ (_09740_, _09739_, _09693_);
  and _18088_ (_09741_, _09740_, _09738_);
  and _18089_ (_09742_, _09675_, word_in[28]);
  or _18090_ (_08413_, _09742_, _09741_);
  or _18091_ (_09743_, _09677_, _08746_);
  not _18092_ (_09744_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _18093_ (_09745_, _09681_, _09744_);
  and _18094_ (_09746_, _09681_, _08612_);
  or _18095_ (_09747_, _09746_, _09745_);
  or _18096_ (_09748_, _09747_, _09679_);
  or _18097_ (_09749_, _09686_, word_in[13]);
  and _18098_ (_09750_, _09749_, _09748_);
  or _18099_ (_09751_, _09750_, _09676_);
  and _18100_ (_09752_, _09751_, _09743_);
  or _18101_ (_09753_, _09752_, _09675_);
  or _18102_ (_09754_, _09693_, word_in[29]);
  and _18103_ (_08416_, _09754_, _09753_);
  or _18104_ (_09755_, _09677_, _08759_);
  not _18105_ (_09756_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _18106_ (_09757_, _09681_, _09756_);
  and _18107_ (_09758_, _09681_, _08628_);
  or _18108_ (_09759_, _09758_, _09757_);
  or _18109_ (_09760_, _09759_, _09679_);
  nand _18110_ (_09761_, _09679_, _09418_);
  and _18111_ (_09762_, _09761_, _09760_);
  or _18112_ (_09763_, _09762_, _09676_);
  and _18113_ (_09764_, _09763_, _09755_);
  and _18114_ (_09765_, _09764_, _09693_);
  and _18115_ (_09766_, _09675_, word_in[30]);
  or _18116_ (_08419_, _09766_, _09765_);
  nor _18117_ (_09767_, _09681_, _07822_);
  and _18118_ (_09768_, _09681_, _08029_);
  or _18119_ (_09769_, _09768_, _09767_);
  or _18120_ (_09770_, _09769_, _09679_);
  nand _18121_ (_09771_, _09679_, _08642_);
  and _18122_ (_09772_, _09771_, _09770_);
  or _18123_ (_09773_, _09772_, _09676_);
  or _18124_ (_09774_, _09677_, _08037_);
  and _18125_ (_09775_, _09774_, _09693_);
  and _18126_ (_09776_, _09775_, _09773_);
  and _18127_ (_09777_, _09675_, word_in[31]);
  or _18128_ (_08421_, _09777_, _09776_);
  and _18129_ (_09778_, _06703_, _05277_);
  not _18130_ (_09779_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _18131_ (_09780_, _05277_, _09779_);
  or _18132_ (_09781_, _09780_, _05572_);
  or _18133_ (_09782_, _09781_, _09778_);
  or _18134_ (_09783_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _18135_ (_09784_, _09783_, _05141_);
  and _18136_ (_08473_, _09784_, _09782_);
  not _18137_ (_09785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  or _18138_ (_09786_, _06695_, _09785_);
  or _18139_ (_09787_, _06697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _18140_ (_09788_, _09787_, _05141_);
  and _18141_ (_08477_, _09788_, _09786_);
  and _18142_ (_09789_, _08917_, _07889_);
  and _18143_ (_09790_, _08022_, _07783_);
  and _18144_ (_09791_, _09790_, word_in[8]);
  and _18145_ (_09792_, _09470_, _08025_);
  and _18146_ (_09793_, _09792_, _08666_);
  not _18147_ (_09794_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor _18148_ (_09795_, _09792_, _09794_);
  nor _18149_ (_09796_, _09795_, _09793_);
  nor _18150_ (_09797_, _09796_, _09790_);
  or _18151_ (_09798_, _09797_, _09791_);
  or _18152_ (_09799_, _09798_, _09789_);
  and _18153_ (_09800_, _09460_, _07761_);
  not _18154_ (_09801_, _09789_);
  nor _18155_ (_09802_, _09801_, _08544_);
  nor _18156_ (_09803_, _09802_, _09800_);
  and _18157_ (_09804_, _09803_, _09799_);
  and _18158_ (_09805_, _09800_, word_in[24]);
  or _18159_ (_08486_, _09805_, _09804_);
  not _18160_ (_09806_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _18161_ (_09807_, _09792_, _09806_);
  and _18162_ (_09808_, _09792_, _08556_);
  or _18163_ (_09809_, _09808_, _09807_);
  or _18164_ (_09810_, _09809_, _09790_);
  not _18165_ (_09811_, _09790_);
  or _18166_ (_09812_, _09811_, word_in[9]);
  and _18167_ (_09813_, _09812_, _09810_);
  or _18168_ (_09814_, _09813_, _09789_);
  not _18169_ (_09815_, _09800_);
  or _18170_ (_09816_, _09801_, _08694_);
  and _18171_ (_09817_, _09816_, _09815_);
  and _18172_ (_09818_, _09817_, _09814_);
  and _18173_ (_09819_, _09800_, _08566_);
  or _18174_ (_08490_, _09819_, _09818_);
  not _18175_ (_09820_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _18176_ (_09821_, _09792_, _09820_);
  and _18177_ (_09822_, _09792_, _08572_);
  or _18178_ (_09823_, _09822_, _09821_);
  or _18179_ (_09824_, _09823_, _09790_);
  or _18180_ (_09825_, _09811_, word_in[10]);
  and _18181_ (_09826_, _09825_, _09824_);
  or _18182_ (_09827_, _09826_, _09789_);
  or _18183_ (_09828_, _09801_, _08707_);
  and _18184_ (_09829_, _09828_, _09815_);
  and _18185_ (_09830_, _09829_, _09827_);
  and _18186_ (_09831_, _09800_, _08568_);
  or _18187_ (_08493_, _09831_, _09830_);
  not _18188_ (_09832_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _18189_ (_09834_, _09792_, _09832_);
  and _18190_ (_09835_, _09792_, _08586_);
  or _18191_ (_09836_, _09835_, _09834_);
  or _18192_ (_09837_, _09836_, _09790_);
  or _18193_ (_09838_, _09811_, word_in[11]);
  and _18194_ (_09839_, _09838_, _09837_);
  or _18195_ (_09840_, _09839_, _09789_);
  or _18196_ (_09841_, _09801_, _08712_);
  and _18197_ (_09842_, _09841_, _09815_);
  and _18198_ (_09843_, _09842_, _09840_);
  and _18199_ (_09844_, _09800_, _08582_);
  or _18200_ (_08495_, _09844_, _09843_);
  not _18201_ (_09845_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _18202_ (_09846_, _09792_, _09845_);
  and _18203_ (_09847_, _09792_, _08598_);
  or _18204_ (_09848_, _09847_, _09846_);
  or _18205_ (_09849_, _09848_, _09790_);
  or _18206_ (_09850_, _09811_, word_in[12]);
  and _18207_ (_09851_, _09850_, _09849_);
  or _18208_ (_09852_, _09851_, _09789_);
  or _18209_ (_09853_, _09801_, _08733_);
  and _18210_ (_09854_, _09853_, _09815_);
  and _18211_ (_09856_, _09854_, _09852_);
  and _18212_ (_09857_, _09800_, _08608_);
  or _18213_ (_08498_, _09857_, _09856_);
  not _18214_ (_09858_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _18215_ (_09860_, _09792_, _09858_);
  and _18216_ (_09861_, _09792_, _08612_);
  or _18217_ (_09863_, _09861_, _09860_);
  or _18218_ (_09864_, _09863_, _09790_);
  or _18219_ (_09865_, _09811_, word_in[13]);
  and _18220_ (_09866_, _09865_, _09864_);
  or _18221_ (_09867_, _09866_, _09789_);
  or _18222_ (_09868_, _09801_, _08746_);
  and _18223_ (_09869_, _09868_, _09815_);
  and _18224_ (_09870_, _09869_, _09867_);
  and _18225_ (_09871_, _09800_, _08622_);
  or _18226_ (_08502_, _09871_, _09870_);
  not _18227_ (_09872_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _18228_ (_09873_, _09792_, _09872_);
  and _18229_ (_09874_, _09792_, _08628_);
  or _18230_ (_09875_, _09874_, _09873_);
  or _18231_ (_09876_, _09875_, _09790_);
  nand _18232_ (_09877_, _09790_, _09418_);
  and _18233_ (_09878_, _09877_, _09876_);
  or _18234_ (_09879_, _09878_, _09789_);
  or _18235_ (_09880_, _09801_, _08759_);
  and _18236_ (_09881_, _09880_, _09815_);
  and _18237_ (_09882_, _09881_, _09879_);
  and _18238_ (_09883_, _09800_, _08624_);
  or _18239_ (_08506_, _09883_, _09882_);
  nor _18240_ (_09884_, _09792_, _07711_);
  and _18241_ (_09885_, _09792_, _08029_);
  or _18242_ (_09886_, _09885_, _09884_);
  or _18243_ (_09887_, _09886_, _09790_);
  nand _18244_ (_09888_, _09790_, _08642_);
  and _18245_ (_09889_, _09888_, _09887_);
  or _18246_ (_09890_, _09889_, _09789_);
  or _18247_ (_09891_, _09801_, _08037_);
  and _18248_ (_09892_, _09891_, _09815_);
  and _18249_ (_09893_, _09892_, _09890_);
  and _18250_ (_09894_, _09800_, _08011_);
  or _18251_ (_08510_, _09894_, _09893_);
  and _18252_ (_09895_, _08382_, _05522_);
  and _18253_ (_09896_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _18254_ (_09897_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _18255_ (_09898_, _09897_, _09896_);
  nor _18256_ (_09899_, _09898_, _08243_);
  and _18257_ (_09900_, _08396_, _06290_);
  or _18258_ (_09901_, _09900_, _09899_);
  or _18259_ (_09902_, _09901_, _09895_);
  and _18260_ (_08517_, _09902_, _05141_);
  and _18261_ (_09903_, _08018_, _07798_);
  not _18262_ (_09904_, _09903_);
  and _18263_ (_09905_, _08021_, _08254_);
  not _18264_ (_09906_, _09905_);
  or _18265_ (_09907_, _09906_, word_in[8]);
  not _18266_ (_09908_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _18267_ (_09909_, _08531_, _08027_);
  nor _18268_ (_09910_, _09909_, _09908_);
  and _18269_ (_09911_, _09909_, word_in[0]);
  or _18270_ (_09912_, _09911_, _09910_);
  or _18271_ (_09913_, _09912_, _09905_);
  and _18272_ (_09914_, _09913_, _09907_);
  and _18273_ (_09915_, _09914_, _09904_);
  not _18274_ (_09916_, _07946_);
  and _18275_ (_09917_, _09034_, _09916_);
  and _18276_ (_09918_, _09917_, _07788_);
  and _18277_ (_09919_, _09903_, _08544_);
  or _18278_ (_09920_, _09919_, _09918_);
  or _18279_ (_09921_, _09920_, _09915_);
  not _18280_ (_09922_, _09918_);
  or _18281_ (_09923_, _09922_, _09040_);
  and _18282_ (_13475_, _09923_, _09921_);
  not _18283_ (_09924_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _18284_ (_09925_, _09909_, _09924_);
  and _18285_ (_09926_, _09909_, word_in[1]);
  or _18286_ (_09927_, _09926_, _09925_);
  and _18287_ (_09928_, _09927_, _09906_);
  and _18288_ (_09929_, _09905_, word_in[9]);
  or _18289_ (_09930_, _09929_, _09928_);
  and _18290_ (_09931_, _09930_, _09904_);
  and _18291_ (_09932_, _09903_, _08694_);
  or _18292_ (_09933_, _09932_, _09918_);
  or _18293_ (_09934_, _09933_, _09931_);
  or _18294_ (_09935_, _09922_, _08566_);
  and _18295_ (_13476_, _09935_, _09934_);
  not _18296_ (_09936_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _18297_ (_09937_, _09909_, _09936_);
  and _18298_ (_09938_, _09909_, word_in[2]);
  or _18299_ (_09939_, _09938_, _09937_);
  and _18300_ (_09940_, _09939_, _09906_);
  and _18301_ (_09941_, _09905_, word_in[10]);
  or _18302_ (_09942_, _09941_, _09940_);
  and _18303_ (_09943_, _09942_, _09904_);
  and _18304_ (_09944_, _09903_, _08707_);
  or _18305_ (_09945_, _09944_, _09918_);
  or _18306_ (_09946_, _09945_, _09943_);
  or _18307_ (_09947_, _09922_, _08568_);
  and _18308_ (_13477_, _09947_, _09946_);
  not _18309_ (_09948_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _18310_ (_09949_, _09909_, _09948_);
  and _18311_ (_09950_, _09909_, word_in[3]);
  or _18312_ (_09951_, _09950_, _09949_);
  and _18313_ (_09952_, _09951_, _09906_);
  and _18314_ (_09953_, _09905_, word_in[11]);
  or _18315_ (_09954_, _09953_, _09952_);
  and _18316_ (_09955_, _09954_, _09904_);
  and _18317_ (_09956_, _09903_, _08712_);
  or _18318_ (_09957_, _09956_, _09918_);
  or _18319_ (_09958_, _09957_, _09955_);
  or _18320_ (_09959_, _09922_, _08582_);
  and _18321_ (_13478_, _09959_, _09958_);
  not _18322_ (_09960_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _18323_ (_09961_, _09909_, _09960_);
  and _18324_ (_09962_, _09909_, word_in[4]);
  or _18325_ (_09963_, _09962_, _09961_);
  and _18326_ (_09964_, _09963_, _09906_);
  and _18327_ (_09965_, _09905_, word_in[12]);
  or _18328_ (_09966_, _09965_, _09964_);
  and _18329_ (_09967_, _09966_, _09904_);
  and _18330_ (_09968_, _09903_, _08733_);
  or _18331_ (_09969_, _09968_, _09918_);
  or _18332_ (_09970_, _09969_, _09967_);
  or _18333_ (_09971_, _09922_, _08608_);
  and _18334_ (_13479_, _09971_, _09970_);
  not _18335_ (_09972_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _18336_ (_09973_, _09909_, _09972_);
  and _18337_ (_09974_, _09909_, word_in[5]);
  or _18338_ (_09975_, _09974_, _09973_);
  or _18339_ (_09976_, _09975_, _09905_);
  or _18340_ (_09977_, _09906_, word_in[13]);
  and _18341_ (_09978_, _09977_, _09976_);
  and _18342_ (_09979_, _09978_, _09904_);
  and _18343_ (_09980_, _09903_, _08746_);
  or _18344_ (_09981_, _09980_, _09918_);
  or _18345_ (_09982_, _09981_, _09979_);
  or _18346_ (_09983_, _09922_, _08622_);
  and _18347_ (_13480_, _09983_, _09982_);
  not _18348_ (_09984_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _18349_ (_09985_, _09909_, _09984_);
  and _18350_ (_09986_, _09909_, word_in[6]);
  or _18351_ (_09987_, _09986_, _09985_);
  and _18352_ (_09988_, _09987_, _09906_);
  and _18353_ (_09989_, _09905_, word_in[14]);
  or _18354_ (_09990_, _09989_, _09988_);
  and _18355_ (_09991_, _09990_, _09904_);
  and _18356_ (_09992_, _09903_, _08759_);
  or _18357_ (_09993_, _09992_, _09918_);
  or _18358_ (_09994_, _09993_, _09991_);
  or _18359_ (_09995_, _09922_, _08624_);
  and _18360_ (_13481_, _09995_, _09994_);
  nor _18361_ (_09996_, _09909_, _07864_);
  and _18362_ (_09997_, _09909_, word_in[7]);
  or _18363_ (_09998_, _09997_, _09996_);
  and _18364_ (_09999_, _09998_, _09906_);
  and _18365_ (_10000_, _09905_, word_in[15]);
  or _18366_ (_10001_, _10000_, _09999_);
  and _18367_ (_10002_, _10001_, _09904_);
  and _18368_ (_10003_, _09903_, _08037_);
  or _18369_ (_10004_, _10003_, _09918_);
  or _18370_ (_10005_, _10004_, _10002_);
  or _18371_ (_10006_, _09922_, _08011_);
  and _18372_ (_13482_, _10006_, _10005_);
  and _18373_ (_10007_, _09917_, _07798_);
  and _18374_ (_10008_, _08018_, _07765_);
  and _18375_ (_10009_, _08664_, _07811_);
  not _18376_ (_10010_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _18377_ (_10011_, _08668_, _08027_);
  nor _18378_ (_10012_, _10011_, _10010_);
  and _18379_ (_10013_, _10011_, _08666_);
  or _18380_ (_10014_, _10013_, _10012_);
  or _18381_ (_10015_, _10014_, _10009_);
  not _18382_ (_10016_, word_in[8]);
  nand _18383_ (_10017_, _10009_, _10016_);
  and _18384_ (_10018_, _10017_, _10015_);
  or _18385_ (_10019_, _10018_, _10008_);
  not _18386_ (_10020_, _10008_);
  or _18387_ (_10021_, _10020_, _08544_);
  and _18388_ (_10022_, _10021_, _10019_);
  or _18389_ (_10023_, _10022_, _10007_);
  not _18390_ (_10024_, _10007_);
  or _18391_ (_10025_, _10024_, word_in[24]);
  and _18392_ (_13483_, _10025_, _10023_);
  not _18393_ (_10026_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _18394_ (_10027_, _10011_, _10026_);
  and _18395_ (_10028_, _10011_, _08556_);
  nor _18396_ (_10029_, _10028_, _10027_);
  nor _18397_ (_10030_, _10029_, _10009_);
  and _18398_ (_10031_, _10009_, word_in[9]);
  or _18399_ (_10032_, _10031_, _10030_);
  and _18400_ (_10033_, _10032_, _10020_);
  and _18401_ (_10034_, _10008_, _08694_);
  or _18402_ (_10035_, _10034_, _10007_);
  or _18403_ (_10036_, _10035_, _10033_);
  or _18404_ (_10037_, _10024_, word_in[25]);
  and _18405_ (_13484_, _10037_, _10036_);
  not _18406_ (_10038_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _18407_ (_10039_, _10011_, _10038_);
  and _18408_ (_10040_, _10011_, _08572_);
  nor _18409_ (_10041_, _10040_, _10039_);
  nor _18410_ (_10042_, _10041_, _10009_);
  and _18411_ (_10043_, _10009_, word_in[10]);
  or _18412_ (_10044_, _10043_, _10042_);
  and _18413_ (_10045_, _10044_, _10020_);
  and _18414_ (_10046_, _10008_, _08707_);
  or _18415_ (_10047_, _10046_, _10007_);
  or _18416_ (_10048_, _10047_, _10045_);
  or _18417_ (_10049_, _10024_, word_in[26]);
  and _18418_ (_13485_, _10049_, _10048_);
  not _18419_ (_10050_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _18420_ (_10051_, _10011_, _10050_);
  and _18421_ (_10052_, _10011_, _08586_);
  nor _18422_ (_10053_, _10052_, _10051_);
  nor _18423_ (_10054_, _10053_, _10009_);
  and _18424_ (_10055_, _10009_, word_in[11]);
  or _18425_ (_10056_, _10055_, _10054_);
  and _18426_ (_10057_, _10056_, _10020_);
  and _18427_ (_10058_, _10008_, _08712_);
  or _18428_ (_10059_, _10058_, _10007_);
  or _18429_ (_10060_, _10059_, _10057_);
  or _18430_ (_10061_, _10024_, word_in[27]);
  and _18431_ (_08679_, _10061_, _10060_);
  and _18432_ (_10062_, _08382_, _06290_);
  and _18433_ (_10063_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _18434_ (_10064_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _18435_ (_10065_, _10064_, _10063_);
  nor _18436_ (_10066_, _10065_, _08243_);
  and _18437_ (_10067_, _08396_, _05561_);
  or _18438_ (_10069_, _10067_, _10066_);
  or _18439_ (_10070_, _10069_, _10062_);
  and _18440_ (_08682_, _10070_, _05141_);
  not _18441_ (_10071_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _18442_ (_10073_, _10011_, _10071_);
  and _18443_ (_10074_, _10011_, _08598_);
  nor _18444_ (_10075_, _10074_, _10073_);
  nor _18445_ (_10076_, _10075_, _10009_);
  and _18446_ (_10077_, _10009_, word_in[12]);
  or _18447_ (_10078_, _10077_, _10076_);
  and _18448_ (_10079_, _10078_, _10020_);
  and _18449_ (_10080_, _10008_, _08733_);
  or _18450_ (_10081_, _10080_, _10007_);
  or _18451_ (_10082_, _10081_, _10079_);
  or _18452_ (_10083_, _10024_, word_in[28]);
  and _18453_ (_13486_, _10083_, _10082_);
  not _18454_ (_10084_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _18455_ (_10085_, _10011_, _10084_);
  and _18456_ (_10086_, _10011_, _08612_);
  nor _18457_ (_10087_, _10086_, _10085_);
  nor _18458_ (_10088_, _10087_, _10009_);
  and _18459_ (_10089_, _10009_, word_in[13]);
  or _18460_ (_10090_, _10089_, _10088_);
  and _18461_ (_10091_, _10090_, _10020_);
  and _18462_ (_10092_, _10008_, _08746_);
  or _18463_ (_10093_, _10092_, _10007_);
  or _18464_ (_10094_, _10093_, _10091_);
  or _18465_ (_10095_, _10024_, word_in[29]);
  and _18466_ (_13487_, _10095_, _10094_);
  not _18467_ (_10096_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _18468_ (_10097_, _10011_, _10096_);
  and _18469_ (_10098_, _10011_, _08628_);
  nor _18470_ (_10099_, _10098_, _10097_);
  nor _18471_ (_10100_, _10099_, _10009_);
  and _18472_ (_10101_, _10009_, word_in[14]);
  or _18473_ (_10102_, _10101_, _10100_);
  and _18474_ (_10103_, _10102_, _10020_);
  and _18475_ (_10104_, _10008_, _08759_);
  or _18476_ (_10105_, _10104_, _10007_);
  or _18477_ (_10106_, _10105_, _10103_);
  or _18478_ (_10107_, _10024_, word_in[30]);
  and _18479_ (_13488_, _10107_, _10106_);
  and _18480_ (_10108_, _08382_, _06283_);
  and _18481_ (_10109_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _18482_ (_10110_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _18483_ (_10111_, _10110_, _10109_);
  nor _18484_ (_10112_, _10111_, _08243_);
  and _18485_ (_10113_, _08396_, _06004_);
  or _18486_ (_10114_, _10113_, _10112_);
  or _18487_ (_10116_, _10114_, _10108_);
  and _18488_ (_08691_, _10116_, _05141_);
  nor _18489_ (_10117_, _10011_, _07717_);
  and _18490_ (_10118_, _10011_, _08029_);
  nor _18491_ (_10119_, _10118_, _10117_);
  nor _18492_ (_10120_, _10119_, _10009_);
  and _18493_ (_10121_, _10009_, word_in[15]);
  or _18494_ (_10122_, _10121_, _10120_);
  and _18495_ (_10123_, _10122_, _10020_);
  and _18496_ (_10124_, _10008_, _08037_);
  or _18497_ (_10125_, _10124_, _10007_);
  or _18498_ (_10126_, _10125_, _10123_);
  or _18499_ (_10127_, _10024_, word_in[31]);
  and _18500_ (_13489_, _10127_, _10126_);
  and _18501_ (_10128_, _09917_, _07765_);
  and _18502_ (_10129_, _08018_, _07761_);
  and _18503_ (_10130_, _08782_, _07811_);
  not _18504_ (_10131_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _18505_ (_10132_, _08786_, _08008_);
  nor _18506_ (_10133_, _10132_, _10131_);
  and _18507_ (_10134_, _10132_, _08666_);
  or _18508_ (_10135_, _10134_, _10133_);
  or _18509_ (_10136_, _10135_, _10130_);
  nand _18510_ (_10137_, _10130_, _10016_);
  and _18511_ (_10138_, _10137_, _10136_);
  or _18512_ (_10139_, _10138_, _10129_);
  not _18513_ (_10140_, _10129_);
  or _18514_ (_10141_, _10140_, _08544_);
  and _18515_ (_10142_, _10141_, _10139_);
  or _18516_ (_10143_, _10142_, _10128_);
  not _18517_ (_10144_, _10128_);
  or _18518_ (_10145_, _10144_, word_in[24]);
  and _18519_ (_08770_, _10145_, _10143_);
  not _18520_ (_10146_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _18521_ (_10147_, _10132_, _10146_);
  and _18522_ (_10148_, _10132_, _08556_);
  nor _18523_ (_10149_, _10148_, _10147_);
  nor _18524_ (_10150_, _10149_, _10130_);
  and _18525_ (_10151_, _10130_, word_in[9]);
  or _18526_ (_10152_, _10151_, _10150_);
  and _18527_ (_10154_, _10152_, _10140_);
  and _18528_ (_10155_, _10129_, _08694_);
  or _18529_ (_10156_, _10155_, _10128_);
  or _18530_ (_10157_, _10156_, _10154_);
  or _18531_ (_10158_, _10144_, word_in[25]);
  and _18532_ (_08775_, _10158_, _10157_);
  not _18533_ (_10159_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _18534_ (_10160_, _10132_, _10159_);
  and _18535_ (_10161_, _10132_, _08572_);
  or _18536_ (_10162_, _10161_, _10160_);
  or _18537_ (_10163_, _10162_, _10130_);
  not _18538_ (_10164_, _10130_);
  or _18539_ (_10165_, _10164_, word_in[10]);
  and _18540_ (_10166_, _10165_, _10163_);
  or _18541_ (_10167_, _10166_, _10129_);
  or _18542_ (_10168_, _10140_, _08707_);
  and _18543_ (_10169_, _10168_, _10144_);
  and _18544_ (_10170_, _10169_, _10167_);
  and _18545_ (_10171_, _10128_, word_in[26]);
  or _18546_ (_08777_, _10171_, _10170_);
  not _18547_ (_10172_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _18548_ (_10173_, _10132_, _10172_);
  and _18549_ (_10174_, _10132_, _08586_);
  nor _18550_ (_10175_, _10174_, _10173_);
  nor _18551_ (_10176_, _10175_, _10130_);
  and _18552_ (_10177_, _10130_, word_in[11]);
  or _18553_ (_10178_, _10177_, _10176_);
  and _18554_ (_10179_, _10178_, _10140_);
  and _18555_ (_10180_, _10129_, _08712_);
  or _18556_ (_10181_, _10180_, _10128_);
  or _18557_ (_10182_, _10181_, _10179_);
  or _18558_ (_10183_, _10144_, word_in[27]);
  and _18559_ (_08781_, _10183_, _10182_);
  not _18560_ (_10184_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _18561_ (_10185_, _10132_, _10184_);
  and _18562_ (_10186_, _10132_, _08598_);
  nor _18563_ (_10187_, _10186_, _10185_);
  nor _18564_ (_10188_, _10187_, _10130_);
  and _18565_ (_10189_, _10130_, word_in[12]);
  or _18566_ (_10190_, _10189_, _10188_);
  and _18567_ (_10192_, _10190_, _10140_);
  and _18568_ (_10193_, _10129_, _08733_);
  or _18569_ (_10194_, _10193_, _10128_);
  or _18570_ (_10195_, _10194_, _10192_);
  or _18571_ (_10196_, _10144_, word_in[28]);
  and _18572_ (_08785_, _10196_, _10195_);
  not _18573_ (_10197_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _18574_ (_10198_, _10132_, _10197_);
  and _18575_ (_10199_, _10132_, _08612_);
  nor _18576_ (_10200_, _10199_, _10198_);
  nor _18577_ (_10201_, _10200_, _10130_);
  and _18578_ (_10202_, _10130_, word_in[13]);
  or _18579_ (_10203_, _10202_, _10201_);
  and _18580_ (_10204_, _10203_, _10140_);
  and _18581_ (_10205_, _10129_, _08746_);
  or _18582_ (_10206_, _10205_, _10128_);
  or _18583_ (_10207_, _10206_, _10204_);
  or _18584_ (_10208_, _10144_, word_in[29]);
  and _18585_ (_08788_, _10208_, _10207_);
  not _18586_ (_10209_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _18587_ (_10210_, _10132_, _10209_);
  and _18588_ (_10211_, _10132_, _08628_);
  nor _18589_ (_10212_, _10211_, _10210_);
  nor _18590_ (_10213_, _10212_, _10130_);
  and _18591_ (_10214_, _10130_, word_in[14]);
  or _18592_ (_10215_, _10214_, _10213_);
  and _18593_ (_10216_, _10215_, _10140_);
  and _18594_ (_10217_, _10129_, _08759_);
  or _18595_ (_10218_, _10217_, _10128_);
  or _18596_ (_10219_, _10218_, _10216_);
  or _18597_ (_10220_, _10144_, word_in[30]);
  and _18598_ (_08792_, _10220_, _10219_);
  nor _18599_ (_10221_, _10132_, _07858_);
  and _18600_ (_10222_, _10132_, _08029_);
  nor _18601_ (_10223_, _10222_, _10221_);
  nor _18602_ (_10224_, _10223_, _10130_);
  and _18603_ (_10225_, _10130_, word_in[15]);
  or _18604_ (_10226_, _10225_, _10224_);
  and _18605_ (_10227_, _10226_, _10140_);
  and _18606_ (_10228_, _10129_, _08037_);
  or _18607_ (_10229_, _10228_, _10128_);
  or _18608_ (_10230_, _10229_, _10227_);
  or _18609_ (_10231_, _10144_, word_in[31]);
  and _18610_ (_08796_, _10231_, _10230_);
  and _18611_ (_10232_, _09040_, _08013_);
  and _18612_ (_10233_, _08028_, word_in[0]);
  not _18613_ (_10234_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _18614_ (_10235_, _08028_, _10234_);
  nor _18615_ (_10237_, _10235_, _10233_);
  nor _18616_ (_10238_, _10237_, _08023_);
  and _18617_ (_10240_, _08023_, word_in[8]);
  or _18618_ (_10241_, _10240_, _10238_);
  and _18619_ (_10242_, _10241_, _08020_);
  and _18620_ (_10243_, _08544_, _08019_);
  or _18621_ (_10244_, _10243_, _10242_);
  and _18622_ (_10246_, _10244_, _08015_);
  or _18623_ (_08867_, _10246_, _10232_);
  and _18624_ (_10247_, _08566_, _08013_);
  not _18625_ (_10248_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _18626_ (_10249_, _08028_, _10248_);
  and _18627_ (_10250_, _08028_, word_in[1]);
  nor _18628_ (_10252_, _10250_, _10249_);
  nor _18629_ (_10253_, _10252_, _08023_);
  and _18630_ (_10254_, _08023_, word_in[9]);
  or _18631_ (_10255_, _10254_, _10253_);
  and _18632_ (_10256_, _10255_, _08020_);
  and _18633_ (_10257_, _08694_, _08019_);
  or _18634_ (_10258_, _10257_, _10256_);
  and _18635_ (_10259_, _10258_, _08015_);
  or _18636_ (_08870_, _10259_, _10247_);
  not _18637_ (_10260_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _18638_ (_10261_, _08028_, _10260_);
  and _18639_ (_10262_, _08028_, word_in[2]);
  nor _18640_ (_10263_, _10262_, _10261_);
  nor _18641_ (_10264_, _10263_, _08023_);
  and _18642_ (_10265_, _08023_, word_in[10]);
  or _18643_ (_10266_, _10265_, _10264_);
  and _18644_ (_10267_, _10266_, _08020_);
  and _18645_ (_10268_, _08707_, _08019_);
  or _18646_ (_10269_, _10268_, _08013_);
  or _18647_ (_10270_, _10269_, _10267_);
  or _18648_ (_10271_, _08015_, word_in[26]);
  and _18649_ (_08873_, _10271_, _10270_);
  not _18650_ (_10272_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _18651_ (_10273_, _08028_, _10272_);
  and _18652_ (_10274_, _08028_, word_in[3]);
  nor _18653_ (_10275_, _10274_, _10273_);
  nor _18654_ (_10276_, _10275_, _08023_);
  and _18655_ (_10277_, _08023_, word_in[11]);
  or _18656_ (_10278_, _10277_, _10276_);
  and _18657_ (_10279_, _10278_, _08020_);
  and _18658_ (_10280_, _08712_, _08019_);
  or _18659_ (_10281_, _10280_, _08013_);
  or _18660_ (_10282_, _10281_, _10279_);
  or _18661_ (_10283_, _08015_, word_in[27]);
  and _18662_ (_08877_, _10283_, _10282_);
  and _18663_ (_10284_, _08608_, _08013_);
  and _18664_ (_10285_, _08028_, word_in[4]);
  not _18665_ (_10286_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _18666_ (_10287_, _08028_, _10286_);
  nor _18667_ (_10288_, _10287_, _10285_);
  nor _18668_ (_10289_, _10288_, _08023_);
  and _18669_ (_10290_, _08023_, word_in[12]);
  or _18670_ (_10291_, _10290_, _10289_);
  and _18671_ (_10292_, _10291_, _08020_);
  and _18672_ (_10293_, _08733_, _08019_);
  or _18673_ (_10294_, _10293_, _10292_);
  and _18674_ (_10295_, _10294_, _08015_);
  or _18675_ (_08879_, _10295_, _10284_);
  and _18676_ (_10296_, _08622_, _08013_);
  and _18677_ (_10297_, _08028_, word_in[5]);
  not _18678_ (_10298_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _18679_ (_10299_, _08028_, _10298_);
  nor _18680_ (_10300_, _10299_, _10297_);
  nor _18681_ (_10301_, _10300_, _08023_);
  and _18682_ (_10302_, _08023_, word_in[13]);
  or _18683_ (_10303_, _10302_, _10301_);
  and _18684_ (_10304_, _10303_, _08020_);
  and _18685_ (_10305_, _08746_, _08019_);
  or _18686_ (_10306_, _10305_, _10304_);
  and _18687_ (_10307_, _10306_, _08015_);
  or _18688_ (_08882_, _10307_, _10296_);
  and _18689_ (_10308_, _08624_, _08013_);
  not _18690_ (_10309_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _18691_ (_10310_, _08028_, _10309_);
  and _18692_ (_10311_, _08028_, word_in[6]);
  nor _18693_ (_10312_, _10311_, _10310_);
  nor _18694_ (_10313_, _10312_, _08023_);
  and _18695_ (_10314_, _08023_, word_in[14]);
  or _18696_ (_10315_, _10314_, _10313_);
  and _18697_ (_10316_, _10315_, _08020_);
  and _18698_ (_10317_, _08759_, _08019_);
  or _18699_ (_10318_, _10317_, _10316_);
  and _18700_ (_10320_, _10318_, _08015_);
  or _18701_ (_08887_, _10320_, _10308_);
  or _18702_ (_08889_, _06811_, _06831_);
  or _18703_ (_10321_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand _18704_ (_10322_, _07619_, _06324_);
  and _18705_ (_10323_, _10322_, _05141_);
  and _18706_ (_08991_, _10323_, _10321_);
  and _18707_ (_10324_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _18708_ (_10325_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _18709_ (_09143_, _10325_, _10324_);
  or _18710_ (_10326_, _05842_, _05840_);
  not _18711_ (_10327_, _05686_);
  nand _18712_ (_10328_, _05840_, _10327_);
  and _18713_ (_10329_, _10328_, _05656_);
  and _18714_ (_10330_, _10329_, _10326_);
  and _18715_ (_10331_, _06600_, ABINPUT000000[0]);
  and _18716_ (_10332_, _06606_, ABINPUT000[0]);
  or _18717_ (_10333_, _10332_, _10331_);
  nand _18718_ (_10334_, _05879_, _05846_);
  and _18719_ (_10335_, _05880_, _05844_);
  and _18720_ (_10336_, _10335_, _10334_);
  or _18721_ (_10337_, _10336_, _10333_);
  or _18722_ (_10338_, _10337_, _10330_);
  and _18723_ (_10339_, _10338_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _18724_ (_10341_, _05256_);
  and _18725_ (_10342_, _06877_, _10341_);
  and _18726_ (_10343_, _05266_, _05228_);
  and _18727_ (_10345_, _10343_, _05647_);
  and _18728_ (_10346_, _10345_, _10342_);
  not _18729_ (_10348_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and _18730_ (_10349_, _10348_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _18731_ (_10350_, _10349_, _10346_);
  or _18732_ (_10351_, _10350_, _10339_);
  and _18733_ (_10352_, _06018_, _05210_);
  and _18734_ (_10353_, _06733_, _05281_);
  and _18735_ (_10354_, _10353_, _10352_);
  not _18736_ (_10355_, _10354_);
  and _18737_ (_10356_, _05922_, _06620_);
  not _18738_ (_10357_, _06620_);
  nand _18739_ (_10358_, _10357_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand _18740_ (_10359_, _10358_, _10346_);
  or _18741_ (_10360_, _10359_, _10356_);
  and _18742_ (_10361_, _10360_, _10355_);
  and _18743_ (_10362_, _10361_, _10351_);
  nor _18744_ (_10363_, _10355_, _05560_);
  or _18745_ (_10364_, _10363_, _10362_);
  and _18746_ (_09170_, _10364_, _05141_);
  and _18747_ (_10365_, _10352_, _06733_);
  and _18748_ (_10366_, _10365_, _05281_);
  and _18749_ (_10367_, _10346_, _05288_);
  nand _18750_ (_10368_, _10367_, _05963_);
  or _18751_ (_10369_, _10367_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _18752_ (_10370_, _10369_, _10368_);
  or _18753_ (_10371_, _10370_, _10366_);
  nand _18754_ (_10372_, _10354_, _06178_);
  and _18755_ (_10373_, _10372_, _05141_);
  and _18756_ (_09173_, _10373_, _10371_);
  nor _18757_ (_10374_, _05209_, _06007_);
  nor _18758_ (_10375_, _10374_, _08469_);
  not _18759_ (_10376_, _10346_);
  or _18760_ (_10378_, _10376_, _10375_);
  and _18761_ (_10379_, _10378_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _18762_ (_10380_, _05922_, _08469_);
  and _18763_ (_10381_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _18764_ (_10383_, _10381_, _10380_);
  and _18765_ (_10384_, _10383_, _10346_);
  or _18766_ (_10385_, _10384_, _10379_);
  and _18767_ (_10386_, _10385_, _10355_);
  and _18768_ (_10387_, _10354_, _05522_);
  or _18769_ (_10389_, _10387_, _10386_);
  and _18770_ (_09564_, _10389_, _05141_);
  and _18771_ (_10390_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and _18772_ (_10391_, _05864_, _05844_);
  and _18773_ (_10392_, _05835_, _05656_);
  or _18774_ (_10393_, _10392_, _10391_);
  and _18775_ (_10394_, _10393_, _10390_);
  nand _18776_ (_10395_, _10390_, _06598_);
  and _18777_ (_10396_, _10395_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _18778_ (_10397_, _10396_, _10346_);
  or _18779_ (_10398_, _10397_, _10394_);
  or _18780_ (_10399_, _06207_, _07328_);
  nand _18781_ (_10400_, _10399_, _10346_);
  or _18782_ (_10401_, _10400_, _06208_);
  and _18783_ (_10402_, _10401_, _10398_);
  or _18784_ (_10403_, _10402_, _10354_);
  nand _18785_ (_10404_, _10354_, _06244_);
  and _18786_ (_10405_, _10404_, _05141_);
  and _18787_ (_09569_, _10405_, _10403_);
  and _18788_ (_10407_, _05275_, _06007_);
  and _18789_ (_10408_, _10346_, _10407_);
  nand _18790_ (_10410_, _10408_, _05963_);
  or _18791_ (_10411_, _10408_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _18792_ (_10413_, _10411_, _10410_);
  or _18793_ (_10414_, _10413_, _10366_);
  or _18794_ (_10415_, _10355_, _06004_);
  and _18795_ (_10416_, _10415_, _05141_);
  and _18796_ (_09572_, _10416_, _10414_);
  or _18797_ (_10418_, _06389_, _07117_);
  or _18798_ (_10419_, _06270_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _18799_ (_10420_, _10419_, _05141_);
  and _18800_ (_09689_, _10420_, _10418_);
  and _18801_ (_10421_, _07758_, word_in[0]);
  nand _18802_ (_10422_, _07613_, _09576_);
  or _18803_ (_10423_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _18804_ (_10424_, _10423_, _10422_);
  and _18805_ (_10425_, _10424_, _07666_);
  nand _18806_ (_10426_, _07613_, _09794_);
  or _18807_ (_10427_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _18808_ (_10428_, _10427_, _10426_);
  and _18809_ (_10429_, _10428_, _07643_);
  nand _18810_ (_10430_, _07613_, _10010_);
  or _18811_ (_10431_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _18812_ (_10432_, _10431_, _10430_);
  and _18813_ (_10433_, _10432_, _07640_);
  or _18814_ (_10434_, _10433_, _10429_);
  or _18815_ (_10435_, _10434_, _10425_);
  nand _18816_ (_10436_, _07613_, _10234_);
  or _18817_ (_10438_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _18818_ (_10439_, _10438_, _10436_);
  and _18819_ (_10440_, _10439_, _07650_);
  or _18820_ (_10441_, _10440_, _07676_);
  or _18821_ (_10442_, _10441_, _10435_);
  nand _18822_ (_10443_, _07613_, _08672_);
  or _18823_ (_10444_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _18824_ (_10445_, _10444_, _10443_);
  and _18825_ (_10446_, _10445_, _07666_);
  nand _18826_ (_10447_, _07613_, _08924_);
  or _18827_ (_10448_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _18828_ (_10449_, _10448_, _10447_);
  and _18829_ (_10450_, _10449_, _07643_);
  nand _18830_ (_10451_, _07613_, _09133_);
  or _18831_ (_10452_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _18832_ (_10453_, _10452_, _10451_);
  and _18833_ (_10454_, _10453_, _07640_);
  or _18834_ (_10455_, _10454_, _10450_);
  or _18835_ (_10456_, _10455_, _10446_);
  nand _18836_ (_10457_, _07613_, _09343_);
  or _18837_ (_10459_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _18838_ (_10460_, _10459_, _10457_);
  and _18839_ (_10462_, _10460_, _07650_);
  or _18840_ (_10463_, _10462_, _07626_);
  or _18841_ (_10464_, _10463_, _10456_);
  and _18842_ (_10465_, _10464_, _10442_);
  and _18843_ (_10466_, _10465_, _07705_);
  or _18844_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _10466_, _10421_);
  and _18845_ (_10467_, _07758_, word_in[1]);
  nand _18846_ (_10468_, _07613_, _09592_);
  or _18847_ (_10469_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _18848_ (_10470_, _10469_, _10468_);
  and _18849_ (_10471_, _10470_, _07666_);
  nand _18850_ (_10472_, _07613_, _09806_);
  or _18851_ (_10473_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _18852_ (_10474_, _10473_, _10472_);
  and _18853_ (_10475_, _10474_, _07643_);
  nand _18854_ (_10477_, _07613_, _10026_);
  or _18855_ (_10478_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _18856_ (_10479_, _10478_, _10477_);
  and _18857_ (_10480_, _10479_, _07640_);
  or _18858_ (_10481_, _10480_, _10475_);
  or _18859_ (_10482_, _10481_, _10471_);
  nand _18860_ (_10483_, _07613_, _10248_);
  or _18861_ (_10484_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _18862_ (_10485_, _10484_, _10483_);
  and _18863_ (_10486_, _10485_, _07650_);
  or _18864_ (_10487_, _10486_, _07676_);
  or _18865_ (_10488_, _10487_, _10482_);
  nand _18866_ (_10490_, _07613_, _08685_);
  or _18867_ (_10491_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _18868_ (_10493_, _10491_, _10490_);
  and _18869_ (_10495_, _10493_, _07666_);
  nand _18870_ (_10496_, _07613_, _08937_);
  or _18871_ (_10497_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _18872_ (_10498_, _10497_, _10496_);
  and _18873_ (_10500_, _10498_, _07643_);
  nand _18874_ (_10501_, _07613_, _09150_);
  or _18875_ (_10502_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _18876_ (_10504_, _10502_, _10501_);
  and _18877_ (_10505_, _10504_, _07640_);
  or _18878_ (_10506_, _10505_, _10500_);
  or _18879_ (_10507_, _10506_, _10495_);
  nand _18880_ (_10508_, _07613_, _09354_);
  or _18881_ (_10509_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _18882_ (_10511_, _10509_, _10508_);
  and _18883_ (_10512_, _10511_, _07650_);
  or _18884_ (_10513_, _10512_, _07626_);
  or _18885_ (_10514_, _10513_, _10507_);
  and _18886_ (_10515_, _10514_, _10488_);
  and _18887_ (_10516_, _10515_, _07705_);
  or _18888_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _10516_, _10467_);
  and _18889_ (_10517_, _07758_, word_in[2]);
  nand _18890_ (_10518_, _07613_, _09604_);
  or _18891_ (_10519_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _18892_ (_10520_, _10519_, _10518_);
  and _18893_ (_10521_, _10520_, _07666_);
  nand _18894_ (_10522_, _07613_, _10038_);
  or _18895_ (_10523_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _18896_ (_10524_, _10523_, _10522_);
  and _18897_ (_10525_, _10524_, _07640_);
  nand _18898_ (_10526_, _07613_, _09820_);
  or _18899_ (_10527_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _18900_ (_10528_, _10527_, _10526_);
  and _18901_ (_10530_, _10528_, _07643_);
  or _18902_ (_10531_, _10530_, _10525_);
  or _18903_ (_10532_, _10531_, _10521_);
  nand _18904_ (_10533_, _07613_, _10260_);
  or _18905_ (_10534_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _18906_ (_10535_, _10534_, _10533_);
  and _18907_ (_10536_, _10535_, _07650_);
  or _18908_ (_10537_, _10536_, _07676_);
  or _18909_ (_10538_, _10537_, _10532_);
  nand _18910_ (_10539_, _07613_, _08700_);
  or _18911_ (_10541_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _18912_ (_10542_, _10541_, _10539_);
  and _18913_ (_10543_, _10542_, _07666_);
  nand _18914_ (_10544_, _07613_, _08949_);
  or _18915_ (_10545_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _18916_ (_10546_, _10545_, _10544_);
  and _18917_ (_10547_, _10546_, _07643_);
  nand _18918_ (_10548_, _07613_, _09161_);
  or _18919_ (_10549_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _18920_ (_10550_, _10549_, _10548_);
  and _18921_ (_10551_, _10550_, _07640_);
  or _18922_ (_10552_, _10551_, _10547_);
  or _18923_ (_10553_, _10552_, _10543_);
  nand _18924_ (_10554_, _07613_, _09366_);
  or _18925_ (_10556_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _18926_ (_10558_, _10556_, _10554_);
  and _18927_ (_10559_, _10558_, _07650_);
  or _18928_ (_10560_, _10559_, _07626_);
  or _18929_ (_10561_, _10560_, _10553_);
  and _18930_ (_10562_, _10561_, _10538_);
  and _18931_ (_10563_, _10562_, _07705_);
  or _18932_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _10563_, _10517_);
  and _18933_ (_10564_, _07758_, word_in[3]);
  nand _18934_ (_10565_, _07613_, _09617_);
  or _18935_ (_10566_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _18936_ (_10567_, _10566_, _10565_);
  and _18937_ (_10568_, _10567_, _07666_);
  nand _18938_ (_10569_, _07613_, _10050_);
  or _18939_ (_10571_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _18940_ (_10572_, _10571_, _10569_);
  and _18941_ (_10573_, _10572_, _07640_);
  nand _18942_ (_10574_, _07613_, _09832_);
  or _18943_ (_10576_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _18944_ (_10577_, _10576_, _10574_);
  and _18945_ (_10578_, _10577_, _07643_);
  or _18946_ (_10579_, _10578_, _10573_);
  or _18947_ (_10580_, _10579_, _10568_);
  nand _18948_ (_10581_, _07613_, _10272_);
  or _18949_ (_10582_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _18950_ (_10584_, _10582_, _10581_);
  and _18951_ (_10585_, _10584_, _07650_);
  or _18952_ (_10586_, _10585_, _07676_);
  or _18953_ (_10587_, _10586_, _10580_);
  nand _18954_ (_10588_, _07613_, _08714_);
  or _18955_ (_10589_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _18956_ (_10590_, _10589_, _10588_);
  and _18957_ (_10591_, _10590_, _07666_);
  nand _18958_ (_10592_, _07613_, _08960_);
  or _18959_ (_10593_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _18960_ (_10594_, _10593_, _10592_);
  and _18961_ (_10595_, _10594_, _07643_);
  nand _18962_ (_10596_, _07613_, _09175_);
  or _18963_ (_10597_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _18964_ (_10598_, _10597_, _10596_);
  and _18965_ (_10599_, _10598_, _07640_);
  or _18966_ (_10600_, _10599_, _10595_);
  or _18967_ (_10601_, _10600_, _10591_);
  nand _18968_ (_10602_, _07613_, _09378_);
  or _18969_ (_10603_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _18970_ (_10604_, _10603_, _10602_);
  and _18971_ (_10605_, _10604_, _07650_);
  or _18972_ (_10606_, _10605_, _07626_);
  or _18973_ (_10607_, _10606_, _10601_);
  and _18974_ (_10608_, _10607_, _10587_);
  and _18975_ (_10609_, _10608_, _07705_);
  or _18976_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _10609_, _10564_);
  and _18977_ (_10611_, _07758_, word_in[4]);
  nand _18978_ (_10612_, _07613_, _09628_);
  or _18979_ (_10613_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _18980_ (_10614_, _10613_, _10612_);
  and _18981_ (_10615_, _10614_, _07666_);
  nand _18982_ (_10616_, _07613_, _09845_);
  or _18983_ (_10617_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _18984_ (_10618_, _10617_, _10616_);
  and _18985_ (_10619_, _10618_, _07643_);
  nand _18986_ (_10620_, _07613_, _10071_);
  or _18987_ (_10621_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _18988_ (_10622_, _10621_, _10620_);
  and _18989_ (_10623_, _10622_, _07640_);
  or _18990_ (_10624_, _10623_, _10619_);
  or _18991_ (_10625_, _10624_, _10615_);
  nand _18992_ (_10626_, _07613_, _10286_);
  or _18993_ (_10627_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _18994_ (_10628_, _10627_, _10626_);
  and _18995_ (_10629_, _10628_, _07650_);
  or _18996_ (_10630_, _10629_, _07676_);
  or _18997_ (_10631_, _10630_, _10625_);
  nand _18998_ (_10632_, _07613_, _08726_);
  or _18999_ (_10633_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _19000_ (_10634_, _10633_, _10632_);
  and _19001_ (_10635_, _10634_, _07666_);
  nand _19002_ (_10636_, _07613_, _08972_);
  or _19003_ (_10637_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _19004_ (_10638_, _10637_, _10636_);
  and _19005_ (_10639_, _10638_, _07643_);
  nand _19006_ (_10641_, _07613_, _09186_);
  or _19007_ (_10642_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _19008_ (_10643_, _10642_, _10641_);
  and _19009_ (_10644_, _10643_, _07640_);
  or _19010_ (_10645_, _10644_, _10639_);
  or _19011_ (_10646_, _10645_, _10635_);
  nand _19012_ (_10648_, _07613_, _09390_);
  or _19013_ (_10649_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _19014_ (_10650_, _10649_, _10648_);
  and _19015_ (_10651_, _10650_, _07650_);
  or _19016_ (_10652_, _10651_, _07626_);
  or _19017_ (_10653_, _10652_, _10646_);
  and _19018_ (_10654_, _10653_, _10631_);
  and _19019_ (_10655_, _10654_, _07705_);
  or _19020_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _10655_, _10611_);
  and _19021_ (_10657_, _07758_, word_in[5]);
  nand _19022_ (_10658_, _07613_, _09858_);
  or _19023_ (_10659_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _19024_ (_10660_, _10659_, _10658_);
  and _19025_ (_10661_, _10660_, _07643_);
  nand _19026_ (_10662_, _07613_, _10084_);
  or _19027_ (_10663_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _19028_ (_10664_, _10663_, _10662_);
  and _19029_ (_10665_, _10664_, _07640_);
  nand _19030_ (_10666_, _07613_, _09640_);
  or _19031_ (_10667_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _19032_ (_10668_, _10667_, _10666_);
  and _19033_ (_10669_, _10668_, _07666_);
  or _19034_ (_10670_, _10669_, _10665_);
  or _19035_ (_10671_, _10670_, _10661_);
  nand _19036_ (_10672_, _07613_, _10298_);
  or _19037_ (_10673_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _19038_ (_10674_, _10673_, _10672_);
  and _19039_ (_10675_, _10674_, _07650_);
  or _19040_ (_10676_, _10675_, _07676_);
  or _19041_ (_10677_, _10676_, _10671_);
  nand _19042_ (_10678_, _07613_, _08984_);
  or _19043_ (_10679_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _19044_ (_10680_, _10679_, _10678_);
  and _19045_ (_10681_, _10680_, _07643_);
  nand _19046_ (_10682_, _07613_, _08739_);
  or _19047_ (_10683_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _19048_ (_10684_, _10683_, _10682_);
  and _19049_ (_10685_, _10684_, _07666_);
  nand _19050_ (_10686_, _07613_, _09198_);
  or _19051_ (_10687_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _19052_ (_10688_, _10687_, _10686_);
  and _19053_ (_10689_, _10688_, _07640_);
  or _19054_ (_10690_, _10689_, _10685_);
  or _19055_ (_10691_, _10690_, _10681_);
  nand _19056_ (_10692_, _07613_, _09402_);
  or _19057_ (_10693_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _19058_ (_10694_, _10693_, _10692_);
  and _19059_ (_10695_, _10694_, _07650_);
  or _19060_ (_10696_, _10695_, _07626_);
  or _19061_ (_10697_, _10696_, _10691_);
  and _19062_ (_10699_, _10697_, _10677_);
  and _19063_ (_10700_, _10699_, _07705_);
  or _19064_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _10700_, _10657_);
  and _19065_ (_10701_, _07758_, word_in[6]);
  nand _19066_ (_10702_, _07613_, _09872_);
  or _19067_ (_10703_, _07613_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _19068_ (_10704_, _10703_, _10702_);
  and _19069_ (_10705_, _10704_, _07643_);
  nand _19070_ (_10706_, _07613_, _10096_);
  or _19071_ (_10707_, _07613_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _19072_ (_10708_, _10707_, _10706_);
  and _19073_ (_10709_, _10708_, _07640_);
  nand _19074_ (_10710_, _07613_, _09652_);
  or _19075_ (_10711_, _07613_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _19076_ (_10712_, _10711_, _10710_);
  and _19077_ (_10713_, _10712_, _07666_);
  or _19078_ (_10714_, _10713_, _10709_);
  or _19079_ (_10716_, _10714_, _10705_);
  nand _19080_ (_10717_, _07613_, _10309_);
  or _19081_ (_10719_, _07613_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _19082_ (_10720_, _10719_, _10717_);
  and _19083_ (_10721_, _10720_, _07650_);
  or _19084_ (_10722_, _10721_, _07676_);
  or _19085_ (_10723_, _10722_, _10716_);
  nand _19086_ (_10724_, _07613_, _08998_);
  or _19087_ (_10725_, _07613_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _19088_ (_10726_, _10725_, _10724_);
  and _19089_ (_10727_, _10726_, _07643_);
  nand _19090_ (_10728_, _07613_, _08752_);
  or _19091_ (_10729_, _07613_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _19092_ (_10730_, _10729_, _10728_);
  and _19093_ (_10731_, _10730_, _07666_);
  nand _19094_ (_10732_, _07613_, _09211_);
  or _19095_ (_10733_, _07613_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _19096_ (_10734_, _10733_, _10732_);
  and _19097_ (_10735_, _10734_, _07640_);
  or _19098_ (_10736_, _10735_, _10731_);
  or _19099_ (_10737_, _10736_, _10727_);
  nand _19100_ (_10738_, _07613_, _09413_);
  or _19101_ (_10739_, _07613_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _19102_ (_10740_, _10739_, _10738_);
  and _19103_ (_10741_, _10740_, _07650_);
  or _19104_ (_10743_, _10741_, _07626_);
  or _19105_ (_10744_, _10743_, _10737_);
  and _19106_ (_10745_, _10744_, _10723_);
  and _19107_ (_10746_, _10745_, _07705_);
  or _19108_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _10746_, _10701_);
  and _19109_ (_10748_, _07819_, word_in[8]);
  nand _19110_ (_10749_, _07613_, _08790_);
  or _19111_ (_10751_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _19112_ (_10752_, _10751_, _10749_);
  and _19113_ (_10753_, _10752_, _07821_);
  nand _19114_ (_10754_, _07613_, _08535_);
  or _19115_ (_10755_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _19116_ (_10756_, _10755_, _10754_);
  and _19117_ (_10757_, _10756_, _07820_);
  or _19118_ (_10758_, _10757_, _10753_);
  and _19119_ (_10759_, _10758_, _07781_);
  nand _19120_ (_10760_, _07613_, _09680_);
  or _19121_ (_10761_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _19122_ (_10762_, _10761_, _10760_);
  and _19123_ (_10763_, _10762_, _07821_);
  nand _19124_ (_10764_, _07613_, _09468_);
  or _19125_ (_10765_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _19126_ (_10766_, _10765_, _10764_);
  and _19127_ (_10767_, _10766_, _07820_);
  or _19128_ (_10768_, _10767_, _10763_);
  and _19129_ (_10769_, _10768_, _07783_);
  nand _19130_ (_10770_, _07613_, _09236_);
  or _19131_ (_10771_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _19132_ (_10772_, _10771_, _10770_);
  and _19133_ (_10773_, _10772_, _07821_);
  nand _19134_ (_10774_, _07613_, _09025_);
  or _19135_ (_10775_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _19136_ (_10776_, _10775_, _10774_);
  and _19137_ (_10777_, _10776_, _07820_);
  or _19138_ (_10778_, _10777_, _10773_);
  and _19139_ (_10779_, _10778_, _07807_);
  nand _19140_ (_10780_, _07613_, _10131_);
  or _19141_ (_10781_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _19142_ (_10782_, _10781_, _10780_);
  and _19143_ (_10783_, _10782_, _07821_);
  nand _19144_ (_10784_, _07613_, _09908_);
  or _19145_ (_10785_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _19146_ (_10786_, _10785_, _10784_);
  and _19147_ (_10787_, _10786_, _07820_);
  or _19148_ (_10788_, _10787_, _10783_);
  and _19149_ (_10789_, _10788_, _07811_);
  or _19150_ (_10790_, _10789_, _10779_);
  or _19151_ (_10791_, _10790_, _10769_);
  nor _19152_ (_10793_, _10791_, _10759_);
  nor _19153_ (_10794_, _10793_, _07819_);
  or _19154_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _10794_, _10748_);
  and _19155_ (_10795_, _07819_, word_in[9]);
  nand _19156_ (_10796_, _07613_, _08810_);
  or _19157_ (_10797_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _19158_ (_10798_, _10797_, _10796_);
  and _19159_ (_10799_, _10798_, _07821_);
  nand _19160_ (_10801_, _07613_, _08554_);
  or _19161_ (_10802_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _19162_ (_10803_, _10802_, _10801_);
  and _19163_ (_10804_, _10803_, _07820_);
  or _19164_ (_10805_, _10804_, _10799_);
  and _19165_ (_10806_, _10805_, _07781_);
  nand _19166_ (_10807_, _07613_, _09695_);
  or _19167_ (_10808_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _19168_ (_10809_, _10808_, _10807_);
  and _19169_ (_10810_, _10809_, _07821_);
  nand _19170_ (_10811_, _07613_, _09483_);
  or _19171_ (_10812_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _19172_ (_10813_, _10812_, _10811_);
  and _19173_ (_10814_, _10813_, _07820_);
  or _19174_ (_10815_, _10814_, _10810_);
  and _19175_ (_10816_, _10815_, _07783_);
  nand _19176_ (_10817_, _07613_, _09253_);
  or _19177_ (_10818_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _19178_ (_10819_, _10818_, _10817_);
  and _19179_ (_10820_, _10819_, _07821_);
  nand _19180_ (_10821_, _07613_, _09043_);
  or _19181_ (_10822_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _19182_ (_10823_, _10822_, _10821_);
  and _19183_ (_10824_, _10823_, _07820_);
  or _19184_ (_10825_, _10824_, _10820_);
  and _19185_ (_10826_, _10825_, _07807_);
  nand _19186_ (_10827_, _07613_, _10146_);
  or _19187_ (_10828_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _19188_ (_10829_, _10828_, _10827_);
  and _19189_ (_10830_, _10829_, _07821_);
  nand _19190_ (_10831_, _07613_, _09924_);
  or _19191_ (_10832_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _19192_ (_10833_, _10832_, _10831_);
  and _19193_ (_10834_, _10833_, _07820_);
  or _19194_ (_10835_, _10834_, _10830_);
  and _19195_ (_10836_, _10835_, _07811_);
  or _19196_ (_10837_, _10836_, _10826_);
  or _19197_ (_10838_, _10837_, _10816_);
  nor _19198_ (_10839_, _10838_, _10806_);
  nor _19199_ (_10840_, _10839_, _07819_);
  or _19200_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _10840_, _10795_);
  and _19201_ (_10841_, _07819_, word_in[10]);
  nand _19202_ (_10842_, _07613_, _08823_);
  or _19203_ (_10843_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _19204_ (_10844_, _10843_, _10842_);
  and _19205_ (_10845_, _10844_, _07821_);
  nand _19206_ (_10846_, _07613_, _08570_);
  or _19207_ (_10847_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _19208_ (_10848_, _10847_, _10846_);
  and _19209_ (_10849_, _10848_, _07820_);
  or _19210_ (_10850_, _10849_, _10845_);
  and _19211_ (_10851_, _10850_, _07781_);
  nand _19212_ (_10852_, _07613_, _09708_);
  or _19213_ (_10853_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _19214_ (_10854_, _10853_, _10852_);
  and _19215_ (_10855_, _10854_, _07821_);
  nand _19216_ (_10856_, _07613_, _09495_);
  or _19217_ (_10857_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _19218_ (_10858_, _10857_, _10856_);
  and _19219_ (_10859_, _10858_, _07820_);
  or _19220_ (_10860_, _10859_, _10855_);
  and _19221_ (_10861_, _10860_, _07783_);
  nand _19222_ (_10862_, _07613_, _09264_);
  or _19223_ (_10863_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _19224_ (_10864_, _10863_, _10862_);
  and _19225_ (_10865_, _10864_, _07821_);
  nand _19226_ (_10866_, _07613_, _09055_);
  or _19227_ (_10867_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _19228_ (_10868_, _10867_, _10866_);
  and _19229_ (_10869_, _10868_, _07820_);
  or _19230_ (_10870_, _10869_, _10865_);
  and _19231_ (_10872_, _10870_, _07807_);
  nand _19232_ (_10873_, _07613_, _10159_);
  or _19233_ (_10874_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _19234_ (_10875_, _10874_, _10873_);
  and _19235_ (_10876_, _10875_, _07821_);
  nand _19236_ (_10877_, _07613_, _09936_);
  or _19237_ (_10878_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _19238_ (_10879_, _10878_, _10877_);
  and _19239_ (_10880_, _10879_, _07820_);
  or _19240_ (_10881_, _10880_, _10876_);
  and _19241_ (_10882_, _10881_, _07811_);
  or _19242_ (_10883_, _10882_, _10872_);
  or _19243_ (_10884_, _10883_, _10861_);
  nor _19244_ (_10885_, _10884_, _10851_);
  nor _19245_ (_10886_, _10885_, _07819_);
  or _19246_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _10886_, _10841_);
  and _19247_ (_10888_, _07819_, word_in[11]);
  nand _19248_ (_10889_, _07613_, _08836_);
  or _19249_ (_10891_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _19250_ (_10892_, _10891_, _10889_);
  and _19251_ (_10893_, _10892_, _07821_);
  nand _19252_ (_10894_, _07613_, _08584_);
  or _19253_ (_10895_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _19254_ (_10896_, _10895_, _10894_);
  and _19255_ (_10897_, _10896_, _07820_);
  or _19256_ (_10898_, _10897_, _10893_);
  and _19257_ (_10899_, _10898_, _07781_);
  nand _19258_ (_10900_, _07613_, _09720_);
  or _19259_ (_10901_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _19260_ (_10902_, _10901_, _10900_);
  and _19261_ (_10903_, _10902_, _07821_);
  nand _19262_ (_10904_, _07613_, _09507_);
  or _19263_ (_10905_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _19264_ (_10906_, _10905_, _10904_);
  and _19265_ (_10907_, _10906_, _07820_);
  or _19266_ (_10908_, _10907_, _10903_);
  and _19267_ (_10909_, _10908_, _07783_);
  nand _19268_ (_10910_, _07613_, _09276_);
  or _19269_ (_10911_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _19270_ (_10912_, _10911_, _10910_);
  and _19271_ (_10913_, _10912_, _07821_);
  nand _19272_ (_10914_, _07613_, _09067_);
  or _19273_ (_10915_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _19274_ (_10916_, _10915_, _10914_);
  and _19275_ (_10917_, _10916_, _07820_);
  or _19276_ (_10918_, _10917_, _10913_);
  and _19277_ (_10919_, _10918_, _07807_);
  nand _19278_ (_10920_, _07613_, _10172_);
  or _19279_ (_10921_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _19280_ (_10922_, _10921_, _10920_);
  and _19281_ (_10923_, _10922_, _07821_);
  nand _19282_ (_10924_, _07613_, _09948_);
  or _19283_ (_10925_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _19284_ (_10926_, _10925_, _10924_);
  and _19285_ (_10927_, _10926_, _07820_);
  or _19286_ (_10928_, _10927_, _10923_);
  and _19287_ (_10929_, _10928_, _07811_);
  or _19288_ (_10930_, _10929_, _10919_);
  or _19289_ (_10931_, _10930_, _10909_);
  nor _19290_ (_10932_, _10931_, _10899_);
  nor _19291_ (_10933_, _10932_, _07819_);
  or _19292_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _10933_, _10888_);
  and _19293_ (_10934_, _07819_, word_in[12]);
  nand _19294_ (_10935_, _07613_, _08850_);
  or _19295_ (_10937_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _19296_ (_10938_, _10937_, _10935_);
  and _19297_ (_10939_, _10938_, _07821_);
  nand _19298_ (_10941_, _07613_, _08596_);
  or _19299_ (_10942_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _19300_ (_10944_, _10942_, _10941_);
  and _19301_ (_10945_, _10944_, _07820_);
  or _19302_ (_10946_, _10945_, _10939_);
  and _19303_ (_10947_, _10946_, _07781_);
  nand _19304_ (_10948_, _07613_, _09731_);
  or _19305_ (_10949_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _19306_ (_10950_, _10949_, _10948_);
  and _19307_ (_10951_, _10950_, _07821_);
  nand _19308_ (_10952_, _07613_, _09519_);
  or _19309_ (_10953_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _19310_ (_10954_, _10953_, _10952_);
  and _19311_ (_10955_, _10954_, _07820_);
  or _19312_ (_10956_, _10955_, _10951_);
  and _19313_ (_10957_, _10956_, _07783_);
  nand _19314_ (_10958_, _07613_, _09289_);
  or _19315_ (_10959_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _19316_ (_10960_, _10959_, _10958_);
  and _19317_ (_10961_, _10960_, _07821_);
  nand _19318_ (_10962_, _07613_, _09079_);
  or _19319_ (_10963_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _19320_ (_10964_, _10963_, _10962_);
  and _19321_ (_10965_, _10964_, _07820_);
  or _19322_ (_10966_, _10965_, _10961_);
  and _19323_ (_10967_, _10966_, _07807_);
  nand _19324_ (_10968_, _07613_, _10184_);
  or _19325_ (_10969_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _19326_ (_10970_, _10969_, _10968_);
  and _19327_ (_10971_, _10970_, _07821_);
  nand _19328_ (_10972_, _07613_, _09960_);
  or _19329_ (_10973_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _19330_ (_10974_, _10973_, _10972_);
  and _19331_ (_10975_, _10974_, _07820_);
  or _19332_ (_10976_, _10975_, _10971_);
  and _19333_ (_10977_, _10976_, _07811_);
  or _19334_ (_10978_, _10977_, _10967_);
  or _19335_ (_10979_, _10978_, _10957_);
  nor _19336_ (_10980_, _10979_, _10947_);
  nor _19337_ (_10981_, _10980_, _07819_);
  or _19338_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _10981_, _10934_);
  and _19339_ (_10982_, _07819_, word_in[13]);
  nand _19340_ (_10983_, _07613_, _08862_);
  or _19341_ (_10984_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _19342_ (_10985_, _10984_, _10983_);
  and _19343_ (_10987_, _10985_, _07821_);
  nand _19344_ (_10988_, _07613_, _08610_);
  or _19345_ (_10989_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _19346_ (_10990_, _10989_, _10988_);
  and _19347_ (_10991_, _10990_, _07820_);
  or _19348_ (_10992_, _10991_, _10987_);
  and _19349_ (_10993_, _10992_, _07781_);
  nand _19350_ (_10994_, _07613_, _09744_);
  or _19351_ (_10995_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _19352_ (_10996_, _10995_, _10994_);
  and _19353_ (_10997_, _10996_, _07821_);
  nand _19354_ (_10998_, _07613_, _09531_);
  or _19355_ (_10999_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _19356_ (_11000_, _10999_, _10998_);
  and _19357_ (_11001_, _11000_, _07820_);
  or _19358_ (_11002_, _11001_, _10997_);
  and _19359_ (_11003_, _11002_, _07783_);
  nand _19360_ (_11004_, _07613_, _09301_);
  or _19361_ (_11005_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _19362_ (_11006_, _11005_, _11004_);
  and _19363_ (_11007_, _11006_, _07821_);
  nand _19364_ (_11008_, _07613_, _09091_);
  or _19365_ (_11009_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _19366_ (_11010_, _11009_, _11008_);
  and _19367_ (_11011_, _11010_, _07820_);
  or _19368_ (_11012_, _11011_, _11007_);
  and _19369_ (_11013_, _11012_, _07807_);
  nand _19370_ (_11014_, _07613_, _10197_);
  or _19371_ (_11015_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _19372_ (_11016_, _11015_, _11014_);
  and _19373_ (_11017_, _11016_, _07821_);
  nand _19374_ (_11018_, _07613_, _09972_);
  or _19375_ (_11019_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _19376_ (_11020_, _11019_, _11018_);
  and _19377_ (_11021_, _11020_, _07820_);
  or _19378_ (_11022_, _11021_, _11017_);
  and _19379_ (_11023_, _11022_, _07811_);
  or _19380_ (_11024_, _11023_, _11013_);
  or _19381_ (_11025_, _11024_, _11003_);
  nor _19382_ (_11026_, _11025_, _10993_);
  nor _19383_ (_11027_, _11026_, _07819_);
  or _19384_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _11027_, _10982_);
  and _19385_ (_11028_, _07819_, word_in[14]);
  nand _19386_ (_11029_, _07613_, _08890_);
  or _19387_ (_11031_, _07613_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _19388_ (_11032_, _11031_, _11029_);
  and _19389_ (_11033_, _11032_, _07821_);
  nand _19390_ (_11035_, _07613_, _08626_);
  or _19391_ (_11036_, _07613_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _19392_ (_11037_, _11036_, _11035_);
  and _19393_ (_11038_, _11037_, _07820_);
  or _19394_ (_11039_, _11038_, _11033_);
  and _19395_ (_11040_, _11039_, _07781_);
  nand _19396_ (_11041_, _07613_, _09756_);
  or _19397_ (_11042_, _07613_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _19398_ (_11043_, _11042_, _11041_);
  and _19399_ (_11044_, _11043_, _07821_);
  nand _19400_ (_11045_, _07613_, _09543_);
  or _19401_ (_11046_, _07613_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _19402_ (_11047_, _11046_, _11045_);
  and _19403_ (_11048_, _11047_, _07820_);
  or _19404_ (_11049_, _11048_, _11044_);
  and _19405_ (_11050_, _11049_, _07783_);
  nand _19406_ (_11051_, _07613_, _09313_);
  or _19407_ (_11052_, _07613_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _19408_ (_11053_, _11052_, _11051_);
  and _19409_ (_11054_, _11053_, _07821_);
  nand _19410_ (_11055_, _07613_, _09103_);
  or _19411_ (_11056_, _07613_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _19412_ (_11057_, _11056_, _11055_);
  and _19413_ (_11058_, _11057_, _07820_);
  or _19414_ (_11059_, _11058_, _11054_);
  and _19415_ (_11060_, _11059_, _07807_);
  nand _19416_ (_11061_, _07613_, _10209_);
  or _19417_ (_11062_, _07613_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _19418_ (_11064_, _11062_, _11061_);
  and _19419_ (_11065_, _11064_, _07821_);
  nand _19420_ (_11066_, _07613_, _09984_);
  or _19421_ (_11067_, _07613_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _19422_ (_11069_, _11067_, _11066_);
  and _19423_ (_11070_, _11069_, _07820_);
  or _19424_ (_11071_, _11070_, _11065_);
  and _19425_ (_11072_, _11071_, _07811_);
  or _19426_ (_11073_, _11072_, _11060_);
  or _19427_ (_11074_, _11073_, _11050_);
  nor _19428_ (_11075_, _11074_, _11040_);
  nor _19429_ (_11076_, _11075_, _07819_);
  or _19430_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _11076_, _11028_);
  and _19431_ (_11078_, _07917_, word_in[16]);
  and _19432_ (_11079_, _10453_, _07643_);
  and _19433_ (_11080_, _10445_, _07650_);
  or _19434_ (_11081_, _11080_, _11079_);
  and _19435_ (_11082_, _10460_, _07640_);
  and _19436_ (_11083_, _10449_, _07666_);
  or _19437_ (_11084_, _11083_, _11082_);
  or _19438_ (_11085_, _11084_, _11081_);
  or _19439_ (_11086_, _11085_, _07888_);
  and _19440_ (_11087_, _10424_, _07650_);
  and _19441_ (_11088_, _10439_, _07640_);
  or _19442_ (_11089_, _11088_, _11087_);
  and _19443_ (_11090_, _10432_, _07643_);
  and _19444_ (_11091_, _10428_, _07666_);
  or _19445_ (_11092_, _11091_, _11090_);
  or _19446_ (_11093_, _11092_, _11089_);
  or _19447_ (_11095_, _11093_, _07927_);
  nand _19448_ (_11096_, _11095_, _11086_);
  nor _19449_ (_11097_, _11096_, _07917_);
  or _19450_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _11097_, _11078_);
  and _19451_ (_11099_, _07917_, word_in[17]);
  and _19452_ (_11101_, _10504_, _07643_);
  and _19453_ (_11102_, _10493_, _07650_);
  or _19454_ (_11103_, _11102_, _11101_);
  and _19455_ (_11105_, _10511_, _07640_);
  and _19456_ (_11106_, _10498_, _07666_);
  or _19457_ (_11108_, _11106_, _11105_);
  or _19458_ (_11109_, _11108_, _11103_);
  or _19459_ (_11110_, _11109_, _07888_);
  and _19460_ (_11111_, _10470_, _07650_);
  and _19461_ (_11112_, _10485_, _07640_);
  or _19462_ (_11113_, _11112_, _11111_);
  and _19463_ (_11114_, _10479_, _07643_);
  and _19464_ (_11115_, _10474_, _07666_);
  or _19465_ (_11116_, _11115_, _11114_);
  or _19466_ (_11117_, _11116_, _11113_);
  or _19467_ (_11118_, _11117_, _07927_);
  nand _19468_ (_11119_, _11118_, _11110_);
  nor _19469_ (_11120_, _11119_, _07917_);
  or _19470_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _11120_, _11099_);
  and _19471_ (_11121_, _07917_, word_in[18]);
  and _19472_ (_11122_, _10542_, _07650_);
  and _19473_ (_11123_, _10558_, _07640_);
  or _19474_ (_11124_, _11123_, _11122_);
  and _19475_ (_11125_, _10550_, _07643_);
  and _19476_ (_11126_, _10546_, _07666_);
  or _19477_ (_11127_, _11126_, _11125_);
  or _19478_ (_11128_, _11127_, _11124_);
  or _19479_ (_11129_, _11128_, _07888_);
  and _19480_ (_11130_, _10524_, _07643_);
  and _19481_ (_11131_, _10520_, _07650_);
  or _19482_ (_11132_, _11131_, _11130_);
  and _19483_ (_11133_, _10535_, _07640_);
  and _19484_ (_11134_, _10528_, _07666_);
  or _19485_ (_11135_, _11134_, _11133_);
  or _19486_ (_11136_, _11135_, _11132_);
  or _19487_ (_11137_, _11136_, _07927_);
  nand _19488_ (_11138_, _11137_, _11129_);
  nor _19489_ (_11139_, _11138_, _07917_);
  or _19490_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _11139_, _11121_);
  and _19491_ (_11140_, _07917_, word_in[19]);
  and _19492_ (_11141_, _10590_, _07650_);
  and _19493_ (_11142_, _10604_, _07640_);
  or _19494_ (_11143_, _11142_, _11141_);
  and _19495_ (_11144_, _10598_, _07643_);
  and _19496_ (_11145_, _10594_, _07666_);
  or _19497_ (_11146_, _11145_, _11144_);
  or _19498_ (_11147_, _11146_, _11143_);
  or _19499_ (_11148_, _11147_, _07888_);
  and _19500_ (_11149_, _10567_, _07650_);
  and _19501_ (_11150_, _10584_, _07640_);
  or _19502_ (_11151_, _11150_, _11149_);
  and _19503_ (_11152_, _10572_, _07643_);
  and _19504_ (_11153_, _10577_, _07666_);
  or _19505_ (_11154_, _11153_, _11152_);
  or _19506_ (_11155_, _11154_, _11151_);
  or _19507_ (_11156_, _11155_, _07927_);
  nand _19508_ (_11157_, _11156_, _11148_);
  nor _19509_ (_11158_, _11157_, _07917_);
  or _19510_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _11158_, _11140_);
  and _19511_ (_11159_, _07917_, word_in[20]);
  and _19512_ (_11160_, _10643_, _07643_);
  and _19513_ (_11162_, _10634_, _07650_);
  or _19514_ (_11164_, _11162_, _11160_);
  and _19515_ (_11165_, _10650_, _07640_);
  and _19516_ (_11167_, _10638_, _07666_);
  or _19517_ (_11168_, _11167_, _11165_);
  or _19518_ (_11169_, _11168_, _11164_);
  or _19519_ (_11170_, _11169_, _07888_);
  and _19520_ (_11171_, _10614_, _07650_);
  and _19521_ (_11172_, _10628_, _07640_);
  or _19522_ (_11173_, _11172_, _11171_);
  and _19523_ (_11174_, _10622_, _07643_);
  and _19524_ (_11175_, _10618_, _07666_);
  or _19525_ (_11176_, _11175_, _11174_);
  or _19526_ (_11177_, _11176_, _11173_);
  or _19527_ (_11178_, _11177_, _07927_);
  nand _19528_ (_11179_, _11178_, _11170_);
  nor _19529_ (_11181_, _11179_, _07917_);
  or _19530_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _11181_, _11159_);
  and _19531_ (_11182_, _07917_, word_in[21]);
  and _19532_ (_11183_, _10688_, _07643_);
  and _19533_ (_11184_, _10684_, _07650_);
  or _19534_ (_11185_, _11184_, _11183_);
  and _19535_ (_11186_, _10694_, _07640_);
  and _19536_ (_11187_, _10680_, _07666_);
  or _19537_ (_11188_, _11187_, _11186_);
  or _19538_ (_11189_, _11188_, _11185_);
  or _19539_ (_11190_, _11189_, _07888_);
  and _19540_ (_11191_, _10664_, _07643_);
  and _19541_ (_11192_, _10668_, _07650_);
  or _19542_ (_11193_, _11192_, _11191_);
  and _19543_ (_11194_, _10674_, _07640_);
  and _19544_ (_11195_, _10660_, _07666_);
  or _19545_ (_11196_, _11195_, _11194_);
  or _19546_ (_11197_, _11196_, _11193_);
  or _19547_ (_11198_, _11197_, _07927_);
  nand _19548_ (_11199_, _11198_, _11190_);
  nor _19549_ (_11200_, _11199_, _07917_);
  or _19550_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11200_, _11182_);
  and _19551_ (_11201_, _07917_, word_in[22]);
  and _19552_ (_11202_, _10734_, _07643_);
  and _19553_ (_11203_, _10730_, _07650_);
  or _19554_ (_11204_, _11203_, _11202_);
  and _19555_ (_11205_, _10740_, _07640_);
  and _19556_ (_11206_, _10726_, _07666_);
  or _19557_ (_11207_, _11206_, _11205_);
  or _19558_ (_11208_, _11207_, _11204_);
  or _19559_ (_11209_, _11208_, _07888_);
  and _19560_ (_11210_, _10712_, _07650_);
  and _19561_ (_11211_, _10720_, _07640_);
  or _19562_ (_11212_, _11211_, _11210_);
  and _19563_ (_11213_, _10708_, _07643_);
  and _19564_ (_11215_, _10704_, _07666_);
  or _19565_ (_11216_, _11215_, _11213_);
  or _19566_ (_11218_, _11216_, _11212_);
  or _19567_ (_11219_, _11218_, _07927_);
  nand _19568_ (_11220_, _11219_, _11209_);
  nor _19569_ (_11222_, _11220_, _07917_);
  or _19570_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11222_, _11201_);
  and _19571_ (_11223_, _07984_, word_in[24]);
  and _19572_ (_11224_, _10766_, _07821_);
  and _19573_ (_11225_, _10762_, _07820_);
  or _19574_ (_11226_, _11225_, _11224_);
  and _19575_ (_11227_, _11226_, _07949_);
  and _19576_ (_11228_, _10756_, _07821_);
  and _19577_ (_11230_, _10752_, _07820_);
  or _19578_ (_11231_, _11230_, _11228_);
  and _19579_ (_11232_, _11231_, _07947_);
  and _19580_ (_11233_, _10776_, _07821_);
  and _19581_ (_11234_, _10772_, _07820_);
  or _19582_ (_11235_, _11234_, _11233_);
  and _19583_ (_11237_, _11235_, _07993_);
  and _19584_ (_11238_, _10786_, _07821_);
  and _19585_ (_11240_, _10782_, _07820_);
  or _19586_ (_11241_, _11240_, _11238_);
  and _19587_ (_11242_, _11241_, _08001_);
  or _19588_ (_11243_, _11242_, _11237_);
  or _19589_ (_11244_, _11243_, _11232_);
  nor _19590_ (_11245_, _11244_, _11227_);
  nor _19591_ (_11246_, _11245_, _07984_);
  or _19592_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11246_, _11223_);
  and _19593_ (_11247_, _07984_, word_in[25]);
  and _19594_ (_11248_, _10813_, _07821_);
  and _19595_ (_11249_, _10809_, _07820_);
  or _19596_ (_11250_, _11249_, _11248_);
  and _19597_ (_11251_, _11250_, _07949_);
  and _19598_ (_11252_, _10803_, _07821_);
  and _19599_ (_11253_, _10798_, _07820_);
  or _19600_ (_11255_, _11253_, _11252_);
  and _19601_ (_11256_, _11255_, _07947_);
  and _19602_ (_11257_, _10823_, _07821_);
  and _19603_ (_11258_, _10819_, _07820_);
  or _19604_ (_11260_, _11258_, _11257_);
  and _19605_ (_11261_, _11260_, _07993_);
  and _19606_ (_11262_, _10833_, _07821_);
  and _19607_ (_11264_, _10829_, _07820_);
  or _19608_ (_11265_, _11264_, _11262_);
  and _19609_ (_11266_, _11265_, _08001_);
  or _19610_ (_11267_, _11266_, _11261_);
  or _19611_ (_11268_, _11267_, _11256_);
  nor _19612_ (_11269_, _11268_, _11251_);
  nor _19613_ (_11270_, _11269_, _07984_);
  or _19614_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _11270_, _11247_);
  and _19615_ (_11271_, _07984_, word_in[26]);
  and _19616_ (_11272_, _10848_, _07821_);
  and _19617_ (_11273_, _10844_, _07820_);
  or _19618_ (_11274_, _11273_, _11272_);
  and _19619_ (_11275_, _11274_, _07947_);
  and _19620_ (_11276_, _10858_, _07821_);
  and _19621_ (_11277_, _10854_, _07820_);
  or _19622_ (_11278_, _11277_, _11276_);
  and _19623_ (_11279_, _11278_, _07949_);
  and _19624_ (_11280_, _10868_, _07821_);
  and _19625_ (_11282_, _10864_, _07820_);
  or _19626_ (_11283_, _11282_, _11280_);
  and _19627_ (_11284_, _11283_, _07993_);
  and _19628_ (_11285_, _10879_, _07821_);
  and _19629_ (_11286_, _10875_, _07820_);
  or _19630_ (_11287_, _11286_, _11285_);
  and _19631_ (_11288_, _11287_, _08001_);
  or _19632_ (_11289_, _11288_, _11284_);
  or _19633_ (_11290_, _11289_, _11279_);
  nor _19634_ (_11291_, _11290_, _11275_);
  nor _19635_ (_11292_, _11291_, _07984_);
  or _19636_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _11292_, _11271_);
  and _19637_ (_11293_, _07984_, word_in[27]);
  and _19638_ (_11294_, _10906_, _07821_);
  and _19639_ (_11295_, _10902_, _07820_);
  or _19640_ (_11296_, _11295_, _11294_);
  and _19641_ (_11297_, _11296_, _07949_);
  and _19642_ (_11298_, _10896_, _07821_);
  and _19643_ (_11299_, _10892_, _07820_);
  or _19644_ (_11301_, _11299_, _11298_);
  and _19645_ (_11302_, _11301_, _07947_);
  and _19646_ (_11303_, _10916_, _07821_);
  and _19647_ (_11304_, _10912_, _07820_);
  or _19648_ (_11305_, _11304_, _11303_);
  and _19649_ (_11306_, _11305_, _07993_);
  and _19650_ (_11307_, _10926_, _07821_);
  and _19651_ (_11308_, _10922_, _07820_);
  or _19652_ (_11309_, _11308_, _11307_);
  and _19653_ (_11311_, _11309_, _08001_);
  or _19654_ (_11312_, _11311_, _11306_);
  or _19655_ (_11313_, _11312_, _11302_);
  nor _19656_ (_11314_, _11313_, _11297_);
  nor _19657_ (_11315_, _11314_, _07984_);
  or _19658_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _11315_, _11293_);
  and _19659_ (_11316_, _07984_, word_in[28]);
  and _19660_ (_11317_, _10954_, _07821_);
  and _19661_ (_11318_, _10950_, _07820_);
  or _19662_ (_11320_, _11318_, _11317_);
  and _19663_ (_11321_, _11320_, _07949_);
  and _19664_ (_11322_, _10944_, _07821_);
  and _19665_ (_11324_, _10938_, _07820_);
  or _19666_ (_11325_, _11324_, _11322_);
  and _19667_ (_11326_, _11325_, _07947_);
  and _19668_ (_11327_, _10964_, _07821_);
  and _19669_ (_11328_, _10960_, _07820_);
  or _19670_ (_11329_, _11328_, _11327_);
  and _19671_ (_11330_, _11329_, _07993_);
  and _19672_ (_11331_, _10974_, _07821_);
  and _19673_ (_11332_, _10970_, _07820_);
  or _19674_ (_11333_, _11332_, _11331_);
  and _19675_ (_11334_, _11333_, _08001_);
  or _19676_ (_11336_, _11334_, _11330_);
  or _19677_ (_11337_, _11336_, _11326_);
  nor _19678_ (_11338_, _11337_, _11321_);
  nor _19679_ (_11339_, _11338_, _07984_);
  or _19680_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _11339_, _11316_);
  and _19681_ (_11340_, _07984_, word_in[29]);
  and _19682_ (_11341_, _11000_, _07821_);
  and _19683_ (_11342_, _10996_, _07820_);
  or _19684_ (_11343_, _11342_, _11341_);
  and _19685_ (_11344_, _11343_, _07949_);
  and _19686_ (_11345_, _10990_, _07821_);
  and _19687_ (_11347_, _10985_, _07820_);
  or _19688_ (_11348_, _11347_, _11345_);
  and _19689_ (_11349_, _11348_, _07947_);
  and _19690_ (_11350_, _11010_, _07821_);
  and _19691_ (_11351_, _11006_, _07820_);
  or _19692_ (_11352_, _11351_, _11350_);
  and _19693_ (_11353_, _11352_, _07993_);
  and _19694_ (_11354_, _11020_, _07821_);
  and _19695_ (_11355_, _11016_, _07820_);
  or _19696_ (_11357_, _11355_, _11354_);
  and _19697_ (_11358_, _11357_, _08001_);
  or _19698_ (_11359_, _11358_, _11353_);
  or _19699_ (_11361_, _11359_, _11349_);
  nor _19700_ (_11362_, _11361_, _11344_);
  nor _19701_ (_11364_, _11362_, _07984_);
  or _19702_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _11364_, _11340_);
  and _19703_ (_11365_, _07984_, word_in[30]);
  and _19704_ (_11366_, _11037_, _07821_);
  and _19705_ (_11367_, _11032_, _07820_);
  or _19706_ (_11368_, _11367_, _11366_);
  and _19707_ (_11369_, _11368_, _07947_);
  and _19708_ (_11370_, _11047_, _07821_);
  and _19709_ (_11371_, _11043_, _07820_);
  or _19710_ (_11372_, _11371_, _11370_);
  and _19711_ (_11373_, _11372_, _07949_);
  and _19712_ (_11374_, _11057_, _07821_);
  and _19713_ (_11375_, _11053_, _07820_);
  or _19714_ (_11377_, _11375_, _11374_);
  and _19715_ (_11378_, _11377_, _07993_);
  and _19716_ (_11379_, _11069_, _07821_);
  and _19717_ (_11380_, _11064_, _07820_);
  or _19718_ (_11381_, _11380_, _11379_);
  and _19719_ (_11382_, _11381_, _08001_);
  or _19720_ (_11383_, _11382_, _11378_);
  or _19721_ (_11384_, _11383_, _11373_);
  nor _19722_ (_11385_, _11384_, _11369_);
  nor _19723_ (_11386_, _11385_, _07984_);
  or _19724_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _11386_, _11365_);
  nand _19725_ (_11387_, _06415_, _06270_);
  or _19726_ (_11388_, _06270_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _19727_ (_11390_, _11388_, _05141_);
  and _19728_ (_09833_, _11390_, _11387_);
  or _19729_ (_11391_, _06497_, _07117_);
  or _19730_ (_11392_, _06270_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _19731_ (_11393_, _11392_, _05141_);
  and _19732_ (_09855_, _11393_, _11391_);
  or _19733_ (_11394_, _06447_, _07117_);
  or _19734_ (_11395_, _06270_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _19735_ (_11396_, _11395_, _05141_);
  and _19736_ (_09859_, _11396_, _11394_);
  or _19737_ (_11397_, _06524_, _07117_);
  or _19738_ (_11398_, _06270_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _19739_ (_11399_, _11398_, _05141_);
  and _19740_ (_09862_, _11399_, _11397_);
  and _19741_ (_11400_, _08382_, _06004_);
  and _19742_ (_11401_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _19743_ (_11402_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _19744_ (_11403_, _11402_, _11401_);
  nor _19745_ (_11404_, _11403_, _08243_);
  and _19746_ (_11405_, _08396_, _05522_);
  or _19747_ (_11406_, _11405_, _11404_);
  or _19748_ (_11407_, _11406_, _11400_);
  and _19749_ (_10068_, _11407_, _05141_);
  nor _19750_ (_11408_, _08656_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _19751_ (_11410_, _11408_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _19752_ (_11411_, _11408_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _19753_ (_11412_, _11411_, _05141_);
  and _19754_ (_10072_, _11412_, _11410_);
  nand _19755_ (_11413_, _07350_, _06624_);
  or _19756_ (_11414_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _19757_ (_11415_, _11414_, _05141_);
  and _19758_ (_10236_, _11415_, _11413_);
  nor _19759_ (_11417_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _19760_ (_11418_, _11417_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _19761_ (_03037_, _11418_, _05141_);
  and _19762_ (_10494_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _05141_);
  and _19763_ (_11419_, _10494_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _19764_ (_10245_, _11419_, _03037_);
  not _19765_ (_11420_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _19766_ (_11421_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , _11420_);
  and _19767_ (_10251_, _11421_, _05141_);
  and _19768_ (_11422_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _19769_ (_11423_, _11422_);
  nand _19770_ (_11424_, _08344_, _05143_);
  and _19771_ (_11425_, _11424_, _11423_);
  and _19772_ (_11426_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _19773_ (_11427_, _11426_);
  or _19774_ (_11428_, _06564_, _06556_);
  and _19775_ (_11429_, _11428_, _06771_);
  and _19776_ (_11430_, _06771_, _06563_);
  and _19777_ (_11431_, _11430_, _06450_);
  nor _19778_ (_11432_, _11431_, _11429_);
  or _19779_ (_11433_, _07053_, _06529_);
  nand _19780_ (_11434_, _11433_, _06771_);
  nand _19781_ (_11435_, _07044_, _06449_);
  and _19782_ (_11436_, _11435_, _11434_);
  and _19783_ (_11437_, _11436_, _11432_);
  nand _19784_ (_11438_, _06556_, _06544_);
  not _19785_ (_11439_, _11438_);
  nor _19786_ (_11440_, _11439_, _07076_);
  and _19787_ (_11441_, _07069_, _06766_);
  nor _19788_ (_11442_, _11441_, _06772_);
  and _19789_ (_11443_, _06771_, _06765_);
  nor _19790_ (_11444_, _11443_, _06979_);
  and _19791_ (_11445_, _11444_, _11442_);
  and _19792_ (_11446_, _11445_, _11440_);
  and _19793_ (_11447_, _11446_, _11437_);
  nand _19794_ (_11448_, _11447_, _08337_);
  nand _19795_ (_11449_, _11448_, _06821_);
  and _19796_ (_11450_, _11439_, _07087_);
  and _19797_ (_11451_, _11450_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _19798_ (_11452_, _07088_, _06575_);
  nor _19799_ (_11453_, _11452_, _11451_);
  nand _19800_ (_11454_, _11453_, _11449_);
  nand _19801_ (_11455_, _11454_, _05143_);
  nand _19802_ (_11456_, _11455_, _11427_);
  and _19803_ (_11457_, _11456_, _11425_);
  and _19804_ (_10319_, _11457_, _05141_);
  and _19805_ (_10340_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _05141_);
  and _19806_ (_11458_, _10343_, _06204_);
  and _19807_ (_11459_, _11458_, _05288_);
  nand _19808_ (_11460_, _11459_, _05963_);
  or _19809_ (_11461_, _11459_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _19810_ (_11462_, _06734_, _05926_);
  not _19811_ (_11463_, _11462_);
  and _19812_ (_11464_, _11463_, _11461_);
  and _19813_ (_11465_, _11464_, _11460_);
  nor _19814_ (_11466_, _11463_, _06178_);
  or _19815_ (_11467_, _11466_, _11465_);
  and _19816_ (_10344_, _11467_, _05141_);
  and _19817_ (_11468_, _11458_, _05210_);
  and _19818_ (_11469_, _11468_, _05963_);
  nor _19819_ (_11470_, _11468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _19820_ (_11471_, _11470_, _11469_);
  nand _19821_ (_11472_, _11471_, _11463_);
  nand _19822_ (_11473_, _11462_, _05604_);
  and _19823_ (_11474_, _11473_, _05141_);
  and _19824_ (_10347_, _11474_, _11472_);
  nor _19825_ (_11475_, _07619_, _07516_);
  nor _19826_ (_11476_, _06363_, _06337_);
  and _19827_ (_11477_, _11476_, _07010_);
  not _19828_ (_11478_, _11477_);
  and _19829_ (_11479_, _06497_, _07023_);
  and _19830_ (_11480_, _11479_, _07007_);
  and _19831_ (_11481_, _06524_, _07006_);
  and _19832_ (_11482_, _11481_, _07014_);
  nor _19833_ (_11483_, _11482_, _11480_);
  nor _19834_ (_11484_, _11483_, _11478_);
  not _19835_ (_11485_, _11484_);
  and _19836_ (_11486_, _06497_, _06447_);
  nor _19837_ (_11487_, _06497_, _06447_);
  nor _19838_ (_11488_, _11487_, _11486_);
  and _19839_ (_11489_, _11488_, _07007_);
  and _19840_ (_11490_, _11489_, _07018_);
  not _19841_ (_11491_, _07021_);
  and _19842_ (_11492_, _06524_, _06472_);
  and _19843_ (_11493_, _11492_, _11479_);
  and _19844_ (_11494_, _07006_, _06447_);
  and _19845_ (_11495_, _11494_, _07007_);
  nor _19846_ (_11496_, _11495_, _11493_);
  nor _19847_ (_11497_, _11496_, _11491_);
  nor _19848_ (_11498_, _11497_, _11490_);
  and _19849_ (_11499_, _11498_, _11485_);
  and _19850_ (_11500_, _11494_, _11492_);
  and _19851_ (_11501_, _11500_, _11477_);
  not _19852_ (_11502_, _11501_);
  nor _19853_ (_11503_, _07017_, _06337_);
  and _19854_ (_11504_, _11503_, _07010_);
  and _19855_ (_11505_, _07023_, _06415_);
  and _19856_ (_11506_, _06389_, _06337_);
  and _19857_ (_11507_, _11506_, _11505_);
  and _19858_ (_11508_, _11507_, _07007_);
  nor _19859_ (_11509_, _11508_, _11504_);
  and _19860_ (_11510_, _11509_, _11502_);
  and _19861_ (_11511_, _11492_, _11486_);
  and _19862_ (_11512_, _11511_, _07022_);
  and _19863_ (_11513_, _11493_, _07011_);
  nor _19864_ (_11514_, _11513_, _11512_);
  and _19865_ (_11516_, _11514_, _11510_);
  and _19866_ (_11517_, _06524_, _07014_);
  and _19867_ (_11518_, _11517_, _11479_);
  and _19868_ (_11519_, _07021_, _06363_);
  and _19869_ (_11520_, _11519_, _11518_);
  not _19870_ (_11521_, _11519_);
  and _19871_ (_11522_, _11517_, _11487_);
  nor _19872_ (_11524_, _11522_, _07015_);
  nor _19873_ (_11525_, _11524_, _11521_);
  nor _19874_ (_11527_, _11525_, _11520_);
  and _19875_ (_11528_, _11527_, _11516_);
  and _19876_ (_11529_, _11528_, _11499_);
  nor _19877_ (_11530_, _07021_, _07018_);
  and _19878_ (_11531_, _11492_, _11487_);
  and _19879_ (_11532_, _11517_, _11486_);
  and _19880_ (_11533_, _11519_, _11532_);
  nor _19881_ (_11534_, _11533_, _11531_);
  nor _19882_ (_11535_, _11534_, _11530_);
  not _19883_ (_11536_, _11535_);
  and _19884_ (_11537_, _07015_, _07006_);
  and _19885_ (_11538_, _11537_, _07018_);
  not _19886_ (_11539_, _11538_);
  and _19887_ (_11540_, _11477_, _07015_);
  nand _19888_ (_11541_, _11540_, _11488_);
  not _19889_ (_11542_, _11541_);
  and _19890_ (_11543_, _11517_, _11494_);
  and _19891_ (_11544_, _11543_, _11519_);
  nor _19892_ (_11545_, _11544_, _11542_);
  and _19893_ (_11546_, _11545_, _11539_);
  and _19894_ (_11547_, _11486_, _07007_);
  and _19895_ (_11548_, _11547_, _07022_);
  and _19896_ (_11549_, _11487_, _07007_);
  nor _19897_ (_11550_, _11511_, _11549_);
  nor _19898_ (_11551_, _11550_, _11521_);
  nor _19899_ (_11552_, _11551_, _11548_);
  and _19900_ (_11553_, _11552_, _11546_);
  and _19901_ (_11554_, _11553_, _11536_);
  and _19902_ (_11555_, _11554_, _11529_);
  and _19903_ (_11556_, _07007_, _06497_);
  not _19904_ (_11557_, _11556_);
  nor _19905_ (_11558_, _11543_, _11511_);
  and _19906_ (_11559_, _11558_, _11557_);
  nor _19907_ (_11560_, _11559_, _06415_);
  not _19908_ (_11561_, _11500_);
  nor _19909_ (_11562_, _11530_, _11561_);
  nor _19910_ (_11563_, _11562_, _11560_);
  and _19911_ (_11564_, _11547_, _11519_);
  and _19912_ (_11565_, _11500_, _07012_);
  nor _19913_ (_11566_, _11565_, _11564_);
  not _19914_ (_11567_, _11566_);
  not _19915_ (_11568_, _07018_);
  nor _19916_ (_11569_, _11522_, _11547_);
  and _19917_ (_11570_, _11569_, _11558_);
  nor _19918_ (_11571_, _11570_, _11568_);
  nor _19919_ (_11572_, _11571_, _11567_);
  and _19920_ (_11573_, _11572_, _11563_);
  not _19921_ (_11574_, _11549_);
  nor _19922_ (_11575_, _11477_, _07009_);
  and _19923_ (_11576_, _11575_, _11568_);
  or _19924_ (_11577_, _11576_, _11574_);
  and _19925_ (_11578_, _06447_, _06415_);
  and _19926_ (_11579_, _11506_, _11578_);
  and _19927_ (_11580_, _11492_, _06497_);
  or _19928_ (_11581_, _11556_, _11580_);
  and _19929_ (_11582_, _11581_, _11579_);
  not _19930_ (_11583_, _11582_);
  nand _19931_ (_11584_, _11580_, _11477_);
  not _19932_ (_11585_, _11584_);
  and _19933_ (_11586_, _07022_, _07016_);
  nor _19934_ (_11587_, _11586_, _11585_);
  and _19935_ (_11588_, _11587_, _11583_);
  and _19936_ (_11589_, _11588_, _11577_);
  and _19937_ (_11590_, _11531_, _07012_);
  and _19938_ (_11591_, _11495_, _11477_);
  nor _19939_ (_11592_, _11591_, _11590_);
  not _19940_ (_11593_, _11592_);
  not _19941_ (_11594_, _11547_);
  and _19942_ (_11595_, _11486_, _07015_);
  nor _19943_ (_11596_, _11531_, _11595_);
  and _19944_ (_11597_, _11596_, _11594_);
  nor _19945_ (_11598_, _11597_, _11478_);
  nor _19946_ (_11599_, _11598_, _11593_);
  and _19947_ (_11600_, _11599_, _11589_);
  and _19948_ (_11601_, _11600_, _11573_);
  and _19949_ (_11602_, _11601_, _11555_);
  nor _19950_ (_11603_, _11602_, _06318_);
  not _19951_ (_11604_, _11602_);
  and _19952_ (_11605_, _11513_, _06363_);
  not _19953_ (_11606_, _11605_);
  and _19954_ (_11607_, _11477_, _11595_);
  or _19955_ (_11608_, _11506_, _07009_);
  and _19956_ (_11609_, _11608_, _11547_);
  nor _19957_ (_11610_, _11609_, _11607_);
  and _19958_ (_11611_, _11610_, _11606_);
  and _19959_ (_11612_, _11611_, _11592_);
  and _19960_ (_11613_, _11612_, _11566_);
  and _19961_ (_11614_, _11613_, _11553_);
  nand _19962_ (_11615_, _11614_, _11604_);
  and _19963_ (_11617_, _11615_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _19964_ (_11618_, _11602_, _06318_);
  nor _19965_ (_11619_, _11618_, _11603_);
  and _19966_ (_11620_, _11619_, _11617_);
  nor _19967_ (_11621_, _11620_, _11603_);
  nor _19968_ (_11622_, _11621_, _07516_);
  and _19969_ (_11623_, _11622_, _06302_);
  nor _19970_ (_11624_, _11622_, _06302_);
  nor _19971_ (_11625_, _11624_, _11623_);
  nor _19972_ (_11626_, _11625_, _11475_);
  and _19973_ (_11627_, _06319_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _19974_ (_11628_, _11627_, _11475_);
  nor _19975_ (_11629_, _11628_, _11614_);
  or _19976_ (_11630_, _11629_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _19977_ (_11631_, _11630_, _11626_);
  and _19978_ (_10377_, _11631_, _05141_);
  and _19979_ (_11633_, _05141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  not _19980_ (_11634_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor _19981_ (_11635_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _19982_ (_11636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _19983_ (_11637_, _11636_, _11635_);
  not _19984_ (_11639_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _19985_ (_11640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _19986_ (_11642_, _11640_, _11639_);
  and _19987_ (_11643_, _11642_, _11637_);
  and _19988_ (_11644_, _11643_, _11634_);
  and _19989_ (_11646_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _05141_);
  and _19990_ (_11647_, _11646_, _11644_);
  or _19991_ (_10382_, _11647_, _11633_);
  nor _19992_ (_11648_, _11644_, rst);
  or _19993_ (_11649_, _07516_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _19994_ (_11650_, _11649_, _10340_);
  or _19995_ (_10388_, _11650_, _11648_);
  not _19996_ (_11651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _19997_ (_11652_, _06725_, _11651_);
  or _19998_ (_11653_, _11652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _19999_ (_11654_, _11653_, _11458_);
  not _20000_ (_11655_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _20001_ (_11656_, _06207_, _11655_);
  nand _20002_ (_11657_, _11656_, _11458_);
  or _20003_ (_11659_, _11657_, _06208_);
  and _20004_ (_11660_, _11659_, _11654_);
  or _20005_ (_11661_, _11660_, _11462_);
  nand _20006_ (_11662_, _11462_, _06244_);
  and _20007_ (_11663_, _11662_, _05141_);
  and _20008_ (_10406_, _11663_, _11661_);
  and _20009_ (_11665_, _05922_, _10407_);
  or _20010_ (_11667_, _05209_, _05186_);
  nor _20011_ (_11668_, _05287_, _08651_);
  and _20012_ (_11669_, _11668_, _11667_);
  or _20013_ (_11671_, _11669_, _11665_);
  and _20014_ (_11672_, _11671_, _11458_);
  nor _20015_ (_11673_, _06209_, _05287_);
  nand _20016_ (_11674_, _11458_, _11673_);
  and _20017_ (_11676_, _11674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _20018_ (_11678_, _11676_, _11462_);
  or _20019_ (_11680_, _11678_, _11672_);
  or _20020_ (_11681_, _11463_, _06004_);
  and _20021_ (_11683_, _11681_, _05141_);
  and _20022_ (_10409_, _11683_, _11680_);
  and _20023_ (_11684_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _20024_ (_11685_, _11684_, _10380_);
  and _20025_ (_11686_, _11685_, _11458_);
  not _20026_ (_11687_, _11458_);
  or _20027_ (_11689_, _11687_, _10375_);
  and _20028_ (_11690_, _11689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _20029_ (_11691_, _11690_, _11462_);
  or _20030_ (_11692_, _11691_, _11686_);
  or _20031_ (_11693_, _11463_, _05522_);
  and _20032_ (_11694_, _11693_, _05141_);
  and _20033_ (_10412_, _11694_, _11692_);
  and _20034_ (_11696_, _08283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _20035_ (_11698_, _11696_, _08281_);
  and _20036_ (_11699_, _11698_, _11458_);
  nand _20037_ (_11701_, _11458_, _05186_);
  and _20038_ (_11702_, _11701_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _20039_ (_11704_, _11702_, _11462_);
  or _20040_ (_11705_, _11704_, _11699_);
  nand _20041_ (_11706_, _11462_, _06062_);
  and _20042_ (_11707_, _11706_, _05141_);
  and _20043_ (_10417_, _11707_, _11705_);
  and _20044_ (_11708_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _20045_ (_11709_, _11708_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  or _20046_ (_11710_, _11709_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _20047_ (_10458_, _11710_, _05141_);
  not _20048_ (_11711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand _20049_ (_11712_, _08463_, _11711_);
  nor _20050_ (_11713_, _06727_, _11711_);
  and _20051_ (_11714_, _11713_, _08439_);
  and _20052_ (_11715_, _11714_, _08457_);
  and _20053_ (_11716_, _08453_, _08439_);
  and _20054_ (_11718_, _11716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor _20055_ (_11720_, _11716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor _20056_ (_11721_, _11720_, _11718_);
  or _20057_ (_11722_, _11721_, _08463_);
  or _20058_ (_11723_, _11722_, _11715_);
  and _20059_ (_11724_, _11723_, _11712_);
  and _20060_ (_11725_, _06736_, _10407_);
  and _20061_ (_11726_, _11725_, _06734_);
  nor _20062_ (_11727_, _11726_, _08471_);
  and _20063_ (_11728_, _11727_, _11724_);
  and _20064_ (_11729_, _08478_, _06703_);
  and _20065_ (_11730_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _20066_ (_11731_, _11730_, _11729_);
  or _20067_ (_11732_, _11731_, _11728_);
  and _20068_ (_10461_, _11732_, _05141_);
  not _20069_ (_11733_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _20070_ (_11734_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor _20071_ (_11735_, _11734_, _11733_);
  and _20072_ (_11736_, _11734_, _11733_);
  nor _20073_ (_11737_, _11736_, _11735_);
  not _20074_ (_11738_, _11737_);
  and _20075_ (_11739_, _11738_, _10458_);
  nor _20076_ (_11740_, _11735_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _20077_ (_11741_, _11735_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _20078_ (_11742_, _11741_, _11740_);
  nor _20079_ (_11743_, _11708_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _20080_ (_11744_, _11743_, _11709_);
  or _20081_ (_11745_, _11744_, _11734_);
  and _20082_ (_11746_, _11745_, _11742_);
  and _20083_ (_10476_, _11746_, _11739_);
  nor _20084_ (_11747_, _08478_, _08471_);
  and _20085_ (_11748_, _11718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _20086_ (_11749_, _11748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand _20087_ (_11750_, _11749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _20088_ (_11751_, _11749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _20089_ (_11752_, _11751_, _11750_);
  not _20090_ (_11753_, _06727_);
  and _20091_ (_11754_, _08439_, _11753_);
  and _20092_ (_11755_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _20093_ (_11756_, _11755_, _08457_);
  or _20094_ (_11757_, _11756_, _08463_);
  or _20095_ (_11758_, _11757_, _11752_);
  or _20096_ (_11759_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _20097_ (_11760_, _11759_, _11758_);
  and _20098_ (_11761_, _11760_, _11747_);
  nor _20099_ (_11762_, _08479_, _06062_);
  and _20100_ (_11763_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _20101_ (_11764_, _11763_, _11762_);
  or _20102_ (_11765_, _11764_, _11761_);
  and _20103_ (_10489_, _11765_, _05141_);
  nor _20104_ (_11766_, _11748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _20105_ (_11767_, _11766_, _11749_);
  or _20106_ (_11768_, _11767_, _08463_);
  and _20107_ (_11769_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _20108_ (_11770_, _11769_, _08457_);
  or _20109_ (_11771_, _11770_, _11768_);
  or _20110_ (_11772_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _20111_ (_11773_, _11772_, _11771_);
  and _20112_ (_11774_, _11773_, _11747_);
  and _20113_ (_11775_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _20114_ (_11776_, _11775_, _11774_);
  nor _20115_ (_11777_, _08479_, _05560_);
  or _20116_ (_11778_, _11777_, _11776_);
  and _20117_ (_10492_, _11778_, _05141_);
  and _20118_ (_11779_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _20119_ (_11780_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _20120_ (_11781_, _11718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _20121_ (_11782_, _11781_, _11748_);
  or _20122_ (_11783_, _11782_, _08463_);
  and _20123_ (_11784_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _20124_ (_11785_, _11784_, _08457_);
  or _20125_ (_11786_, _11785_, _11783_);
  and _20126_ (_11787_, _11786_, _11780_);
  and _20127_ (_11788_, _11787_, _11727_);
  not _20128_ (_11789_, _11726_);
  nor _20129_ (_11790_, _11789_, _06178_);
  or _20130_ (_11791_, _11790_, _11788_);
  or _20131_ (_11792_, _11791_, _11779_);
  and _20132_ (_10499_, _11792_, _05141_);
  and _20133_ (_11793_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07611_);
  and _20134_ (_11794_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _20135_ (_11795_, _11794_, _11793_);
  and _20136_ (_10503_, _11795_, _05141_);
  and _20137_ (_11796_, _06520_, _06468_);
  and _20138_ (_11797_, _11796_, _06442_);
  and _20139_ (_11798_, _06269_, _06317_);
  and _20140_ (_11799_, _11798_, _06296_);
  and _20141_ (_11800_, _11799_, _06332_);
  and _20142_ (_11801_, _06493_, _06410_);
  and _20143_ (_11802_, _11801_, _11800_);
  and _20144_ (_11803_, _06385_, _06358_);
  and _20145_ (_11804_, _11803_, _11802_);
  and _20146_ (_10510_, _11804_, _11797_);
  and _20147_ (_11805_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _20148_ (_11806_, _08478_, _06004_);
  or _20149_ (_11807_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _20150_ (_11808_, _08453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _20151_ (_11809_, _11808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _20152_ (_11810_, _11809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _20153_ (_11811_, _11810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _20154_ (_11812_, _11811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _20155_ (_11813_, _11812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _20156_ (_11814_, _11813_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _20157_ (_11815_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _20158_ (_11816_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _20159_ (_11817_, _11816_, _11815_);
  and _20160_ (_11818_, _08455_, _08439_);
  or _20161_ (_11819_, _11818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand _20162_ (_11820_, _11818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _20163_ (_11821_, _11820_, _11819_);
  or _20164_ (_11822_, _11821_, _08463_);
  or _20165_ (_11823_, _11822_, _11817_);
  and _20166_ (_11824_, _11823_, _11807_);
  and _20167_ (_11825_, _11824_, _11747_);
  or _20168_ (_11826_, _11825_, _11806_);
  or _20169_ (_11827_, _11826_, _11805_);
  and _20170_ (_10529_, _11827_, _05141_);
  nand _20171_ (_11828_, _11726_, _06244_);
  and _20172_ (_11829_, _08456_, _08439_);
  and _20173_ (_11830_, _11829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _20174_ (_11831_, _11829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _20175_ (_11832_, _11831_, _11830_);
  and _20176_ (_11833_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _20177_ (_11834_, _11833_, _08439_);
  and _20178_ (_11835_, _11834_, _08457_);
  or _20179_ (_11836_, _11835_, _08463_);
  or _20180_ (_11837_, _11836_, _11832_);
  nor _20181_ (_11838_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _20182_ (_11839_, _11838_, _08471_);
  and _20183_ (_11840_, _11839_, _11837_);
  and _20184_ (_11841_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _20185_ (_11842_, _11841_, _08478_);
  or _20186_ (_11843_, _11842_, _11840_);
  and _20187_ (_11844_, _11843_, _05141_);
  and _20188_ (_10540_, _11844_, _11828_);
  not _20189_ (_11845_, _05522_);
  and _20190_ (_11846_, _05256_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _20191_ (_11847_, _10355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _20192_ (_11848_, _11847_, _10387_);
  and _20193_ (_11849_, _11848_, _10341_);
  nor _20194_ (_11850_, _11849_, _11846_);
  and _20195_ (_11851_, _06531_, _05197_);
  not _20196_ (_11852_, _11851_);
  and _20197_ (_11853_, _06365_, _05286_);
  nand _20198_ (_11854_, _05266_, _05287_);
  nor _20199_ (_11855_, _11854_, _11853_);
  and _20200_ (_11856_, _11855_, _11852_);
  and _20201_ (_11857_, _11856_, _05242_);
  and _20202_ (_11858_, _11857_, _05297_);
  nand _20203_ (_11859_, _10355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _20204_ (_11860_, _10355_, _06062_);
  nand _20205_ (_11861_, _11860_, _11859_);
  or _20206_ (_11862_, _11861_, _05172_);
  and _20207_ (_11863_, _11860_, _11859_);
  or _20208_ (_11864_, _11863_, _05173_);
  and _20209_ (_11865_, _11864_, _11862_);
  and _20210_ (_11866_, _11865_, _11858_);
  and _20211_ (_11867_, _11866_, _11850_);
  nand _20212_ (_11868_, _11867_, _05960_);
  not _20213_ (_11869_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or _20214_ (_11870_, _11847_, _10387_);
  and _20215_ (_11871_, _11863_, _06365_);
  nand _20216_ (_11872_, _11871_, _11870_);
  or _20217_ (_11873_, _11872_, _11869_);
  and _20218_ (_11874_, _11861_, _06365_);
  and _20219_ (_11875_, _11874_, _11848_);
  nand _20220_ (_11876_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _20221_ (_11877_, _11876_, _11873_);
  and _20222_ (_11878_, _11863_, _06531_);
  and _20223_ (_11879_, _11878_, _11870_);
  nand _20224_ (_11880_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _20225_ (_11881_, _11878_, _11848_);
  nand _20226_ (_11882_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _20227_ (_11883_, _11882_, _11880_);
  and _20228_ (_11884_, _11883_, _11877_);
  not _20229_ (_11885_, _11867_);
  and _20230_ (_11886_, _11861_, _06531_);
  and _20231_ (_11887_, _11886_, _11870_);
  nand _20232_ (_11888_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _20233_ (_11889_, _11874_, _11870_);
  nand _20234_ (_11891_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _20235_ (_11892_, _11891_, _11888_);
  and _20236_ (_11893_, _11886_, _11848_);
  nand _20237_ (_11894_, _11893_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _20238_ (_11895_, _11871_, _11848_);
  nand _20239_ (_11896_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _20240_ (_11897_, _11896_, _11894_);
  and _20241_ (_11898_, _11897_, _11892_);
  and _20242_ (_11899_, _11898_, _11885_);
  nand _20243_ (_11900_, _11899_, _11884_);
  and _20244_ (_11901_, _11900_, _11868_);
  and _20245_ (_10555_, _11901_, _05141_);
  and _20246_ (_10557_, _11870_, _05141_);
  not _20247_ (_11902_, _08471_);
  or _20248_ (_11903_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _20249_ (_11904_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _20250_ (_11905_, _11904_, _08439_);
  and _20251_ (_11906_, _11905_, _08457_);
  nand _20252_ (_11907_, _08448_, _08439_);
  nor _20253_ (_11908_, _11907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _20254_ (_11909_, _11907_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _20255_ (_11910_, _11909_, _08463_);
  or _20256_ (_11911_, _11910_, _11908_);
  or _20257_ (_11912_, _11911_, _11906_);
  nand _20258_ (_11913_, _11912_, _11903_);
  nand _20259_ (_11914_, _11913_, _11902_);
  nand _20260_ (_11915_, _08471_, _06062_);
  and _20261_ (_11916_, _11915_, _11914_);
  or _20262_ (_11917_, _11916_, _11726_);
  or _20263_ (_11918_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _20264_ (_11919_, _11918_, _05141_);
  and _20265_ (_10570_, _11919_, _11917_);
  nor _20266_ (_11920_, _11902_, _06244_);
  and _20267_ (_11922_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _20268_ (_11923_, _11922_, _08439_);
  and _20269_ (_11924_, _11923_, _08457_);
  nand _20270_ (_11925_, _08451_, _08439_);
  nor _20271_ (_11926_, _11925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _20272_ (_11927_, _11925_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _20273_ (_11928_, _11927_, _08463_);
  or _20274_ (_11929_, _11928_, _11926_);
  or _20275_ (_11930_, _11929_, _11924_);
  nor _20276_ (_11931_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _20277_ (_11932_, _11931_, _08471_);
  and _20278_ (_11933_, _11932_, _11930_);
  or _20279_ (_11934_, _11933_, _11726_);
  or _20280_ (_11935_, _11934_, _11920_);
  or _20281_ (_11936_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _20282_ (_11937_, _11936_, _05141_);
  and _20283_ (_10575_, _11937_, _11935_);
  and _20284_ (_11938_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _20285_ (_11939_, _11938_, _08439_);
  and _20286_ (_11940_, _11939_, _08457_);
  and _20287_ (_11941_, _08450_, _08439_);
  or _20288_ (_11942_, _11941_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _20289_ (_11943_, _11942_, _11925_);
  or _20290_ (_11944_, _11943_, _08463_);
  or _20291_ (_11945_, _11944_, _11940_);
  nor _20292_ (_11946_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor _20293_ (_11948_, _11946_, _08471_);
  and _20294_ (_11949_, _11948_, _11945_);
  and _20295_ (_11950_, _08471_, _06004_);
  or _20296_ (_11951_, _11950_, _08478_);
  or _20297_ (_11952_, _11951_, _11949_);
  or _20298_ (_11953_, _08479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _20299_ (_11954_, _11953_, _05141_);
  and _20300_ (_10583_, _11954_, _11952_);
  and _20301_ (_11955_, _05651_, _05209_);
  and _20302_ (_11956_, _11955_, _06734_);
  and _20303_ (_11957_, _11956_, _05925_);
  or _20304_ (_11958_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _20305_ (_11959_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _20306_ (_11960_, _11959_, _08439_);
  and _20307_ (_11961_, _11960_, _08457_);
  and _20308_ (_11962_, _08449_, _08439_);
  nor _20309_ (_11963_, _11962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _20310_ (_11964_, _11963_, _11941_);
  or _20311_ (_11965_, _11964_, _08463_);
  or _20312_ (_11966_, _11965_, _11961_);
  nand _20313_ (_11967_, _11966_, _11958_);
  nor _20314_ (_11969_, _11967_, _11957_);
  and _20315_ (_11970_, _11957_, _05522_);
  or _20316_ (_11971_, _11970_, _11969_);
  or _20317_ (_11972_, _11971_, _11726_);
  or _20318_ (_11973_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _20319_ (_11974_, _11973_, _05141_);
  and _20320_ (_10610_, _11974_, _11972_);
  and _20321_ (_11976_, _05141_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _20322_ (_11977_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _20323_ (_11978_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _20324_ (_11980_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _20325_ (_11981_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _20326_ (_11982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _20327_ (_11983_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _20328_ (_11984_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _20329_ (_11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _20330_ (_11986_, _11985_, _11983_);
  and _20331_ (_11988_, _11986_, _11984_);
  nor _20332_ (_11989_, _11988_, _11983_);
  nor _20333_ (_11990_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _20334_ (_11991_, _11990_, _11982_);
  not _20335_ (_11992_, _11991_);
  nor _20336_ (_11994_, _11992_, _11989_);
  nor _20337_ (_11996_, _11994_, _11982_);
  not _20338_ (_11997_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _20339_ (_11998_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _20340_ (_11999_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _20341_ (_12000_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _20342_ (_12001_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _20343_ (_12003_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _20344_ (_12004_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _20345_ (_12005_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _20346_ (_12006_, _12005_, _12004_);
  and _20347_ (_12007_, _12006_, _12003_);
  and _20348_ (_12009_, _12007_, _12001_);
  and _20349_ (_12010_, _12009_, _12000_);
  and _20350_ (_12011_, _12010_, _11999_);
  and _20351_ (_12012_, _12011_, _11998_);
  and _20352_ (_12014_, _12012_, _11997_);
  and _20353_ (_12015_, _12014_, _11996_);
  and _20354_ (_12017_, _12015_, _11981_);
  and _20355_ (_12019_, _12017_, _11980_);
  and _20356_ (_12020_, _12019_, _11978_);
  and _20357_ (_12021_, _12020_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _20358_ (_12022_, _12020_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _20359_ (_12023_, _12022_, _12021_);
  nor _20360_ (_12024_, _12019_, _11978_);
  nor _20361_ (_12025_, _12024_, _12020_);
  nor _20362_ (_12026_, _12017_, _11980_);
  nor _20363_ (_12027_, _12026_, _12019_);
  nor _20364_ (_12028_, _12015_, _11981_);
  nor _20365_ (_12029_, _12028_, _12017_);
  not _20366_ (_12030_, _12029_);
  and _20367_ (_12031_, _12012_, _11996_);
  nor _20368_ (_12032_, _12031_, _11997_);
  nor _20369_ (_12033_, _12032_, _12015_);
  not _20370_ (_12034_, _12033_);
  and _20371_ (_12035_, _12011_, _11996_);
  nor _20372_ (_12036_, _12035_, _11998_);
  nor _20373_ (_12037_, _12036_, _12031_);
  not _20374_ (_12038_, _12037_);
  and _20375_ (_12039_, _12010_, _11996_);
  nor _20376_ (_12040_, _12039_, _11999_);
  nor _20377_ (_12041_, _12040_, _12035_);
  not _20378_ (_12042_, _12041_);
  and _20379_ (_12043_, _11996_, _12009_);
  nor _20380_ (_12044_, _12043_, _12000_);
  nor _20381_ (_12045_, _12044_, _12039_);
  not _20382_ (_12046_, _12045_);
  and _20383_ (_12047_, _11996_, _12007_);
  nor _20384_ (_12048_, _12047_, _12001_);
  nor _20385_ (_12049_, _12048_, _12043_);
  not _20386_ (_12050_, _12049_);
  and _20387_ (_12051_, _11996_, _12006_);
  nor _20388_ (_12052_, _12051_, _12003_);
  or _20389_ (_12053_, _12052_, _12047_);
  not _20390_ (_12054_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  not _20391_ (_12055_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _20392_ (_12056_, _11996_, _12055_);
  and _20393_ (_12057_, _12056_, _12054_);
  nor _20394_ (_12059_, _12057_, _12004_);
  or _20395_ (_12060_, _12059_, _12051_);
  nor _20396_ (_12061_, _11996_, _12055_);
  nor _20397_ (_12062_, _12061_, _12056_);
  not _20398_ (_12063_, _12062_);
  nor _20399_ (_12064_, _11986_, _11984_);
  nor _20400_ (_12065_, _12064_, _11988_);
  nand _20401_ (_12066_, _12065_, _11604_);
  not _20402_ (_12068_, _12066_);
  nor _20403_ (_12069_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _20404_ (_12071_, _12069_, _11984_);
  and _20405_ (_12072_, _12071_, _11615_);
  or _20406_ (_12074_, _12065_, _11604_);
  and _20407_ (_12075_, _12074_, _12066_);
  and _20408_ (_12077_, _12075_, _12072_);
  or _20409_ (_12078_, _12077_, _12068_);
  and _20410_ (_12079_, _11992_, _11989_);
  nor _20411_ (_12081_, _12079_, _11994_);
  and _20412_ (_12083_, _12081_, _12078_);
  and _20413_ (_12084_, _12083_, _12063_);
  nor _20414_ (_12086_, _12056_, _12054_);
  or _20415_ (_12087_, _12086_, _12057_);
  and _20416_ (_12088_, _12087_, _12084_);
  and _20417_ (_12089_, _12088_, _12060_);
  and _20418_ (_12091_, _12089_, _12053_);
  and _20419_ (_12092_, _12091_, _12050_);
  and _20420_ (_12093_, _12092_, _12046_);
  and _20421_ (_12094_, _12093_, _12042_);
  and _20422_ (_12095_, _12094_, _12038_);
  and _20423_ (_12096_, _12095_, _12034_);
  nand _20424_ (_12097_, _12096_, _12030_);
  or _20425_ (_12099_, _12097_, _12027_);
  or _20426_ (_12100_, _12099_, _12025_);
  or _20427_ (_12101_, _12100_, _12023_);
  nand _20428_ (_12103_, _12100_, _12023_);
  and _20429_ (_12105_, _12103_, _12101_);
  or _20430_ (_12106_, _12105_, _07135_);
  or _20431_ (_12107_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _20432_ (_12108_, rst, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _20433_ (_12110_, _12108_, _12107_);
  and _20434_ (_12111_, _12110_, _12106_);
  or _20435_ (_10640_, _12111_, _11977_);
  and _20436_ (_12112_, _06782_, _06550_);
  and _20437_ (_12114_, _08333_, _06544_);
  nor _20438_ (_12115_, _12114_, _12112_);
  and _20439_ (_12117_, _06760_, _06565_);
  and _20440_ (_12118_, _06767_, _06550_);
  nor _20441_ (_12120_, _12118_, _12117_);
  nand _20442_ (_12121_, _12120_, _12115_);
  nor _20443_ (_12123_, _12121_, _07040_);
  and _20444_ (_12124_, _06566_, _06550_);
  or _20445_ (_12126_, _12124_, _06559_);
  nor _20446_ (_12127_, _12126_, _07056_);
  or _20447_ (_12129_, _07047_, _06990_);
  and _20448_ (_12130_, _06544_, _06572_);
  or _20449_ (_12131_, _12130_, _07073_);
  nor _20450_ (_12132_, _12131_, _12129_);
  and _20451_ (_12133_, _12132_, _12127_);
  nand _20452_ (_12135_, _06768_, _06760_);
  and _20453_ (_12136_, _06760_, _07053_);
  or _20454_ (_12138_, _12136_, _06994_);
  and _20455_ (_12139_, _11428_, _06760_);
  nor _20456_ (_12141_, _12139_, _12138_);
  and _20457_ (_12142_, _12141_, _12135_);
  and _20458_ (_12144_, _06760_, _06529_);
  or _20459_ (_12145_, _07067_, _07044_);
  nor _20460_ (_12147_, _12145_, _12144_);
  nor _20461_ (_12148_, _07063_, _06799_);
  and _20462_ (_12149_, _12148_, _11438_);
  and _20463_ (_12150_, _12149_, _12147_);
  and _20464_ (_12151_, _12150_, _12142_);
  and _20465_ (_12152_, _12151_, _12133_);
  nand _20466_ (_12153_, _12152_, _12123_);
  nand _20467_ (_12155_, _12153_, _06821_);
  nor _20468_ (_12156_, _11451_, _08341_);
  nand _20469_ (_12158_, _12156_, _12155_);
  nand _20470_ (_12159_, _12158_, _05143_);
  and _20471_ (_12161_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _20472_ (_12162_, _12161_);
  nand _20473_ (_12164_, _12162_, _12159_);
  not _20474_ (_12165_, _11425_);
  or _20475_ (_12166_, _11456_, _12165_);
  or _20476_ (_12167_, _12166_, _12164_);
  or _20477_ (_12168_, _12167_, _11848_);
  and _20478_ (_12169_, _12162_, _12159_);
  or _20479_ (_12170_, _12166_, _12169_);
  nor _20480_ (_12171_, _06271_, _05312_);
  nor _20481_ (_12172_, _06308_, _06427_);
  nor _20482_ (_12173_, _06314_, _06429_);
  nor _20483_ (_12174_, _12173_, _12172_);
  and _20484_ (_12175_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _20485_ (_12176_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _20486_ (_12177_, _12176_, _12175_);
  and _20487_ (_12178_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _20488_ (_12179_, _06320_, _06438_);
  nor _20489_ (_12181_, _12179_, _12178_);
  and _20490_ (_12182_, _12181_, _12177_);
  and _20491_ (_12184_, _12182_, _12174_);
  nor _20492_ (_12185_, _12184_, _07135_);
  nor _20493_ (_12186_, _12185_, _12171_);
  or _20494_ (_12188_, _12186_, _12170_);
  and _20495_ (_12189_, _12188_, _12168_);
  and _20496_ (_12191_, _12169_, _11456_);
  and _20497_ (_12192_, _12191_, _11425_);
  and _20498_ (_12193_, _11867_, _11845_);
  not _20499_ (_12194_, _11872_);
  nand _20500_ (_12195_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nand _20501_ (_12196_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _20502_ (_12197_, _12196_, _12195_);
  nand _20503_ (_12199_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nand _20504_ (_12200_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _20505_ (_12201_, _12200_, _12199_);
  and _20506_ (_12202_, _12201_, _12197_);
  or _20507_ (_12204_, _11863_, _06365_);
  or _20508_ (_12205_, _12204_, _11870_);
  or _20509_ (_12207_, _12205_, _08129_);
  nand _20510_ (_12208_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _20511_ (_12209_, _12208_, _12207_);
  nand _20512_ (_12211_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nand _20513_ (_12213_, _11878_, _11848_);
  or _20514_ (_12214_, _12213_, _06719_);
  and _20515_ (_12215_, _12214_, _12211_);
  and _20516_ (_12216_, _12215_, _12209_);
  and _20517_ (_12217_, _12216_, _11885_);
  and _20518_ (_12219_, _12217_, _12202_);
  nor _20519_ (_12220_, _12219_, _12193_);
  nand _20520_ (_12221_, _12220_, _12192_);
  or _20521_ (_12222_, _11456_, _11425_);
  nand _20522_ (_12223_, _12164_, _11456_);
  nor _20523_ (_12224_, _12223_, _12165_);
  and _20524_ (_12225_, _06621_, _05288_);
  and _20525_ (_12226_, _12225_, _05522_);
  nand _20526_ (_12228_, _06621_, _05288_);
  or _20527_ (_12229_, _12228_, _06062_);
  or _20528_ (_12230_, _12225_, _05152_);
  nand _20529_ (_12231_, _12230_, _12229_);
  or _20530_ (_12232_, _12225_, _05153_);
  or _20531_ (_12233_, _12228_, _05560_);
  nand _20532_ (_12234_, _12233_, _12232_);
  nand _20533_ (_12235_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  or _20534_ (_12236_, _12228_, _06178_);
  and _20535_ (_12237_, _12236_, _12235_);
  not _20536_ (_12238_, _12237_);
  not _20537_ (_12239_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  or _20538_ (_12240_, _12225_, _05192_);
  or _20539_ (_12241_, _12228_, _05604_);
  nand _20540_ (_12243_, _12241_, _12240_);
  or _20541_ (_12244_, _12243_, _12239_);
  or _20542_ (_12245_, _12244_, _12238_);
  or _20543_ (_12247_, _12245_, _12234_);
  nor _20544_ (_12248_, _12247_, _12231_);
  and _20545_ (_12249_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _20546_ (_12250_, _12249_, _12226_);
  and _20547_ (_12251_, _12250_, _12248_);
  nor _20548_ (_12252_, _12250_, _12248_);
  or _20549_ (_12253_, _12252_, _12251_);
  nand _20550_ (_12254_, _12253_, _05243_);
  nand _20551_ (_12255_, _12254_, _05246_);
  and _20552_ (_12256_, _12255_, _12228_);
  or _20553_ (_12257_, _12256_, _12226_);
  nand _20554_ (_12258_, _12257_, _12224_);
  and _20555_ (_12259_, _12258_, _12222_);
  and _20556_ (_12260_, _12259_, _12221_);
  and _20557_ (_12261_, _12260_, _12189_);
  or _20558_ (_12262_, _12261_, _10341_);
  nand _20559_ (_12263_, _12260_, _12189_);
  or _20560_ (_12264_, _12263_, _05256_);
  and _20561_ (_12265_, _12264_, _12262_);
  and _20562_ (_12266_, _11456_, _12165_);
  nand _20563_ (_12267_, _12266_, _12164_);
  or _20564_ (_12268_, _12170_, _07514_);
  nor _20565_ (_12269_, _11885_, _06004_);
  nand _20566_ (_12270_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand _20567_ (_12271_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _20568_ (_12272_, _12271_, _12270_);
  nand _20569_ (_12273_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _20570_ (_12274_, _12205_, _08237_);
  and _20571_ (_12275_, _12274_, _12273_);
  and _20572_ (_12276_, _12275_, _12272_);
  or _20573_ (_12277_, _11872_, _07096_);
  nand _20574_ (_12278_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _20575_ (_12279_, _12278_, _12277_);
  nand _20576_ (_12280_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nand _20577_ (_12281_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _20578_ (_12282_, _12281_, _12280_);
  and _20579_ (_12283_, _12282_, _12279_);
  and _20580_ (_12285_, _12283_, _11885_);
  and _20581_ (_12286_, _12285_, _12276_);
  or _20582_ (_12287_, _12286_, _12269_);
  not _20583_ (_12288_, _12287_);
  nand _20584_ (_12289_, _12288_, _12192_);
  and _20585_ (_12290_, _12289_, _12268_);
  or _20586_ (_12291_, _12223_, _12165_);
  and _20587_ (_12292_, _12225_, _06004_);
  not _20588_ (_12293_, _12292_);
  and _20589_ (_12294_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _20590_ (_12296_, _12294_, _12292_);
  nand _20591_ (_12297_, _12296_, _12251_);
  or _20592_ (_12299_, _12296_, _12251_);
  and _20593_ (_12300_, _12299_, _12297_);
  or _20594_ (_12301_, _12300_, _05159_);
  and _20595_ (_12302_, _12301_, _05259_);
  or _20596_ (_12303_, _12302_, _12225_);
  and _20597_ (_12304_, _12303_, _12293_);
  or _20598_ (_12305_, _12304_, _12291_);
  or _20599_ (_12306_, _12222_, _12164_);
  and _20600_ (_12308_, _12306_, _12305_);
  and _20601_ (_12309_, _12308_, _12290_);
  and _20602_ (_12310_, _12309_, _12267_);
  and _20603_ (_12312_, _12310_, _05280_);
  nand _20604_ (_12313_, _12309_, _12267_);
  and _20605_ (_12314_, _12313_, _05266_);
  nor _20606_ (_12315_, _12314_, _12312_);
  and _20607_ (_12317_, _12315_, _12265_);
  and _20608_ (_12318_, _12247_, _12231_);
  nor _20609_ (_12319_, _12318_, _12248_);
  nor _20610_ (_12320_, _12319_, _05159_);
  not _20611_ (_12321_, _12320_);
  nand _20612_ (_12322_, _12321_, _05162_);
  nand _20613_ (_12323_, _12322_, _12228_);
  nand _20614_ (_12325_, _12323_, _12229_);
  nand _20615_ (_12326_, _12325_, _12224_);
  or _20616_ (_12327_, _12167_, _11863_);
  nand _20617_ (_12329_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nand _20618_ (_12330_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _20619_ (_12331_, _12330_, _12329_);
  nand _20620_ (_12332_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nand _20621_ (_12333_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _20622_ (_12335_, _12333_, _12332_);
  and _20623_ (_12336_, _12335_, _12331_);
  or _20624_ (_12338_, _12205_, _08076_);
  or _20625_ (_12339_, _12213_, _08487_);
  and _20626_ (_12340_, _12339_, _12338_);
  nand _20627_ (_12341_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nand _20628_ (_12343_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _20629_ (_12344_, _12343_, _12341_);
  and _20630_ (_12346_, _12344_, _12340_);
  and _20631_ (_12347_, _12346_, _11885_);
  nand _20632_ (_12349_, _12347_, _12336_);
  nand _20633_ (_12350_, _11867_, _06062_);
  and _20634_ (_12351_, _12350_, _12349_);
  nand _20635_ (_12352_, _12351_, _12192_);
  nor _20636_ (_12354_, _06271_, _05385_);
  nor _20637_ (_12355_, _06308_, _06403_);
  nor _20638_ (_12356_, _06314_, _06395_);
  nor _20639_ (_12357_, _12356_, _12355_);
  and _20640_ (_12358_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _20641_ (_12359_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _20642_ (_12361_, _12359_, _12358_);
  nor _20643_ (_12362_, _06304_, _06399_);
  nor _20644_ (_12363_, _06320_, _06406_);
  nor _20645_ (_12364_, _12363_, _12362_);
  and _20646_ (_12365_, _12364_, _12361_);
  and _20647_ (_12366_, _12365_, _12357_);
  nor _20648_ (_12367_, _12366_, _07135_);
  nor _20649_ (_12368_, _12367_, _12354_);
  or _20650_ (_12369_, _12368_, _12170_);
  and _20651_ (_12370_, _12369_, _12352_);
  and _20652_ (_12371_, _12370_, _12327_);
  and _20653_ (_12372_, _12371_, _12326_);
  or _20654_ (_12373_, _12372_, _05173_);
  nand _20655_ (_12374_, _12371_, _12326_);
  or _20656_ (_12375_, _12374_, _05172_);
  and _20657_ (_12376_, _12375_, _12373_);
  and _20658_ (_12377_, _12225_, _05960_);
  not _20659_ (_12378_, _12297_);
  nor _20660_ (_12379_, _12228_, _06244_);
  and _20661_ (_12380_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _20662_ (_12381_, _12380_, _12379_);
  and _20663_ (_12382_, _12381_, _12378_);
  and _20664_ (_12383_, _12228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand _20665_ (_12384_, _12383_, _12382_);
  or _20666_ (_12385_, _12383_, _12382_);
  and _20667_ (_12386_, _12385_, _05243_);
  nand _20668_ (_12387_, _12386_, _12384_);
  and _20669_ (_12388_, _12228_, _05232_);
  and _20670_ (_12389_, _12388_, _12387_);
  nor _20671_ (_12390_, _12389_, _12377_);
  nand _20672_ (_12391_, _12390_, _12224_);
  and _20673_ (_12392_, _11901_, _12192_);
  and _20674_ (_12393_, _12223_, _12165_);
  nor _20675_ (_12394_, _12393_, _12392_);
  or _20676_ (_12395_, _12170_, _07137_);
  and _20677_ (_12396_, _12395_, _12267_);
  and _20678_ (_12397_, _12396_, _12394_);
  and _20679_ (_12398_, _12397_, _12391_);
  nand _20680_ (_12399_, _12398_, _05241_);
  or _20681_ (_12400_, _12398_, _05241_);
  and _20682_ (_12401_, _12400_, _12399_);
  nand _20683_ (_12402_, _12381_, _12378_);
  or _20684_ (_12403_, _12381_, _12378_);
  nand _20685_ (_12404_, _12403_, _12402_);
  nand _20686_ (_12405_, _12404_, _05243_);
  nand _20687_ (_12407_, _12405_, _05218_);
  and _20688_ (_12408_, _12407_, _12228_);
  or _20689_ (_12409_, _12408_, _12379_);
  nand _20690_ (_12410_, _12409_, _12224_);
  and _20691_ (_12411_, _12267_, _12222_);
  nor _20692_ (_12412_, _06271_, _05692_);
  nor _20693_ (_12413_, _06308_, _06514_);
  nor _20694_ (_12414_, _06314_, _06510_);
  nor _20695_ (_12415_, _12414_, _12413_);
  and _20696_ (_12416_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor _20697_ (_12417_, _06320_, _06516_);
  nor _20698_ (_12418_, _12417_, _12416_);
  and _20699_ (_12419_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _20700_ (_12420_, _06304_, _06508_);
  nor _20701_ (_12421_, _12420_, _12419_);
  and _20702_ (_12422_, _12421_, _12418_);
  and _20703_ (_12423_, _12422_, _12415_);
  nor _20704_ (_12424_, _12423_, _07135_);
  nor _20705_ (_12425_, _12424_, _12412_);
  or _20706_ (_12426_, _12425_, _12170_);
  nand _20707_ (_12427_, _11867_, _06244_);
  nand _20708_ (_12428_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nand _20709_ (_12429_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _20710_ (_12430_, _12429_, _12428_);
  nand _20711_ (_12431_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nand _20712_ (_12432_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _20713_ (_12433_, _12432_, _12431_);
  and _20714_ (_12434_, _12433_, _12430_);
  nand _20715_ (_12435_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nand _20716_ (_12436_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _20717_ (_12437_, _12436_, _12435_);
  nand _20718_ (_12438_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nand _20719_ (_12439_, _11893_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _20720_ (_12440_, _12439_, _12438_);
  and _20721_ (_12441_, _12440_, _12437_);
  and _20722_ (_12442_, _12441_, _11885_);
  nand _20723_ (_12443_, _12442_, _12434_);
  and _20724_ (_12444_, _12443_, _12427_);
  nand _20725_ (_12445_, _12444_, _12192_);
  and _20726_ (_12446_, _12445_, _12426_);
  and _20727_ (_12447_, _12446_, _12411_);
  nand _20728_ (_12448_, _12447_, _12410_);
  and _20729_ (_12449_, _12448_, _05227_);
  and _20730_ (_12450_, _12447_, _12410_);
  and _20731_ (_12451_, _12450_, _05228_);
  nor _20732_ (_12452_, _12451_, _12449_);
  and _20733_ (_12453_, _12452_, _12401_);
  and _20734_ (_12454_, _12453_, _12376_);
  and _20735_ (_12455_, _12454_, _12317_);
  nor _20736_ (_12456_, _12243_, _12239_);
  and _20737_ (_12457_, _12243_, _12239_);
  nor _20738_ (_12458_, _12457_, _12456_);
  nor _20739_ (_12459_, _12458_, _05159_);
  nor _20740_ (_12460_, _12459_, _05193_);
  nor _20741_ (_12461_, _12460_, _12225_);
  not _20742_ (_12462_, _12461_);
  and _20743_ (_12463_, _12462_, _12241_);
  or _20744_ (_12464_, _12463_, _12291_);
  or _20745_ (_12465_, _12167_, _06365_);
  nand _20746_ (_12466_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or _20747_ (_12467_, _12213_, _09779_);
  and _20748_ (_12468_, _12467_, _12466_);
  nand _20749_ (_12469_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or _20750_ (_12470_, _12205_, _05621_);
  and _20751_ (_12471_, _12470_, _12469_);
  and _20752_ (_12472_, _12471_, _12468_);
  nand _20753_ (_12473_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand _20754_ (_12474_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _20755_ (_12475_, _12474_, _12473_);
  nand _20756_ (_12476_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nand _20757_ (_12477_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _20758_ (_12478_, _12477_, _12476_);
  and _20759_ (_12479_, _12478_, _12475_);
  and _20760_ (_12480_, _12479_, _11885_);
  nand _20761_ (_12481_, _12480_, _12472_);
  nand _20762_ (_12482_, _11867_, _05604_);
  and _20763_ (_12483_, _12482_, _12481_);
  nand _20764_ (_12484_, _12483_, _12192_);
  nor _20765_ (_12485_, _06271_, _05406_);
  nor _20766_ (_12486_, _06308_, _06351_);
  nor _20767_ (_12487_, _06314_, _06343_);
  nor _20768_ (_12488_, _12487_, _12486_);
  and _20769_ (_12489_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _20770_ (_12490_, _06320_, _06353_);
  nor _20771_ (_12491_, _12490_, _12489_);
  and _20772_ (_12492_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _20773_ (_12493_, _06304_, _06347_);
  nor _20774_ (_12494_, _12493_, _12492_);
  and _20775_ (_12495_, _12494_, _12491_);
  and _20776_ (_12496_, _12495_, _12488_);
  nor _20777_ (_12497_, _12496_, _07135_);
  nor _20778_ (_12498_, _12497_, _12485_);
  or _20779_ (_12499_, _12498_, _12170_);
  and _20780_ (_12500_, _12499_, _12484_);
  and _20781_ (_12501_, _12500_, _12465_);
  and _20782_ (_12502_, _12501_, _12464_);
  or _20783_ (_12503_, _12502_, _05197_);
  nand _20784_ (_12504_, _12501_, _12464_);
  or _20785_ (_12505_, _12504_, _05286_);
  nand _20786_ (_12506_, _12505_, _12503_);
  and _20787_ (_12507_, _12506_, _05646_);
  and _20788_ (_12508_, _12244_, _12238_);
  not _20789_ (_12509_, _12508_);
  and _20790_ (_12510_, _12509_, _12245_);
  nor _20791_ (_12511_, _12510_, _05159_);
  nor _20792_ (_12512_, _12511_, _05200_);
  nor _20793_ (_12513_, _12512_, _12225_);
  not _20794_ (_12514_, _12513_);
  and _20795_ (_12515_, _12514_, _12236_);
  or _20796_ (_12516_, _12515_, _12291_);
  nand _20797_ (_12517_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nand _20798_ (_12518_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _20799_ (_12519_, _12518_, _12517_);
  nand _20800_ (_12520_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand _20801_ (_12521_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _20802_ (_12522_, _12521_, _12520_);
  and _20803_ (_12523_, _12522_, _12519_);
  nand _20804_ (_12524_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nand _20805_ (_12525_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _20806_ (_12526_, _12525_, _12524_);
  or _20807_ (_12527_, _12205_, _08155_);
  nand _20808_ (_12528_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _20809_ (_12529_, _12528_, _12527_);
  and _20810_ (_12530_, _12529_, _12526_);
  and _20811_ (_12531_, _12530_, _11885_);
  nand _20812_ (_12532_, _12531_, _12523_);
  nand _20813_ (_12533_, _11867_, _06178_);
  and _20814_ (_12534_, _12533_, _12532_);
  nand _20815_ (_12535_, _12534_, _12192_);
  nor _20816_ (_12537_, _06271_, _05430_);
  nor _20817_ (_12538_, _06308_, _06301_);
  nor _20818_ (_12539_, _06314_, _06306_);
  nor _20819_ (_12540_, _12539_, _12538_);
  and _20820_ (_12541_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _20821_ (_12542_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _20822_ (_12543_, _12542_, _12541_);
  nor _20823_ (_12544_, _06304_, _06324_);
  nor _20824_ (_12545_, _06320_, _06311_);
  nor _20825_ (_12546_, _12545_, _12544_);
  and _20826_ (_12547_, _12546_, _12543_);
  and _20827_ (_12548_, _12547_, _12540_);
  nor _20828_ (_12549_, _12548_, _07135_);
  nor _20829_ (_12550_, _12549_, _12537_);
  or _20830_ (_12551_, _12550_, _12170_);
  and _20831_ (_12552_, _12551_, _12535_);
  nand _20832_ (_12553_, _12266_, _12169_);
  or _20833_ (_12554_, _12167_, _06339_);
  and _20834_ (_12555_, _12554_, _12553_);
  and _20835_ (_12556_, _12555_, _12552_);
  and _20836_ (_12557_, _12556_, _12516_);
  and _20837_ (_12558_, _12557_, _05274_);
  nand _20838_ (_12559_, _12556_, _12516_);
  and _20839_ (_12560_, _12559_, _05208_);
  nor _20840_ (_12561_, _12560_, _12558_);
  and _20841_ (_12562_, _12245_, _12234_);
  not _20842_ (_12563_, _12562_);
  and _20843_ (_12564_, _12563_, _12247_);
  nor _20844_ (_12565_, _12564_, _05159_);
  nor _20845_ (_12566_, _12565_, _05178_);
  nor _20846_ (_12567_, _12566_, _12225_);
  not _20847_ (_12568_, _12567_);
  and _20848_ (_12569_, _12568_, _12233_);
  or _20849_ (_12570_, _12569_, _12291_);
  nand _20850_ (_12571_, _12194_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nand _20851_ (_12572_, _11881_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _20852_ (_12573_, _12572_, _12571_);
  nand _20853_ (_12574_, _11887_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or _20854_ (_12575_, _12205_, _08132_);
  and _20855_ (_12576_, _12575_, _12574_);
  and _20856_ (_12577_, _12576_, _12573_);
  nand _20857_ (_12578_, _11879_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nand _20858_ (_12579_, _11895_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _20859_ (_12580_, _12579_, _12578_);
  nand _20860_ (_12581_, _11889_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nand _20861_ (_12582_, _11875_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _20862_ (_12583_, _12582_, _12581_);
  and _20863_ (_12584_, _12583_, _12580_);
  and _20864_ (_12585_, _12584_, _11885_);
  and _20865_ (_12586_, _12585_, _12577_);
  and _20866_ (_12587_, _11867_, _05560_);
  nor _20867_ (_12588_, _12587_, _12586_);
  nand _20868_ (_12589_, _12588_, _12192_);
  or _20869_ (_12590_, _12167_, _06533_);
  nor _20870_ (_12591_, _06271_, _05447_);
  nor _20871_ (_12592_, _06308_, _06376_);
  nor _20872_ (_12593_, _06314_, _06374_);
  nor _20873_ (_12594_, _12593_, _12592_);
  and _20874_ (_12595_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _20875_ (_12596_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _20876_ (_12597_, _12596_, _12595_);
  nor _20877_ (_12598_, _06304_, _06379_);
  nor _20878_ (_12599_, _06320_, _06370_);
  nor _20879_ (_12600_, _12599_, _12598_);
  and _20880_ (_12601_, _12600_, _12597_);
  and _20881_ (_12602_, _12601_, _12594_);
  nor _20882_ (_12603_, _12602_, _07135_);
  nor _20883_ (_12604_, _12603_, _12591_);
  or _20884_ (_12605_, _12604_, _12170_);
  and _20885_ (_12606_, _12605_, _12590_);
  and _20886_ (_12607_, _12606_, _12589_);
  and _20887_ (_12608_, _12607_, _12570_);
  or _20888_ (_12609_, _12608_, _05186_);
  nand _20889_ (_12610_, _12607_, _12570_);
  or _20890_ (_12611_, _12610_, _06007_);
  nand _20891_ (_12612_, _12611_, _12609_);
  and _20892_ (_12613_, _12612_, _12561_);
  and _20893_ (_12614_, _12613_, _12507_);
  and _20894_ (_12615_, _12614_, _12455_);
  and _20895_ (_12616_, _05241_, _05295_);
  nand _20896_ (_12617_, _12616_, _12615_);
  not _20897_ (_12618_, _08171_);
  and _20898_ (_12619_, _11452_, _12618_);
  not _20899_ (_12621_, _06846_);
  and _20900_ (_12622_, _06563_, _06550_);
  nor _20901_ (_12624_, _12622_, _06575_);
  not _20902_ (_12625_, _12624_);
  and _20903_ (_12626_, _12625_, _07088_);
  not _20904_ (_12627_, _06558_);
  nor _20905_ (_12628_, _12124_, _06554_);
  and _20906_ (_12629_, _12628_, _12627_);
  and _20907_ (_12631_, _12622_, _07088_);
  not _20908_ (_12632_, _12631_);
  and _20909_ (_12633_, _12632_, _12629_);
  nor _20910_ (_12634_, _12633_, _06791_);
  nor _20911_ (_12635_, _12634_, _12626_);
  and _20912_ (_12636_, _06588_, _05824_);
  nand _20913_ (_12637_, _12636_, _07322_);
  nor _20914_ (_12638_, _12637_, _07233_);
  and _20915_ (_12639_, _12638_, _07171_);
  and _20916_ (_12640_, _12639_, _06662_);
  and _20917_ (_12642_, _12640_, _07487_);
  and _20918_ (_12643_, _12642_, _12635_);
  and _20919_ (_12644_, _12643_, _12621_);
  and _20920_ (_12645_, _07088_, _06563_);
  and _20921_ (_12646_, _12645_, _06550_);
  not _20922_ (_12647_, _12646_);
  nor _20923_ (_12649_, _12646_, _12126_);
  nor _20924_ (_12650_, _12649_, _06791_);
  and _20925_ (_12651_, _12650_, _12647_);
  and _20926_ (_12652_, _12651_, _05379_);
  nor _20927_ (_12653_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _20928_ (_12654_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _20929_ (_12655_, _12654_, _12653_);
  nor _20930_ (_12657_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _20931_ (_12658_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _20932_ (_12659_, _12658_, _12657_);
  and _20933_ (_12660_, _12659_, _12655_);
  and _20934_ (_12662_, _12660_, _11452_);
  and _20935_ (_12663_, _12646_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _20936_ (_12664_, _12663_, _12662_);
  or _20937_ (_12665_, _12664_, _12652_);
  nor _20938_ (_12666_, _12665_, _12644_);
  and _20939_ (_12667_, _08340_, _06450_);
  nor _20940_ (_12668_, _12667_, _06559_);
  nor _20941_ (_12669_, _12668_, _12666_);
  or _20942_ (_12670_, _08334_, _06573_);
  and _20943_ (_12671_, _06767_, _06755_);
  nor _20944_ (_12672_, _12671_, _06981_);
  nor _20945_ (_12673_, _06774_, _12124_);
  nand _20946_ (_12674_, _12673_, _12672_);
  and _20947_ (_12675_, _06570_, _06417_);
  and _20948_ (_12676_, _08340_, _06449_);
  or _20949_ (_12677_, _12676_, _12675_);
  or _20950_ (_12678_, _12677_, _12674_);
  and _20951_ (_12679_, _12678_, _12666_);
  or _20952_ (_12680_, _12679_, _12670_);
  or _20953_ (_12681_, _12680_, _12669_);
  and _20954_ (_12682_, _12681_, _07088_);
  and _20955_ (_12683_, _06552_, _06544_);
  nor _20956_ (_12684_, _12683_, _06816_);
  nor _20957_ (_12685_, _12684_, _08330_);
  nor _20958_ (_12686_, _12685_, _11450_);
  not _20959_ (_12687_, _12686_);
  nor _20960_ (_12688_, _12687_, _12682_);
  nor _20961_ (_12689_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _20962_ (_12690_, _12689_);
  nor _20963_ (_12691_, _10354_, _12690_);
  and _20964_ (_12692_, _12691_, _10376_);
  nor _20965_ (_12693_, _12692_, _12632_);
  or _20966_ (_12694_, _12693_, _12688_);
  nor _20967_ (_12695_, _12694_, _12619_);
  nor _20968_ (_12696_, _06735_, _06008_);
  and _20969_ (_12697_, _12696_, _12455_);
  nand _20970_ (_12698_, _12697_, _12651_);
  and _20971_ (_12699_, _12698_, _12695_);
  and _20972_ (_12700_, _12699_, _12617_);
  and _20973_ (_12701_, _08334_, _07088_);
  and _20974_ (_12702_, _12701_, _06975_);
  not _20975_ (_12703_, _11451_);
  nor _20976_ (_12704_, _12703_, _06875_);
  and _20977_ (_12705_, _06821_, _06556_);
  and _20978_ (_12706_, _12705_, _06550_);
  and _20979_ (_12707_, _12683_, _06821_);
  or _20980_ (_12708_, _12707_, _12706_);
  nor _20981_ (_12709_, _12708_, _11451_);
  or _20982_ (_12710_, _12674_, _06559_);
  nand _20983_ (_12711_, _12710_, _07088_);
  and _20984_ (_12712_, _12711_, _12709_);
  and _20985_ (_12713_, _12712_, _12685_);
  nand _20986_ (_12714_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _20987_ (_12715_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or _20988_ (_12716_, _12715_, _12714_);
  nand _20989_ (_12717_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand _20990_ (_12718_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _20991_ (_12719_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _20992_ (_12720_, _12719_, _12718_);
  or _20993_ (_12721_, _12720_, _12717_);
  or _20994_ (_12723_, _12721_, _12716_);
  or _20995_ (_12724_, _12723_, _05390_);
  or _20996_ (_12725_, _12724_, _05317_);
  or _20997_ (_12726_, _12725_, _05739_);
  or _20998_ (_12727_, _12726_, _05699_);
  and _20999_ (_12728_, _12727_, _05663_);
  nor _21000_ (_12729_, _12727_, _05663_);
  nor _21001_ (_12730_, _12729_, _12728_);
  and _21002_ (_12731_, _12730_, _12713_);
  not _21003_ (_12732_, _07137_);
  and _21004_ (_12733_, _12707_, _12732_);
  nor _21005_ (_12735_, _12701_, _12685_);
  nand _21006_ (_12736_, _12735_, _12712_);
  or _21007_ (_12737_, _08340_, _12675_);
  nor _21008_ (_12739_, _12737_, _06774_);
  nand _21009_ (_12740_, _12739_, _12672_);
  or _21010_ (_12741_, _12670_, _12126_);
  or _21011_ (_12742_, _12741_, _12740_);
  and _21012_ (_12743_, _12742_, _07088_);
  or _21013_ (_12744_, _12743_, _12706_);
  nor _21014_ (_12745_, _12744_, _12736_);
  and _21015_ (_12746_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _21016_ (_12747_, _12746_, _12733_);
  or _21017_ (_12748_, _12747_, _12731_);
  or _21018_ (_12749_, _12748_, _12704_);
  nor _21019_ (_12750_, _12749_, _12702_);
  nand _21020_ (_12751_, _12750_, _12700_);
  nand _21021_ (_12752_, _12712_, _12732_);
  nor _21022_ (_12753_, _06271_, _05658_);
  and _21023_ (_12754_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21024_ (_12755_, _06308_, _06457_);
  nor _21025_ (_12756_, _06320_, _06462_);
  nor _21026_ (_12757_, _12756_, _12755_);
  and _21027_ (_12758_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _21028_ (_12759_, _06314_, _06459_);
  nor _21029_ (_12760_, _12759_, _12758_);
  and _21030_ (_12761_, _12760_, _12757_);
  and _21031_ (_12762_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _21032_ (_12763_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _21033_ (_12764_, _12763_, _12762_);
  and _21034_ (_12765_, _12764_, _12761_);
  nor _21035_ (_12766_, _12765_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21036_ (_12768_, _12766_, _12754_);
  nor _21037_ (_12769_, _12768_, _07516_);
  nor _21038_ (_12770_, _12769_, _12753_);
  or _21039_ (_12771_, _12770_, _12712_);
  and _21040_ (_12772_, _12771_, _12752_);
  not _21041_ (_12773_, _12772_);
  nor _21042_ (_12774_, \oc8051_top_1.oc8051_memory_interface1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _21043_ (_12775_, _12772_, _05665_);
  not _21044_ (_12776_, _12425_);
  nand _21045_ (_12777_, _12712_, _12776_);
  nor _21046_ (_12778_, _06271_, _05694_);
  and _21047_ (_12779_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21048_ (_12780_, _06308_, _06508_);
  nor _21049_ (_12781_, _06320_, _06510_);
  nor _21050_ (_12782_, _12781_, _12780_);
  and _21051_ (_12783_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor _21052_ (_12784_, _06314_, _06514_);
  nor _21053_ (_12785_, _12784_, _12783_);
  and _21054_ (_12786_, _12785_, _12782_);
  and _21055_ (_12787_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _21056_ (_12789_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _21057_ (_12790_, _12789_, _12787_);
  and _21058_ (_12792_, _12790_, _12786_);
  nor _21059_ (_12793_, _12792_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21060_ (_12794_, _12793_, _12779_);
  nor _21061_ (_12795_, _12794_, _07516_);
  nor _21062_ (_12796_, _12795_, _12778_);
  or _21063_ (_12797_, _12796_, _12712_);
  nand _21064_ (_12798_, _12797_, _12777_);
  nand _21065_ (_12799_, _12798_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _21066_ (_12800_, _12799_);
  nand _21067_ (_12801_, _12772_, _05665_);
  and _21068_ (_12802_, _12801_, _12775_);
  nand _21069_ (_12803_, _12802_, _12800_);
  nand _21070_ (_12804_, _12803_, _12775_);
  or _21071_ (_12805_, _12798_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _21072_ (_12806_, _12805_, _12799_);
  and _21073_ (_12807_, _12806_, _12802_);
  not _21074_ (_12808_, _07514_);
  nand _21075_ (_12809_, _12712_, _12808_);
  nor _21076_ (_12810_, _06271_, _05734_);
  and _21077_ (_12811_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21078_ (_12812_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor _21079_ (_12813_, _06320_, _06484_);
  nor _21080_ (_12814_, _12813_, _12812_);
  nor _21081_ (_12816_, _06308_, _06482_);
  and _21082_ (_12817_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _21083_ (_12818_, _12817_, _12816_);
  and _21084_ (_12819_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _21085_ (_12820_, _06314_, _06487_);
  nor _21086_ (_12821_, _12820_, _12819_);
  and _21087_ (_12822_, _12821_, _12818_);
  and _21088_ (_12823_, _12822_, _12814_);
  nor _21089_ (_12824_, _12823_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21090_ (_12825_, _12824_, _12811_);
  nor _21091_ (_12826_, _12825_, _07516_);
  nor _21092_ (_12827_, _12826_, _12810_);
  or _21093_ (_12828_, _12827_, _12712_);
  and _21094_ (_12829_, _12828_, _12809_);
  or _21095_ (_12830_, _12829_, _05742_);
  not _21096_ (_12831_, _12186_);
  nand _21097_ (_12832_, _12712_, _12831_);
  or _21098_ (_12833_, _12712_, _07593_);
  nand _21099_ (_12834_, _12833_, _12832_);
  nand _21100_ (_12835_, _12834_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand _21101_ (_12836_, _12829_, _05742_);
  and _21102_ (_12837_, _12836_, _12830_);
  not _21103_ (_12838_, _12837_);
  or _21104_ (_12839_, _12838_, _12835_);
  nand _21105_ (_12840_, _12839_, _12830_);
  and _21106_ (_12841_, _12840_, _12807_);
  or _21107_ (_12842_, _12841_, _12804_);
  not _21108_ (_12843_, _12368_);
  and _21109_ (_12844_, _12712_, _12843_);
  nor _21110_ (_12845_, _12712_, _07572_);
  nor _21111_ (_12846_, _12845_, _12844_);
  and _21112_ (_12847_, _12846_, _05388_);
  nor _21113_ (_12848_, _12846_, _05388_);
  not _21114_ (_12849_, _12604_);
  nand _21115_ (_12850_, _12712_, _12849_);
  or _21116_ (_12851_, _12712_, _07550_);
  and _21117_ (_12852_, _12851_, _12850_);
  nor _21118_ (_12853_, _12852_, _05453_);
  not _21119_ (_12855_, _12550_);
  nand _21120_ (_12857_, _12712_, _12855_);
  nor _21121_ (_12859_, _06271_, _05432_);
  and _21122_ (_12860_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _21123_ (_12862_, _07524_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor _21124_ (_12863_, _06320_, _06306_);
  nor _21125_ (_12864_, _12863_, _12862_);
  and _21126_ (_12865_, _06425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor _21127_ (_12866_, _06314_, _06301_);
  nor _21128_ (_12867_, _12866_, _12865_);
  and _21129_ (_12868_, _06328_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _21130_ (_12869_, _06308_, _06324_);
  nor _21131_ (_12870_, _12869_, _12868_);
  and _21132_ (_12871_, _12870_, _12867_);
  and _21133_ (_12872_, _12871_, _12864_);
  nor _21134_ (_12873_, _12872_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21135_ (_12874_, _12873_, _12860_);
  nor _21136_ (_12875_, _12874_, _07516_);
  nor _21137_ (_12876_, _12875_, _12859_);
  or _21138_ (_12877_, _12876_, _12712_);
  and _21139_ (_12878_, _12877_, _12857_);
  nor _21140_ (_12879_, _12878_, _05438_);
  not _21141_ (_12880_, _12498_);
  and _21142_ (_12881_, _12712_, _12880_);
  nor _21143_ (_12882_, _12712_, _07533_);
  or _21144_ (_12883_, _12882_, _12881_);
  and _21145_ (_12884_, _12883_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _21146_ (_12885_, _12879_);
  nand _21147_ (_12886_, _12878_, _05438_);
  and _21148_ (_12887_, _12886_, _12885_);
  and _21149_ (_12888_, _12887_, _12884_);
  or _21150_ (_12889_, _12888_, _12879_);
  not _21151_ (_12890_, _12853_);
  nand _21152_ (_12891_, _12852_, _05453_);
  and _21153_ (_12892_, _12891_, _12890_);
  and _21154_ (_12893_, _12892_, _12889_);
  or _21155_ (_12894_, _12893_, _12853_);
  nor _21156_ (_12895_, _12894_, _12848_);
  nor _21157_ (_12896_, _12895_, _12847_);
  or _21158_ (_12897_, _12834_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _21159_ (_12898_, _12897_, _12835_);
  and _21160_ (_12899_, _12837_, _12898_);
  and _21161_ (_12900_, _12899_, _12807_);
  and _21162_ (_12901_, _12900_, _12896_);
  or _21163_ (_12902_, _12901_, _12842_);
  or _21164_ (_12903_, _12902_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _21165_ (_12904_, _12903_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _21166_ (_12905_, _12904_, _12774_);
  and _21167_ (_12906_, _12905_, _05317_);
  and _21168_ (_12907_, _12906_, _05739_);
  nand _21169_ (_12908_, _12907_, _05699_);
  nand _21170_ (_12909_, _12908_, _12773_);
  and _21171_ (_12910_, \oc8051_top_1.oc8051_memory_interface1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _21172_ (_12911_, _12910_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _21173_ (_12912_, _12902_, _12911_);
  nand _21174_ (_12913_, _12912_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _21175_ (_12914_, _12913_, _05317_);
  nor _21176_ (_12915_, _12914_, _05739_);
  nand _21177_ (_12916_, _12915_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _21178_ (_12917_, _12916_, _12772_);
  nand _21179_ (_12918_, _12917_, _12909_);
  nand _21180_ (_12919_, _12918_, _05663_);
  or _21181_ (_12920_, _12918_, _05663_);
  and _21182_ (_12921_, _12920_, _12919_);
  not _21183_ (_12922_, _12712_);
  or _21184_ (_12923_, _12735_, _12922_);
  and _21185_ (_12924_, _06821_, _06550_);
  and _21186_ (_12926_, _12924_, _06556_);
  and _21187_ (_12927_, _06778_, _06766_);
  nor _21188_ (_12928_, _12927_, _11441_);
  nand _21189_ (_12929_, _12928_, _12624_);
  or _21190_ (_12930_, _12929_, _12670_);
  and _21191_ (_12931_, _06767_, _06420_);
  and _21192_ (_12932_, _06767_, _06760_);
  or _21193_ (_12933_, _12932_, _12931_);
  or _21194_ (_12934_, _12933_, _06981_);
  nor _21195_ (_12935_, _12934_, _06988_);
  nand _21196_ (_12936_, _12935_, _12629_);
  or _21197_ (_12937_, _12936_, _12930_);
  and _21198_ (_12938_, _12937_, _07088_);
  or _21199_ (_12939_, _12938_, _12926_);
  and _21200_ (_12940_, _12939_, _12923_);
  and _21201_ (_12941_, _12940_, _12921_);
  or _21202_ (_12942_, _12941_, _12751_);
  and _21203_ (_12943_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _21204_ (_12944_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _21205_ (_12945_, _12944_, _12943_);
  and _21206_ (_12946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _21207_ (_12947_, _12946_, _12945_);
  and _21208_ (_12948_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _21209_ (_12949_, _12948_, _12947_);
  and _21210_ (_12950_, _12949_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _21211_ (_12951_, _07619_);
  and _21212_ (_12952_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _21213_ (_12953_, _12952_, _12951_);
  and _21214_ (_12954_, _12953_, _12950_);
  and _21215_ (_12955_, _12954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _21216_ (_12956_, _12955_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _21217_ (_12957_, _12956_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _21218_ (_12958_, _12956_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _21219_ (_12959_, _12958_, _12957_);
  or _21220_ (_12960_, _12959_, _12700_);
  and _21221_ (_12961_, _12960_, _05141_);
  and _21222_ (_10647_, _12961_, _12942_);
  and _21223_ (_10656_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _05141_);
  nor _21224_ (_12962_, _12089_, _12053_);
  nor _21225_ (_12963_, _12962_, _12091_);
  or _21226_ (_12964_, _12963_, _07135_);
  or _21227_ (_12965_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _21228_ (_12966_, _12965_, _12108_);
  and _21229_ (_12967_, _12966_, _12964_);
  and _21230_ (_12968_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _21231_ (_10698_, _12968_, _12967_);
  or _21232_ (_12969_, _12905_, _12772_);
  nand _21233_ (_12970_, _12913_, _12772_);
  nand _21234_ (_12971_, _12970_, _12969_);
  nand _21235_ (_12972_, _12971_, _05317_);
  and _21236_ (_12973_, _12744_, _12923_);
  or _21237_ (_12974_, _12971_, _05317_);
  and _21238_ (_12975_, _12974_, _12973_);
  and _21239_ (_12976_, _12975_, _12972_);
  and _21240_ (_12977_, _12701_, _07229_);
  and _21241_ (_12978_, _12707_, _12831_);
  and _21242_ (_12979_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _21243_ (_12980_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _21244_ (_12981_, _12980_, _12979_);
  and _21245_ (_12982_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _21246_ (_12983_, _12982_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _21247_ (_12984_, _12983_, _12911_);
  and _21248_ (_12985_, _12984_, _12981_);
  and _21249_ (_12986_, _12985_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _21250_ (_12987_, _12986_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _21251_ (_12988_, _12987_, _12725_);
  and _21252_ (_12989_, _12988_, _12713_);
  or _21253_ (_12990_, _12989_, _12978_);
  and _21254_ (_12991_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _21255_ (_12992_, _12703_, _07259_);
  or _21256_ (_12993_, _12992_, _12991_);
  or _21257_ (_12995_, _12993_, _12990_);
  nor _21258_ (_12996_, _12995_, _12977_);
  nand _21259_ (_12997_, _12996_, _12700_);
  or _21260_ (_12998_, _12997_, _12976_);
  and _21261_ (_12999_, _12947_, _12951_);
  and _21262_ (_13000_, _12999_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _21263_ (_13001_, _13000_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _21264_ (_13002_, _13001_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _21265_ (_13003_, _13002_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _21266_ (_13004_, _13003_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nand _21267_ (_13005_, _13003_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _21268_ (_13006_, _13005_, _13004_);
  or _21269_ (_13007_, _13006_, _12700_);
  and _21270_ (_13008_, _13007_, _05141_);
  and _21271_ (_10715_, _13008_, _12998_);
  nand _21272_ (_13009_, _08396_, _05960_);
  and _21273_ (_13010_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _21274_ (_13011_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _21275_ (_13012_, _13011_, _13010_);
  or _21276_ (_13013_, _13012_, _08243_);
  and _21277_ (_13014_, _13013_, _05141_);
  and _21278_ (_10718_, _13014_, _13009_);
  and _21279_ (_13015_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _21280_ (_13016_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or _21281_ (_13017_, _13016_, _13015_);
  and _21282_ (_10742_, _13017_, _05141_);
  or _21283_ (_13018_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand _21284_ (_13019_, _07619_, _06508_);
  and _21285_ (_13020_, _13019_, _05141_);
  and _21286_ (_10747_, _13020_, _13018_);
  or _21287_ (_13022_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand _21288_ (_13023_, _07619_, _06301_);
  and _21289_ (_13024_, _13023_, _05141_);
  and _21290_ (_10750_, _13024_, _13022_);
  and _21291_ (_13025_, _08396_, _06283_);
  and _21292_ (_13026_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _21293_ (_13027_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _21294_ (_13028_, _13027_, _13026_);
  nor _21295_ (_13029_, _13028_, _08243_);
  not _21296_ (_13031_, _05960_);
  and _21297_ (_13032_, _08382_, _13031_);
  or _21298_ (_13033_, _13032_, _13029_);
  or _21299_ (_13034_, _13033_, _13025_);
  and _21300_ (_10792_, _13034_, _05141_);
  and _21301_ (_13035_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _21302_ (_13036_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _21303_ (_13037_, pc_log_change, _13036_);
  or _21304_ (_13038_, _13037_, _13035_);
  and _21305_ (_10800_, _13038_, _05141_);
  and _21306_ (_13039_, _08391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _21307_ (_13040_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor _21308_ (_13041_, _13040_, _13039_);
  nor _21309_ (_13042_, _13041_, _08243_);
  or _21310_ (_13043_, _08653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _21311_ (_13044_, _13043_, _08396_);
  or _21312_ (_13045_, _13044_, _13042_);
  and _21313_ (_10871_, _13045_, _05141_);
  and _21314_ (_13046_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _21315_ (_13047_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  or _21316_ (_13048_, _13047_, _13046_);
  and _21317_ (_10887_, _13048_, _05141_);
  or _21318_ (_13049_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _21319_ (_13050_, _07619_, _06376_);
  and _21320_ (_13051_, _13050_, _05141_);
  and _21321_ (_10890_, _13051_, _13049_);
  not _21322_ (_13052_, _12700_);
  or _21323_ (_13053_, _12883_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _21324_ (_13054_, _12884_);
  and _21325_ (_13055_, _12973_, _13054_);
  and _21326_ (_13056_, _13055_, _13053_);
  not _21327_ (_13057_, _07496_);
  or _21328_ (_13058_, _12745_, _12701_);
  and _21329_ (_13059_, _13058_, _13057_);
  not _21330_ (_13060_, _07533_);
  and _21331_ (_13061_, _12707_, _13060_);
  and _21332_ (_13062_, _12713_, _12880_);
  and _21333_ (_13063_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _21334_ (_13064_, _13063_, _13062_);
  or _21335_ (_13065_, _13064_, _13061_);
  or _21336_ (_13066_, _13065_, _13059_);
  or _21337_ (_13068_, _13066_, _13056_);
  or _21338_ (_13069_, _13068_, _13052_);
  or _21339_ (_13070_, _12700_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _21340_ (_13071_, _13070_, _05141_);
  and _21341_ (_10936_, _13071_, _13069_);
  nor _21342_ (_10940_, _12498_, rst);
  and _21343_ (_13072_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _21344_ (_13073_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or _21345_ (_13074_, _13073_, _13072_);
  and _21346_ (_10943_, _13074_, _05141_);
  nor _21347_ (_10986_, _12550_, rst);
  nand _21348_ (_13075_, _11418_, _07434_);
  or _21349_ (_13076_, _11418_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _21350_ (_13077_, _13076_, _05141_);
  and _21351_ (_11030_, _13077_, _13075_);
  and _21352_ (_13078_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _21353_ (_13079_, _12091_, _12050_);
  nor _21354_ (_13080_, _13079_, _12092_);
  or _21355_ (_13081_, _13080_, _07135_);
  or _21356_ (_13082_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _21357_ (_13083_, _13082_, _12108_);
  and _21358_ (_13084_, _13083_, _13081_);
  or _21359_ (_11034_, _13084_, _13078_);
  and _21360_ (_13085_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _21361_ (_13086_, _12094_, _12038_);
  nor _21362_ (_13087_, _13086_, _12095_);
  or _21363_ (_13088_, _13087_, _07135_);
  or _21364_ (_13089_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _21365_ (_13090_, _13089_, _12108_);
  and _21366_ (_13091_, _13090_, _13088_);
  or _21367_ (_11063_, _13091_, _13085_);
  nor _21368_ (_13092_, _12093_, _12042_);
  nor _21369_ (_13093_, _13092_, _12094_);
  or _21370_ (_13094_, _13093_, _07135_);
  or _21371_ (_13095_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _21372_ (_13096_, _13095_, _12108_);
  and _21373_ (_13097_, _13096_, _13094_);
  and _21374_ (_13098_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _21375_ (_11068_, _13098_, _13097_);
  and _21376_ (_13099_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _21377_ (_13100_, _12092_, _12046_);
  nor _21378_ (_13101_, _13100_, _12093_);
  or _21379_ (_13102_, _13101_, _07135_);
  or _21380_ (_13103_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _21381_ (_13104_, _13103_, _12108_);
  and _21382_ (_13105_, _13104_, _13102_);
  or _21383_ (_11077_, _13105_, _13099_);
  or _21384_ (_13106_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand _21385_ (_13107_, _07619_, _06353_);
  and _21386_ (_13108_, _13107_, _05141_);
  and _21387_ (_11094_, _13108_, _13106_);
  and _21388_ (_13109_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _21389_ (_13110_, _07619_, _06379_);
  or _21390_ (_13111_, _13110_, _13109_);
  and _21391_ (_11098_, _13111_, _05141_);
  and _21392_ (_13112_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor _21393_ (_13113_, _07619_, _06459_);
  or _21394_ (_13114_, _13113_, _13112_);
  and _21395_ (_11100_, _13114_, _05141_);
  and _21396_ (_13115_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not _21397_ (_13116_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _21398_ (_13117_, pc_log_change, _13116_);
  or _21399_ (_13118_, _13117_, _13115_);
  and _21400_ (_11104_, _13118_, _05141_);
  and _21401_ (_13119_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _21402_ (_13120_, _07619_, _06376_);
  or _21403_ (_13121_, _13120_, _13119_);
  and _21404_ (_11107_, _13121_, _05141_);
  or _21405_ (_13122_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _21406_ (_13123_, _07619_, _06306_);
  and _21407_ (_13124_, _13123_, _05141_);
  and _21408_ (_11161_, _13124_, _13122_);
  or _21409_ (_13125_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand _21410_ (_13126_, _07619_, _06516_);
  and _21411_ (_13127_, _13126_, _05141_);
  and _21412_ (_11163_, _13127_, _13125_);
  or _21413_ (_13128_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _21414_ (_13129_, _07619_, _06484_);
  and _21415_ (_13130_, _13129_, _05141_);
  and _21416_ (_11166_, _13130_, _13128_);
  or _21417_ (_13131_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not _21418_ (_13132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _21419_ (_13133_, _06728_, _13132_);
  and _21420_ (_13134_, _13133_, _13131_);
  or _21421_ (_13135_, _13134_, _06738_);
  nand _21422_ (_13136_, _06738_, _05604_);
  and _21423_ (_13137_, _13136_, _13135_);
  or _21424_ (_13138_, _13137_, _06743_);
  nand _21425_ (_13139_, _06743_, _08441_);
  and _21426_ (_13140_, _13139_, _05141_);
  and _21427_ (_11180_, _13140_, _13138_);
  or _21428_ (_13141_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _21429_ (_13142_, _07619_, _06311_);
  and _21430_ (_13143_, _13142_, _05141_);
  and _21431_ (_11214_, _13143_, _13141_);
  and _21432_ (_13144_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _21433_ (_13145_, _07619_, _06399_);
  or _21434_ (_13146_, _13145_, _13144_);
  and _21435_ (_11217_, _13146_, _05141_);
  and _21436_ (_13147_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _21437_ (_13148_, _07619_, _06403_);
  or _21438_ (_13149_, _13148_, _13147_);
  and _21439_ (_11221_, _13149_, _05141_);
  and _21440_ (_11229_, _11737_, _05141_);
  or _21441_ (_13150_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand _21442_ (_13151_, _07619_, _06374_);
  and _21443_ (_13152_, _13151_, _05141_);
  and _21444_ (_11236_, _13152_, _13150_);
  or _21445_ (_13153_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not _21446_ (_13154_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _21447_ (_13155_, pc_log_change, _13154_);
  and _21448_ (_13156_, _13155_, _05141_);
  and _21449_ (_11239_, _13156_, _13153_);
  and _21450_ (_13157_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _21451_ (_13158_, _13157_, _11815_);
  not _21452_ (_13159_, _08439_);
  nor _21453_ (_13160_, _11811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _21454_ (_13161_, _13160_, _11812_);
  or _21455_ (_13162_, _13161_, _13159_);
  or _21456_ (_13163_, _13162_, _13158_);
  or _21457_ (_13164_, _08439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _21458_ (_13165_, _13164_, _13163_);
  or _21459_ (_13166_, _13165_, _08463_);
  nor _21460_ (_13167_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _21461_ (_13168_, _13167_, _08471_);
  and _21462_ (_13169_, _13168_, _13166_);
  and _21463_ (_13170_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _21464_ (_13171_, _13170_, _08478_);
  or _21465_ (_13172_, _13171_, _13169_);
  or _21466_ (_13173_, _11789_, _05522_);
  and _21467_ (_13175_, _13173_, _05141_);
  and _21468_ (_11254_, _13175_, _13172_);
  or _21469_ (_13176_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand _21470_ (_13177_, _07619_, _06370_);
  and _21471_ (_13178_, _13177_, _05141_);
  and _21472_ (_11259_, _13178_, _13176_);
  and _21473_ (_13179_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _21474_ (_13180_, _07619_, _06427_);
  or _21475_ (_13181_, _13180_, _13179_);
  and _21476_ (_11263_, _13181_, _05141_);
  or _21477_ (_13182_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand _21478_ (_13183_, _07619_, _06510_);
  and _21479_ (_13184_, _13183_, _05141_);
  and _21480_ (_11281_, _13184_, _13182_);
  nand _21481_ (_13185_, _11418_, _06617_);
  or _21482_ (_13186_, _11418_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _21483_ (_13187_, _13186_, _05141_);
  and _21484_ (_11300_, _13187_, _13185_);
  or _21485_ (_13188_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand _21486_ (_13189_, _07619_, _06406_);
  and _21487_ (_13190_, _13189_, _05141_);
  and _21488_ (_11310_, _13190_, _13188_);
  and _21489_ (_13191_, _07611_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _21490_ (_13192_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [3]);
  or _21491_ (_13193_, _13192_, _13191_);
  and _21492_ (_11319_, _13193_, _05141_);
  and _21493_ (_13194_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _07611_);
  and _21494_ (_13195_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21495_ (_13196_, _13195_, _13194_);
  and _21496_ (_11323_, _13196_, _05141_);
  and _21497_ (_13197_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07611_);
  and _21498_ (_13198_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21499_ (_13199_, _13198_, _13197_);
  and _21500_ (_11335_, _13199_, _05141_);
  and _21501_ (_13200_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07611_);
  and _21502_ (_13201_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21503_ (_13202_, _13201_, _13200_);
  and _21504_ (_11346_, _13202_, _05141_);
  or _21505_ (_13203_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand _21506_ (_13204_, _07619_, _06429_);
  and _21507_ (_13206_, _13204_, _05141_);
  and _21508_ (_11356_, _13206_, _13203_);
  and _21509_ (_13208_, _06290_, _05617_);
  and _21510_ (_13209_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or _21511_ (_13210_, _13209_, _13208_);
  and _21512_ (_11360_, _13210_, _05141_);
  or _21513_ (_13211_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand _21514_ (_13212_, _07619_, _06395_);
  and _21515_ (_13213_, _13212_, _05141_);
  and _21516_ (_11363_, _13213_, _13211_);
  or _21517_ (_13214_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand _21518_ (_13215_, _07619_, _06489_);
  and _21519_ (_13216_, _13215_, _05141_);
  and _21520_ (_11376_, _13216_, _13214_);
  or _21521_ (_13217_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand _21522_ (_13218_, _07619_, _06438_);
  and _21523_ (_13219_, _13218_, _05141_);
  and _21524_ (_11389_, _13219_, _13217_);
  or _21525_ (_13220_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand _21526_ (_13221_, _07619_, _06343_);
  and _21527_ (_13222_, _13221_, _05141_);
  and _21528_ (_11409_, _13222_, _13220_);
  or _21529_ (_13223_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _21530_ (_13224_, _07619_, _06464_);
  and _21531_ (_13225_, _13224_, _05141_);
  and _21532_ (_11416_, _13225_, _13223_);
  and _21533_ (_11515_, _11745_, _05141_);
  nor _21534_ (_11523_, _11742_, rst);
  nand _21535_ (_13226_, _08305_, _05560_);
  or _21536_ (_13227_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _21537_ (_13228_, _13227_, _05141_);
  and _21538_ (_11526_, _13228_, _13226_);
  nor _21539_ (_13229_, _11619_, _11617_);
  nor _21540_ (_13230_, _13229_, _11620_);
  or _21541_ (_13231_, _13230_, _07516_);
  or _21542_ (_13232_, _06271_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _21543_ (_13233_, _13232_, _12108_);
  and _21544_ (_11616_, _13233_, _13231_);
  and _21545_ (_13234_, _11615_, _06271_);
  nand _21546_ (_13235_, _13234_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _21547_ (_13236_, _13234_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _21548_ (_13237_, _13236_, _12108_);
  and _21549_ (_11632_, _13237_, _13235_);
  or _21550_ (_13238_, _11477_, _07011_);
  and _21551_ (_13239_, _06524_, _06497_);
  and _21552_ (_13240_, _13239_, _07014_);
  or _21553_ (_13241_, _13240_, _11501_);
  and _21554_ (_13242_, _13241_, _13238_);
  not _21555_ (_13243_, _11546_);
  or _21556_ (_13244_, _13243_, _07029_);
  or _21557_ (_13245_, _13244_, _13242_);
  and _21558_ (_13246_, _11511_, _07012_);
  nor _21559_ (_13247_, _11596_, _11478_);
  or _21560_ (_13248_, _13247_, _07013_);
  or _21561_ (_13249_, _13248_, _13246_);
  and _21562_ (_13250_, _11477_, _11549_);
  and _21563_ (_13251_, _11543_, _07009_);
  or _21564_ (_13252_, _11609_, _13251_);
  or _21565_ (_13253_, _13252_, _13250_);
  or _21566_ (_13254_, _11504_, _11585_);
  or _21567_ (_13255_, _11564_, _11548_);
  or _21568_ (_13256_, _13255_, _13254_);
  or _21569_ (_13257_, _13256_, _13253_);
  or _21570_ (_13258_, _13257_, _13249_);
  or _21571_ (_13259_, _13258_, _13245_);
  and _21572_ (_13261_, _13259_, _06272_);
  nor _21573_ (_13262_, _07005_, _06790_);
  or _21574_ (_13263_, _13262_, rst);
  or _21575_ (_11638_, _13263_, _13261_);
  and _21576_ (_13264_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _21577_ (_13265_, _07619_, _06301_);
  or _21578_ (_13266_, _13265_, _13264_);
  and _21579_ (_11641_, _13266_, _05141_);
  and _21580_ (_13267_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor _21581_ (_13268_, _07619_, _06351_);
  or _21582_ (_13269_, _13268_, _13267_);
  and _21583_ (_11645_, _13269_, _05141_);
  nand _21584_ (_13270_, _06832_, _06449_);
  and _21585_ (_13271_, _13270_, _06830_);
  or _21586_ (_13272_, _06541_, _06831_);
  or _21587_ (_11658_, _13272_, _13271_);
  and _21588_ (_13273_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _21589_ (_13274_, _07619_, _06514_);
  or _21590_ (_13275_, _13274_, _13273_);
  and _21591_ (_11664_, _13275_, _05141_);
  and _21592_ (_13276_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _21593_ (_13277_, _07619_, _06487_);
  or _21594_ (_13278_, _13277_, _13276_);
  and _21595_ (_11666_, _13278_, _05141_);
  and _21596_ (_13279_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _21597_ (_13280_, _07619_, _06324_);
  or _21598_ (_13281_, _13280_, _13279_);
  and _21599_ (_11670_, _13281_, _05141_);
  and _21600_ (_13282_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _21601_ (_13283_, _07619_, _06347_);
  or _21602_ (_13284_, _13283_, _13282_);
  and _21603_ (_11675_, _13284_, _05141_);
  nand _21604_ (_13285_, _06472_, _06270_);
  or _21605_ (_13286_, _06270_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _21606_ (_13287_, _13286_, _05141_);
  and _21607_ (_11677_, _13287_, _13285_);
  and _21608_ (_13288_, _06755_, _06547_);
  or _21609_ (_13289_, _13288_, _07060_);
  or _21610_ (_13290_, _13289_, _06785_);
  and _21611_ (_13291_, _13290_, _06296_);
  and _21612_ (_13292_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _21613_ (_13293_, _13292_, _06798_);
  and _21614_ (_13294_, _13293_, _05141_);
  or _21615_ (_11679_, _13294_, _13291_);
  and _21616_ (_13295_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _21617_ (_13296_, _07619_, _06482_);
  or _21618_ (_13297_, _13296_, _13295_);
  and _21619_ (_11682_, _13297_, _05141_);
  or _21620_ (_13298_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand _21621_ (_13299_, _07619_, _06434_);
  and _21622_ (_13300_, _13299_, _05141_);
  and _21623_ (_11688_, _13300_, _13298_);
  and _21624_ (_13301_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _21625_ (_13302_, _07619_, _06457_);
  or _21626_ (_13303_, _13302_, _13301_);
  and _21627_ (_11695_, _13303_, _05141_);
  and _21628_ (_11697_, _11454_, _05141_);
  nand _21629_ (_13304_, _08305_, _06178_);
  or _21630_ (_13305_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _21631_ (_13306_, _13305_, _05141_);
  and _21632_ (_11700_, _13306_, _13304_);
  and _21633_ (_13307_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _21634_ (_13308_, _07619_, _06508_);
  or _21635_ (_13309_, _13308_, _13307_);
  and _21636_ (_11703_, _13309_, _05141_);
  or _21637_ (_13310_, _08306_, _05522_);
  or _21638_ (_13311_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _21639_ (_13312_, _13311_, _05141_);
  and _21640_ (_11717_, _13312_, _13310_);
  and _21641_ (_11719_, _12158_, _05141_);
  nand _21642_ (_13313_, _06707_, _06062_);
  or _21643_ (_13314_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _21644_ (_13315_, _13314_, _05141_);
  and _21645_ (_11890_, _13315_, _13313_);
  nand _21646_ (_13316_, _11418_, _07496_);
  or _21647_ (_13317_, _11418_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _21648_ (_13318_, _13317_, _05141_);
  and _21649_ (_11921_, _13318_, _13316_);
  nand _21650_ (_13319_, _11418_, _07350_);
  or _21651_ (_13320_, _11418_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _21652_ (_13321_, _13320_, _05141_);
  and _21653_ (_11947_, _13321_, _13319_);
  and _21654_ (_13322_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _21655_ (_13323_, _13322_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _21656_ (_11968_, _13323_, _05141_);
  and _21657_ (_13324_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _21658_ (_13325_, _13324_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _21659_ (_11975_, _13325_, _05141_);
  or _21660_ (_13326_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _21661_ (_13327_, _07619_, _06351_);
  and _21662_ (_13328_, _13327_, _05141_);
  and _21663_ (_11979_, _13328_, _13326_);
  or _21664_ (_13329_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand _21665_ (_13330_, _07619_, _06482_);
  and _21666_ (_13331_, _13330_, _05141_);
  and _21667_ (_11987_, _13331_, _13329_);
  and _21668_ (_13333_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _21669_ (_13334_, _13333_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _21670_ (_11993_, _13334_, _05141_);
  or _21671_ (_13335_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _21672_ (_13336_, _07619_, _06459_);
  and _21673_ (_13337_, _13336_, _05141_);
  and _21674_ (_11995_, _13337_, _13335_);
  and _21675_ (_13338_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _21676_ (_13339_, _13338_, _10356_);
  and _21677_ (_13340_, _13339_, _11458_);
  nand _21678_ (_13341_, _11458_, _08283_);
  and _21679_ (_13342_, _13341_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _21680_ (_13343_, _13342_, _11462_);
  or _21681_ (_13344_, _13343_, _13340_);
  nand _21682_ (_13345_, _11462_, _05560_);
  and _21683_ (_13346_, _13345_, _05141_);
  and _21684_ (_12002_, _13346_, _13344_);
  and _21685_ (_13347_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _21686_ (_13348_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or _21687_ (_13349_, _13348_, _13347_);
  and _21688_ (_12008_, _13349_, _05141_);
  and _21689_ (_13350_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _05141_);
  and _21690_ (_13351_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _05141_);
  and _21691_ (_13353_, _13351_, _11643_);
  or _21692_ (_12013_, _13353_, _13350_);
  and _21693_ (_13354_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _21694_ (_13355_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or _21695_ (_13356_, _13355_, _13354_);
  and _21696_ (_12016_, _13356_, _05141_);
  and _21697_ (_13357_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _21698_ (_13358_, _13357_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _21699_ (_12018_, _13358_, _05141_);
  or _21700_ (_13359_, _06745_, _06004_);
  and _21701_ (_13360_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _21702_ (_13361_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _21703_ (_13362_, _13361_, _13360_);
  or _21704_ (_13363_, _13362_, _06743_);
  and _21705_ (_13364_, _13363_, _05141_);
  and _21706_ (_12058_, _13364_, _13359_);
  and _21707_ (_13365_, _06742_, _05649_);
  not _21708_ (_13366_, _13365_);
  or _21709_ (_13368_, _13366_, _06004_);
  not _21710_ (_13369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _21711_ (_13370_, _13369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _21712_ (_13371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _21713_ (_13372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13371_);
  nor _21714_ (_13373_, _13372_, _13370_);
  not _21715_ (_13374_, _13373_);
  nand _21716_ (_13375_, _08476_, _05649_);
  and _21717_ (_13376_, _13375_, _13374_);
  not _21718_ (_13377_, _13376_);
  and _21719_ (_13378_, _13377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  not _21720_ (_13379_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _21721_ (_13381_, _13379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not _21722_ (_13382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _21723_ (_13383_, \oc8051_top_1.oc8051_sfr1.pres_ow , _13382_);
  not _21724_ (_13384_, t1_i);
  and _21725_ (_13385_, _13384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _21726_ (_13386_, _13385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or _21727_ (_13388_, _13386_, _13383_);
  and _21728_ (_13389_, _13388_, _13381_);
  and _21729_ (_13391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _21730_ (_13392_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _21731_ (_13393_, _13392_, _13391_);
  and _21732_ (_13394_, _13393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _21733_ (_13395_, _13394_, _13389_);
  nor _21734_ (_13396_, _13395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _21735_ (_13397_, _13395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _21736_ (_13398_, _13397_, _13396_);
  and _21737_ (_13399_, _13374_, _13398_);
  and _21738_ (_13400_, _13397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _21739_ (_13401_, _13400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _21740_ (_13402_, _13401_, _13370_);
  and _21741_ (_13403_, _13402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _21742_ (_13404_, _13403_, _13399_);
  and _21743_ (_13405_, _13404_, _13375_);
  or _21744_ (_13406_, _13405_, _13378_);
  or _21745_ (_13407_, _13365_, _13406_);
  and _21746_ (_13408_, _13407_, _05141_);
  and _21747_ (_12067_, _13408_, _13368_);
  and _21748_ (_13409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _21749_ (_13410_, _13409_);
  and _21750_ (_13412_, _13410_, _13375_);
  and _21751_ (_13413_, _13393_, _13389_);
  and _21752_ (_13414_, _13413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _21753_ (_13415_, _13413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _21754_ (_13416_, _13415_, _13414_);
  and _21755_ (_13417_, _13416_, _13412_);
  not _21756_ (_13418_, _13412_);
  and _21757_ (_13419_, _13418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _21758_ (_13420_, _13419_, _13417_);
  and _21759_ (_13421_, _13402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _21760_ (_13422_, _13421_, _13375_);
  or _21761_ (_13423_, _13422_, _13365_);
  or _21762_ (_13424_, _13423_, _13420_);
  or _21763_ (_13425_, _13366_, _05522_);
  and _21764_ (_13426_, _13425_, _05141_);
  and _21765_ (_12070_, _13426_, _13424_);
  and _21766_ (_13427_, _13389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _21767_ (_13428_, _13427_, _13391_);
  nor _21768_ (_13429_, _13428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _21769_ (_13430_, _13429_, _13413_);
  nand _21770_ (_13432_, _13430_, _13412_);
  or _21771_ (_13433_, _13412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _21772_ (_13434_, _13433_, _13432_);
  and _21773_ (_13435_, _05649_, _05173_);
  and _21774_ (_13437_, _13435_, _06032_);
  and _21775_ (_13438_, _13437_, _05925_);
  and _21776_ (_13439_, _05965_, _05925_);
  and _21777_ (_13440_, _13414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _21778_ (_13441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _21779_ (_13442_, _13441_, _13440_);
  and _21780_ (_13443_, _13442_, _13370_);
  nand _21781_ (_13444_, _13443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _21782_ (_13445_, _13444_, _13439_);
  or _21783_ (_13446_, _13445_, _13438_);
  or _21784_ (_13447_, _13446_, _13434_);
  nand _21785_ (_13448_, _13438_, _06062_);
  and _21786_ (_13449_, _13448_, _05141_);
  and _21787_ (_12073_, _13449_, _13447_);
  nor _21788_ (_12076_, _12287_, rst);
  nand _21789_ (_13450_, _13365_, _06244_);
  nor _21790_ (_13451_, _13397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _21791_ (_13452_, _13451_, _13400_);
  and _21792_ (_13453_, _13452_, _13376_);
  and _21793_ (_13454_, _13377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _21794_ (_13455_, _13443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _21795_ (_13456_, _13455_, _13439_);
  or _21796_ (_13457_, _13456_, _13454_);
  or _21797_ (_13458_, _13457_, _13453_);
  or _21798_ (_13459_, _13458_, _13365_);
  and _21799_ (_13460_, _13459_, _05141_);
  and _21800_ (_12080_, _13460_, _13450_);
  nor _21801_ (_12082_, _12425_, rst);
  nand _21802_ (_13461_, _08305_, _06062_);
  or _21803_ (_13462_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _21804_ (_13463_, _13462_, _05141_);
  and _21805_ (_12085_, _13463_, _13461_);
  not _21806_ (_13464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _21807_ (_13465_, _13412_, _13464_);
  or _21808_ (_13466_, _13389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _21809_ (_13467_, _13427_, _13409_);
  and _21810_ (_13468_, _13467_, _13466_);
  and _21811_ (_13469_, _13370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _21812_ (_13470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _21813_ (_13471_, _13470_, _13441_);
  and _21814_ (_13472_, _13471_, _13393_);
  and _21815_ (_13473_, _13472_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _21816_ (_13474_, _13473_, _13469_);
  or _21817_ (_00003_, _13474_, _13468_);
  and _21818_ (_00004_, _00003_, _13375_);
  or _21819_ (_00005_, _00004_, _13365_);
  or _21820_ (_00006_, _00005_, _13465_);
  nand _21821_ (_00007_, _13365_, _05604_);
  and _21822_ (_00008_, _00007_, _05141_);
  and _21823_ (_12090_, _00008_, _00006_);
  and _21824_ (_00009_, _13427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _21825_ (_00010_, _13427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _21826_ (_00011_, _00010_, _00009_);
  and _21827_ (_00012_, _00011_, _13412_);
  nand _21828_ (_00013_, _13443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _21829_ (_00014_, _00013_, _13439_);
  or _21830_ (_00015_, _00014_, _00012_);
  and _21831_ (_00016_, _13418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _21832_ (_00017_, _00016_, _13365_);
  or _21833_ (_00018_, _00017_, _00015_);
  nand _21834_ (_00019_, _13365_, _06178_);
  and _21835_ (_00020_, _00019_, _05141_);
  and _21836_ (_12098_, _00020_, _00018_);
  nor _21837_ (_00021_, _00009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _21838_ (_00022_, _00021_, _13428_);
  and _21839_ (_00023_, _00022_, _13412_);
  and _21840_ (_00024_, _13418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _21841_ (_00025_, _00024_, _00023_);
  and _21842_ (_00026_, _13402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21843_ (_00027_, _00026_, _13375_);
  or _21844_ (_00028_, _00027_, _13365_);
  or _21845_ (_00029_, _00028_, _00025_);
  nand _21846_ (_00030_, _13365_, _05560_);
  and _21847_ (_00031_, _00030_, _05141_);
  and _21848_ (_12102_, _00031_, _00029_);
  nor _21849_ (_12104_, _12186_, rst);
  nor _21850_ (_12109_, _12796_, rst);
  nor _21851_ (_12113_, _12368_, rst);
  nor _21852_ (_12116_, _12604_, rst);
  or _21853_ (_00032_, _13375_, _06179_);
  not _21854_ (_00033_, _13372_);
  and _21855_ (_00034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _21856_ (_00035_, _13441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _21857_ (_00036_, _00035_, _00034_);
  and _21858_ (_00037_, _00036_, _13393_);
  and _21859_ (_00038_, _00037_, _13389_);
  nor _21860_ (_00039_, _00038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _21861_ (_00040_, _13473_, _13389_);
  and _21862_ (_00041_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _21863_ (_00042_, _00041_, _00039_);
  or _21864_ (_00043_, _00042_, _00033_);
  and _21865_ (_00044_, _00034_, _13393_);
  and _21866_ (_00045_, _00044_, _13389_);
  nor _21867_ (_00046_, _00045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _21868_ (_00047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _21869_ (_00048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _21870_ (_00049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _21871_ (_00050_, _00049_, _13414_);
  nand _21872_ (_00051_, _00050_, _00048_);
  and _21873_ (_00052_, _00051_, _00047_);
  or _21874_ (_00053_, _00052_, _00046_);
  and _21875_ (_00054_, _00053_, _00043_);
  nand _21876_ (_00055_, _00054_, _13375_);
  and _21877_ (_00056_, _00055_, _13366_);
  and _21878_ (_00057_, _00056_, _00032_);
  and _21879_ (_00058_, _13438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _21880_ (_00059_, _00058_, _00057_);
  and _21881_ (_12119_, _00059_, _05141_);
  not _21882_ (_00060_, _13438_);
  and _21883_ (_00061_, _13439_, _05560_);
  or _21884_ (_00062_, _00041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21885_ (_00063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21886_ (_00064_, _00063_, _00040_);
  nor _21887_ (_00065_, _00064_, _00033_);
  nand _21888_ (_00066_, _00065_, _00062_);
  nor _21889_ (_00067_, _00050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _21890_ (_00068_, _00067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21891_ (_00069_, _00034_, _13413_);
  and _21892_ (_00070_, _00063_, _13371_);
  and _21893_ (_00071_, _00070_, _00069_);
  nor _21894_ (_00072_, _00071_, _13372_);
  nand _21895_ (_00073_, _00072_, _00068_);
  and _21896_ (_00074_, _00073_, _00066_);
  and _21897_ (_00075_, _00074_, _13375_);
  or _21898_ (_00076_, _00075_, _00061_);
  nand _21899_ (_00077_, _00076_, _00060_);
  or _21900_ (_00078_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21901_ (_00079_, _00078_, _05141_);
  and _21902_ (_12122_, _00079_, _00077_);
  not _21903_ (_00080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _21904_ (_00081_, _00048_, _13414_);
  and _21905_ (_00082_, _13442_, _13372_);
  nor _21906_ (_00083_, _00082_, _00081_);
  nand _21907_ (_00084_, _00083_, _00080_);
  or _21908_ (_00085_, _00083_, _00080_);
  nand _21909_ (_00086_, _00085_, _00084_);
  nor _21910_ (_00087_, _00086_, _13439_);
  and _21911_ (_00088_, _13439_, _06703_);
  or _21912_ (_00089_, _00088_, _00087_);
  or _21913_ (_00090_, _00089_, _13365_);
  nand _21914_ (_00091_, _13365_, _00080_);
  and _21915_ (_00092_, _00091_, _05141_);
  and _21916_ (_12125_, _00092_, _00090_);
  and _21917_ (_00093_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _21918_ (_00094_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _21919_ (_00095_, _00094_, _00093_);
  or _21920_ (_00096_, _00095_, _06743_);
  nand _21921_ (_00097_, _06743_, _05560_);
  and _21922_ (_00098_, _00097_, _05141_);
  and _21923_ (_12128_, _00098_, _00096_);
  or _21924_ (_00099_, _13375_, _05522_);
  nand _21925_ (_00100_, _00071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _21926_ (_00101_, _00100_, _00033_);
  and _21927_ (_00102_, _00063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _21928_ (_00103_, _00102_, _00038_);
  nor _21929_ (_00104_, _00103_, _00033_);
  nor _21930_ (_00105_, _00104_, _00101_);
  or _21931_ (_00106_, _00105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _21932_ (_00107_, _00105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _21933_ (_00108_, _00107_, _00106_);
  and _21934_ (_00109_, _00108_, _13375_);
  nor _21935_ (_00110_, _00109_, _13365_);
  and _21936_ (_00111_, _00110_, _00099_);
  and _21937_ (_00112_, _06034_, _05925_);
  and _21938_ (_00113_, _00112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _21939_ (_00114_, _00113_, _00111_);
  and _21940_ (_12134_, _00114_, _05141_);
  and _21941_ (_00115_, _13439_, _06244_);
  not _21942_ (_00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _21943_ (_00117_, _00107_, _00116_);
  and _21944_ (_00118_, _00117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _21945_ (_00119_, _00117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _21946_ (_00120_, _00119_, _00118_);
  nor _21947_ (_00121_, _00120_, _13439_);
  or _21948_ (_00122_, _00121_, _00115_);
  nand _21949_ (_00123_, _00122_, _00060_);
  or _21950_ (_00124_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _21951_ (_00125_, _00124_, _05141_);
  and _21952_ (_12137_, _00125_, _00123_);
  or _21953_ (_00126_, _13375_, _06004_);
  nand _21954_ (_00127_, _00107_, _00116_);
  and _21955_ (_00128_, _00127_, _00117_);
  nor _21956_ (_00129_, _00128_, _13439_);
  nor _21957_ (_00130_, _00129_, _13365_);
  and _21958_ (_00131_, _00130_, _00126_);
  and _21959_ (_00132_, _00112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _21960_ (_00133_, _00132_, _00131_);
  and _21961_ (_12140_, _00133_, _05141_);
  and _21962_ (_00134_, _13439_, _06062_);
  nor _21963_ (_00135_, _00072_, _00065_);
  not _21964_ (_00136_, _00135_);
  nand _21965_ (_00137_, _00136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _21966_ (_00138_, _00136_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _21967_ (_00139_, _00138_, _00137_);
  and _21968_ (_00140_, _00139_, _13375_);
  or _21969_ (_00141_, _00140_, _00134_);
  nand _21970_ (_00142_, _00141_, _00060_);
  or _21971_ (_00143_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _21972_ (_00144_, _00143_, _05141_);
  and _21973_ (_12143_, _00144_, _00142_);
  or _21974_ (_00145_, _12912_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _21975_ (_00146_, _00145_, _12913_);
  or _21976_ (_00148_, _00146_, _12773_);
  nand _21977_ (_00149_, _12904_, _05455_);
  and _21978_ (_00150_, _00149_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _21979_ (_00151_, _00150_, _12969_);
  and _21980_ (_00152_, _00151_, _12973_);
  and _21981_ (_00153_, _00152_, _00148_);
  and _21982_ (_00154_, _12701_, _07319_);
  and _21983_ (_00155_, _12707_, _12843_);
  nor _21984_ (_00156_, _12703_, _07350_);
  or _21985_ (_00157_, _00156_, _00155_);
  or _21986_ (_00159_, _12985_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _21987_ (_00160_, _00159_, _12724_);
  and _21988_ (_00161_, _00160_, _12713_);
  and _21989_ (_00162_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _21990_ (_00163_, _00162_, _00161_);
  or _21991_ (_00164_, _00163_, _00157_);
  nor _21992_ (_00165_, _00164_, _00154_);
  nand _21993_ (_00166_, _00165_, _12700_);
  or _21994_ (_00167_, _00166_, _00153_);
  nor _21995_ (_00168_, _13002_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _21996_ (_00169_, _00168_, _13003_);
  or _21997_ (_00170_, _00169_, _12700_);
  and _21998_ (_00171_, _00170_, _05141_);
  and _21999_ (_12146_, _00171_, _00167_);
  not _22000_ (_00173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _22001_ (_00174_, t0_i);
  and _22002_ (_00175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00174_);
  nor _22003_ (_00176_, _00175_, _00173_);
  not _22004_ (_00177_, _00176_);
  not _22005_ (_00178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _22006_ (_00179_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _22007_ (_00180_, _00179_, _00178_);
  and _22008_ (_00181_, _00180_, _00177_);
  and _22009_ (_00182_, _00181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _22010_ (_00183_, _00182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _22011_ (_00184_, _00182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _22012_ (_00185_, _00184_, _00183_);
  not _22013_ (_00186_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22014_ (_00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _00186_);
  and _22015_ (_00188_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22016_ (_00189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _22017_ (_00190_, _00189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _22018_ (_00191_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _22019_ (_00192_, _00191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _22020_ (_00193_, _00192_, _00181_);
  and _22021_ (_00194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _22022_ (_00195_, _00194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _22023_ (_00196_, _00195_, _00193_);
  and _22024_ (_00197_, _00196_, _00188_);
  nor _22025_ (_00198_, _00197_, _00185_);
  and _22026_ (_00199_, _08470_, _05649_);
  nor _22027_ (_00200_, _00199_, _00198_);
  and _22028_ (_00201_, _00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _22029_ (_00202_, _00201_, _00200_);
  and _22030_ (_00203_, _06737_, _05649_);
  not _22031_ (_00204_, _00203_);
  and _22032_ (_00205_, _00204_, _00202_);
  nor _22033_ (_00206_, _00204_, _06178_);
  or _22034_ (_00207_, _00206_, _00205_);
  and _22035_ (_12154_, _00207_, _05141_);
  not _22036_ (_00208_, _12796_);
  and _22037_ (_00210_, _00208_, _12707_);
  and _22038_ (_00211_, _13058_, _06669_);
  and _22039_ (_00212_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _22040_ (_00213_, _12713_, _12776_);
  or _22041_ (_00214_, _00213_, _00212_);
  or _22042_ (_00215_, _00214_, _00211_);
  and _22043_ (_00216_, _12899_, _12896_);
  or _22044_ (_00217_, _00216_, _12840_);
  or _22045_ (_00218_, _00217_, _12806_);
  and _22046_ (_00219_, _00217_, _12806_);
  not _22047_ (_00220_, _00219_);
  and _22048_ (_00221_, _00220_, _12940_);
  and _22049_ (_00222_, _00221_, _00218_);
  or _22050_ (_00223_, _00222_, _00215_);
  or _22051_ (_00224_, _00223_, _00210_);
  and _22052_ (_00225_, _00224_, _12700_);
  and _22053_ (_00226_, _07622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _22054_ (_00227_, _00226_, _12943_);
  and _22055_ (_00228_, _00226_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _22056_ (_00229_, _00228_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _22057_ (_00230_, _00229_, _00227_);
  nor _22058_ (_00231_, _00230_, _12700_);
  or _22059_ (_00232_, _00231_, _00225_);
  and _22060_ (_12157_, _00232_, _05141_);
  not _22061_ (_00233_, _00181_);
  nor _22062_ (_00234_, _00199_, _00233_);
  or _22063_ (_00235_, _00234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _22064_ (_00236_, _00195_, _00192_);
  and _22065_ (_00237_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _22066_ (_00238_, _00237_, _00236_);
  nand _22067_ (_00239_, _00238_, _00182_);
  or _22068_ (_00240_, _00239_, _00199_);
  and _22069_ (_00241_, _00240_, _00235_);
  or _22070_ (_00242_, _00241_, _00203_);
  nand _22071_ (_00243_, _00203_, _05604_);
  and _22072_ (_00244_, _00243_, _05141_);
  and _22073_ (_12160_, _00244_, _00242_);
  or _22074_ (_00245_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _22075_ (_00246_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _22076_ (_00247_, _00246_, _00245_);
  or _22077_ (_00248_, _00247_, _06743_);
  nand _22078_ (_00249_, _06743_, _06178_);
  and _22079_ (_00250_, _00249_, _05141_);
  and _22080_ (_12163_, _00250_, _00248_);
  and _22081_ (_00251_, _00190_, _00181_);
  nor _22082_ (_00252_, _00184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _22083_ (_00253_, _00252_, _00251_);
  and _22084_ (_00254_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22085_ (_00255_, _00254_, _00196_);
  nor _22086_ (_00256_, _00255_, _00253_);
  nor _22087_ (_00257_, _00256_, _00199_);
  and _22088_ (_00258_, _00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _22089_ (_00259_, _00258_, _00257_);
  and _22090_ (_00260_, _00259_, _00204_);
  nor _22091_ (_00261_, _00204_, _05560_);
  or _22092_ (_00262_, _00261_, _00260_);
  and _22093_ (_12180_, _00262_, _05141_);
  or _22094_ (_00263_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not _22095_ (_00264_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _22096_ (_00265_, _08417_, _00264_);
  and _22097_ (_00266_, _00265_, _00263_);
  or _22098_ (_00267_, _00266_, _06743_);
  nand _22099_ (_00268_, _06743_, _05604_);
  and _22100_ (_00269_, _00268_, _05141_);
  and _22101_ (_12183_, _00269_, _00267_);
  and _22102_ (_00270_, _00251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _22103_ (_00271_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _22104_ (_00272_, _00271_, _00193_);
  and _22105_ (_00273_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22106_ (_00274_, _00273_, _00196_);
  nor _22107_ (_00275_, _00274_, _00272_);
  nor _22108_ (_00276_, _00275_, _00199_);
  and _22109_ (_00277_, _00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _22110_ (_00278_, _00277_, _00276_);
  and _22111_ (_00279_, _00278_, _00204_);
  and _22112_ (_00280_, _00203_, _05522_);
  or _22113_ (_00281_, _00280_, _00279_);
  and _22114_ (_12187_, _00281_, _05141_);
  nor _22115_ (_00282_, _00251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _22116_ (_00283_, _00282_, _00270_);
  and _22117_ (_00284_, _00187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22118_ (_00285_, _00284_, _00196_);
  nor _22119_ (_00286_, _00285_, _00283_);
  nor _22120_ (_00287_, _00286_, _00199_);
  and _22121_ (_00288_, _00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _22122_ (_00289_, _00288_, _00287_);
  and _22123_ (_00290_, _00289_, _00204_);
  nor _22124_ (_00291_, _00204_, _06062_);
  or _22125_ (_00292_, _00291_, _00290_);
  and _22126_ (_12190_, _00292_, _05141_);
  or _22127_ (_00293_, _08345_, _06004_);
  and _22128_ (_00294_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _22129_ (_00295_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _22130_ (_00296_, _00295_, _00294_);
  or _22131_ (_00297_, _00296_, _06738_);
  and _22132_ (_00298_, _00297_, _06745_);
  and _22133_ (_00299_, _00298_, _00293_);
  and _22134_ (_00300_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _22135_ (_00301_, _00300_, _00299_);
  and _22136_ (_12198_, _00301_, _05141_);
  or _22137_ (_00303_, _08345_, _05522_);
  and _22138_ (_00304_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _22139_ (_00305_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _22140_ (_00306_, _00305_, _00304_);
  or _22141_ (_00307_, _00306_, _06738_);
  and _22142_ (_00308_, _00307_, _06745_);
  and _22143_ (_00309_, _00308_, _00303_);
  and _22144_ (_00310_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _22145_ (_00311_, _00310_, _00309_);
  and _22146_ (_12203_, _00311_, _05141_);
  nand _22147_ (_00312_, _06738_, _06062_);
  and _22148_ (_00313_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _22149_ (_00314_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _22150_ (_00315_, _00314_, _00313_);
  or _22151_ (_00316_, _00315_, _06738_);
  and _22152_ (_00317_, _00316_, _06745_);
  and _22153_ (_00318_, _00317_, _00312_);
  and _22154_ (_00319_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _22155_ (_00320_, _00319_, _00318_);
  and _22156_ (_12206_, _00320_, _05141_);
  nand _22157_ (_00321_, _06738_, _05560_);
  and _22158_ (_00322_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _22159_ (_00323_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _22160_ (_00324_, _00323_, _00322_);
  or _22161_ (_00325_, _00324_, _06738_);
  and _22162_ (_00326_, _00325_, _06745_);
  and _22163_ (_00327_, _00326_, _00321_);
  and _22164_ (_00328_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _22165_ (_00329_, _00328_, _00327_);
  and _22166_ (_12210_, _00329_, _05141_);
  nor _22167_ (_00330_, _12088_, _12060_);
  nor _22168_ (_00331_, _00330_, _12089_);
  or _22169_ (_00332_, _00331_, _07135_);
  or _22170_ (_00333_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _22171_ (_00334_, _00333_, _12108_);
  and _22172_ (_00335_, _00334_, _00332_);
  and _22173_ (_00336_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _22174_ (_12212_, _00336_, _00335_);
  nor _22175_ (_00337_, _12071_, _11615_);
  nor _22176_ (_00338_, _00337_, _12072_);
  or _22177_ (_00339_, _00338_, _07135_);
  or _22178_ (_00340_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _22179_ (_00342_, _00340_, _12108_);
  and _22180_ (_00344_, _00342_, _00339_);
  and _22181_ (_00346_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _22182_ (_12218_, _00346_, _00344_);
  nor _22183_ (_00347_, _12095_, _12034_);
  nor _22184_ (_00348_, _00347_, _12096_);
  or _22185_ (_00350_, _00348_, _07135_);
  or _22186_ (_00351_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _22187_ (_00352_, _00351_, _12108_);
  and _22188_ (_00353_, _00352_, _00350_);
  and _22189_ (_00354_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _22190_ (_12227_, _00354_, _00353_);
  nor _22191_ (_00356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not _22192_ (_00358_, _00356_);
  and _22193_ (_00359_, _00358_, _00193_);
  and _22194_ (_00360_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _22195_ (_00361_, _00360_);
  nor _22196_ (_00362_, _00361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _22197_ (_00363_, _00196_, _00187_);
  and _22198_ (_00364_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _22199_ (_00365_, _00364_, _00362_);
  nor _22200_ (_00367_, _00365_, _00199_);
  or _22201_ (_00368_, _00361_, _00199_);
  and _22202_ (_00369_, _00368_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _22203_ (_00371_, _00369_, _00367_);
  and _22204_ (_00372_, _00371_, _00204_);
  nor _22205_ (_00373_, _00204_, _06244_);
  or _22206_ (_00375_, _00373_, _00372_);
  and _22207_ (_12242_, _00375_, _05141_);
  not _22208_ (_00378_, _00199_);
  or _22209_ (_00380_, _00378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _22210_ (_00381_, _00380_, _00204_);
  and _22211_ (_00382_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _22212_ (_00383_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _22213_ (_00384_, _00383_, _00368_);
  or _22214_ (_00385_, _00384_, _00382_);
  and _22215_ (_00386_, _00385_, _00381_);
  and _22216_ (_00388_, _00203_, _06004_);
  or _22217_ (_00389_, _00388_, _00386_);
  and _22218_ (_12246_, _00389_, _05141_);
  nand _22219_ (_00390_, _00199_, _06244_);
  not _22220_ (_00391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22221_ (_00392_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22222_ (_00393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22223_ (_00394_, _00393_, _00193_);
  and _22224_ (_00395_, _00394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22225_ (_00396_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22226_ (_00397_, _00396_, _00392_);
  nor _22227_ (_00398_, _00397_, _00391_);
  and _22228_ (_00399_, _00397_, _00391_);
  or _22229_ (_00400_, _00399_, _00398_);
  and _22230_ (_00401_, _00400_, _00356_);
  and _22231_ (_00402_, _00393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22232_ (_00403_, _00402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22233_ (_00404_, _00403_, _00392_);
  and _22234_ (_00405_, _00236_, _00181_);
  and _22235_ (_00406_, _00405_, _00404_);
  or _22236_ (_00407_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _22237_ (_00408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22238_ (_00409_, _00408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22239_ (_00410_, _00404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _22240_ (_00411_, _00410_, _00405_);
  and _22241_ (_00412_, _00411_, _00409_);
  and _22242_ (_00413_, _00412_, _00407_);
  and _22243_ (_00414_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _22244_ (_00415_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22245_ (_00416_, _00415_, _00404_);
  nand _22246_ (_00417_, _00416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _22247_ (_00418_, _00416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22248_ (_00419_, _00418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22249_ (_00420_, _00419_, _00417_);
  or _22250_ (_00421_, _00420_, _00413_);
  or _22251_ (_00422_, _00421_, _00401_);
  or _22252_ (_00423_, _00422_, _00199_);
  and _22253_ (_00424_, _00423_, _00204_);
  and _22254_ (_00425_, _00424_, _00390_);
  and _22255_ (_00426_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _22256_ (_00427_, _00426_, _00425_);
  and _22257_ (_12284_, _00427_, _05141_);
  nand _22258_ (_00428_, _00199_, _05560_);
  or _22259_ (_00429_, _00394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _22260_ (_00430_, _00395_, _00358_);
  and _22261_ (_00431_, _00430_, _00429_);
  and _22262_ (_00432_, _00405_, _00393_);
  or _22263_ (_00433_, _00432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _22264_ (_00434_, _00405_, _00402_);
  and _22265_ (_00435_, _00434_, _00409_);
  and _22266_ (_00436_, _00435_, _00433_);
  and _22267_ (_00437_, _00414_, _00402_);
  nand _22268_ (_00438_, _00437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22269_ (_00439_, _00414_, _00393_);
  and _22270_ (_00440_, _00439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _22271_ (_00441_, _00440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22272_ (_00442_, _00441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22273_ (_00443_, _00442_, _00438_);
  or _22274_ (_00444_, _00443_, _00436_);
  or _22275_ (_00445_, _00444_, _00431_);
  or _22276_ (_00446_, _00445_, _00199_);
  and _22277_ (_00447_, _00446_, _00204_);
  and _22278_ (_00448_, _00447_, _00428_);
  and _22279_ (_00449_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _22280_ (_00450_, _00449_, _00448_);
  and _22281_ (_12295_, _00450_, _05141_);
  nand _22282_ (_00451_, _00199_, _06062_);
  and _22283_ (_00452_, _00405_, _00408_);
  and _22284_ (_00453_, _00452_, _00402_);
  nand _22285_ (_00454_, _00453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _22286_ (_00455_, _00409_, _00187_);
  or _22287_ (_00456_, _00453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22288_ (_00458_, _00456_, _00455_);
  and _22289_ (_00459_, _00458_, _00454_);
  or _22290_ (_00460_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _22291_ (_00461_, _00396_, _00358_);
  and _22292_ (_00462_, _00461_, _00460_);
  or _22293_ (_00463_, _00437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22294_ (_00464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22295_ (_00465_, _00414_, _00403_);
  not _22296_ (_00466_, _00465_);
  and _22297_ (_00467_, _00466_, _00464_);
  and _22298_ (_00468_, _00467_, _00463_);
  or _22299_ (_00469_, _00468_, _00462_);
  or _22300_ (_00470_, _00469_, _00459_);
  or _22301_ (_00471_, _00470_, _00199_);
  and _22302_ (_00472_, _00471_, _00204_);
  and _22303_ (_00473_, _00472_, _00451_);
  and _22304_ (_00474_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _22305_ (_00475_, _00474_, _00473_);
  and _22306_ (_12298_, _00475_, _05141_);
  or _22307_ (_00476_, _00378_, _05522_);
  and _22308_ (_00477_, _00403_, _00193_);
  or _22309_ (_00478_, _00477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22310_ (_00479_, _00477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _22311_ (_00480_, _00479_, _00358_);
  and _22312_ (_00481_, _00480_, _00478_);
  and _22313_ (_00482_, _00192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _22314_ (_00483_, _00482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _22315_ (_00484_, _00483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _22316_ (_00485_, _00403_, _00181_);
  and _22317_ (_00487_, _00485_, _00484_);
  and _22318_ (_00488_, _00487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _22319_ (_00489_, _00487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _22320_ (_00490_, _00489_, _00409_);
  nor _22321_ (_00491_, _00490_, _00488_);
  and _22322_ (_00492_, _00415_, _00403_);
  nand _22323_ (_00493_, _00492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _22324_ (_00494_, _00492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22325_ (_00495_, _00494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22326_ (_00496_, _00495_, _00493_);
  or _22327_ (_00497_, _00496_, _00491_);
  or _22328_ (_00498_, _00497_, _00481_);
  or _22329_ (_00499_, _00498_, _00199_);
  and _22330_ (_00500_, _00499_, _00204_);
  and _22331_ (_00501_, _00500_, _00476_);
  and _22332_ (_00502_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _22333_ (_00503_, _00502_, _00501_);
  and _22334_ (_12307_, _00503_, _05141_);
  or _22335_ (_00504_, _00378_, _06004_);
  and _22336_ (_00505_, _00488_, _00408_);
  nor _22337_ (_00506_, _00505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22338_ (_00507_, _00505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _22339_ (_00508_, _00507_, _00506_);
  and _22340_ (_00509_, _00508_, _00455_);
  and _22341_ (_00510_, _00465_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _22342_ (_00511_, _00510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _22343_ (_00512_, _00510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22344_ (_00513_, _00512_, _00511_);
  and _22345_ (_00514_, _00513_, _00464_);
  or _22346_ (_00515_, _00479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _22347_ (_00516_, _00397_, _00358_);
  and _22348_ (_00517_, _00516_, _00515_);
  or _22349_ (_00518_, _00517_, _00514_);
  or _22350_ (_00519_, _00518_, _00509_);
  or _22351_ (_00520_, _00519_, _00199_);
  and _22352_ (_00521_, _00520_, _00204_);
  and _22353_ (_00522_, _00521_, _00504_);
  and _22354_ (_00523_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _22355_ (_00524_, _00523_, _00522_);
  and _22356_ (_12311_, _00524_, _05141_);
  nand _22357_ (_00525_, _00199_, _06178_);
  and _22358_ (_00526_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _22359_ (_00527_, _00526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _22360_ (_00528_, _00432_);
  and _22361_ (_00529_, _00528_, _00409_);
  or _22362_ (_00530_, _00529_, _00187_);
  and _22363_ (_00531_, _00530_, _00527_);
  and _22364_ (_00532_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _22365_ (_00533_, _00532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _22366_ (_00534_, _00533_, _00464_);
  nor _22367_ (_00535_, _00534_, _00439_);
  and _22368_ (_00536_, _00193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _22369_ (_00537_, _00536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _22370_ (_00538_, _00394_, _00358_);
  and _22371_ (_00539_, _00538_, _00537_);
  or _22372_ (_00540_, _00539_, _00535_);
  or _22373_ (_00541_, _00540_, _00531_);
  or _22374_ (_00542_, _00541_, _00199_);
  and _22375_ (_00543_, _00542_, _00525_);
  or _22376_ (_00544_, _00543_, _00203_);
  or _22377_ (_00545_, _00204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22378_ (_00546_, _00545_, _05141_);
  and _22379_ (_12324_, _00546_, _00544_);
  or _22380_ (_00547_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not _22381_ (_00548_, _00526_);
  and _22382_ (_00549_, _00548_, _00455_);
  and _22383_ (_00550_, _00549_, _00547_);
  nor _22384_ (_00551_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _22385_ (_00552_, _00551_, _00532_);
  and _22386_ (_00553_, _00552_, _00464_);
  or _22387_ (_00554_, _00193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _22388_ (_00555_, _00536_, _00358_);
  and _22389_ (_00556_, _00555_, _00554_);
  or _22390_ (_00557_, _00556_, _00553_);
  or _22391_ (_00558_, _00557_, _00550_);
  or _22392_ (_00559_, _00558_, _00199_);
  nand _22393_ (_00560_, _00199_, _05604_);
  and _22394_ (_00561_, _00560_, _00559_);
  or _22395_ (_00562_, _00561_, _00203_);
  not _22396_ (_00563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _22397_ (_00564_, _00203_, _00563_);
  and _22398_ (_00565_, _00564_, _05141_);
  and _22399_ (_12328_, _00565_, _00562_);
  and _22400_ (_00566_, _08242_, _05649_);
  nand _22401_ (_00567_, _00566_, _05604_);
  or _22402_ (_00568_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22403_ (_00569_, _00568_, _05141_);
  and _22404_ (_12334_, _00569_, _00567_);
  nand _22405_ (_00570_, _00566_, _06178_);
  or _22406_ (_00571_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22407_ (_00572_, _00571_, _05141_);
  and _22408_ (_12337_, _00572_, _00570_);
  or _22409_ (_00573_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _22410_ (_00574_, _00573_, _05141_);
  and _22411_ (_00575_, _06184_, _05925_);
  nand _22412_ (_00576_, _00575_, _06062_);
  and _22413_ (_12342_, _00576_, _00574_);
  or _22414_ (_00577_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _22415_ (_00578_, _00577_, _05141_);
  not _22416_ (_00579_, _00575_);
  or _22417_ (_00580_, _00579_, _05522_);
  and _22418_ (_12345_, _00580_, _00578_);
  nand _22419_ (_00581_, _00566_, _05560_);
  or _22420_ (_00582_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _22421_ (_00583_, _00582_, _05141_);
  and _22422_ (_12348_, _00583_, _00581_);
  or _22423_ (_00584_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _22424_ (_00585_, _00584_, _05141_);
  nand _22425_ (_00586_, _00575_, _06244_);
  and _22426_ (_12353_, _00586_, _00585_);
  or _22427_ (_00587_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _22428_ (_00588_, _00587_, _05141_);
  or _22429_ (_00589_, _00579_, _06004_);
  and _22430_ (_12360_, _00589_, _00588_);
  nand _22431_ (_00590_, _08305_, _06244_);
  or _22432_ (_00591_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _22433_ (_00592_, _00591_, _05141_);
  and _22434_ (_12406_, _00592_, _00590_);
  and _22435_ (_00593_, _05614_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _22436_ (_00594_, _06179_, _05617_);
  nand _22437_ (_00595_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _22438_ (_00596_, _00595_, _05609_);
  or _22439_ (_00597_, _00596_, _00594_);
  or _22440_ (_00598_, _00597_, _00593_);
  and _22441_ (_12536_, _00598_, _05141_);
  not _22442_ (_00599_, _05576_);
  nor _22443_ (_00600_, _05960_, _00599_);
  and _22444_ (_00601_, _00599_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or _22445_ (_00602_, _00601_, _05572_);
  or _22446_ (_00603_, _00602_, _00600_);
  or _22447_ (_00604_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _22448_ (_00605_, _00604_, _05141_);
  and _22449_ (_12620_, _00605_, _00603_);
  or _22450_ (_00606_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand _22451_ (_00607_, _07619_, _06427_);
  and _22452_ (_00608_, _00607_, _05141_);
  and _22453_ (_12623_, _00608_, _00606_);
  nor _22454_ (_00609_, _12628_, _06791_);
  not _22455_ (_00610_, _12115_);
  or _22456_ (_00611_, _12118_, _12130_);
  or _22457_ (_00612_, _00611_, _00610_);
  and _22458_ (_00613_, _07051_, _12627_);
  nand _22459_ (_00614_, _00613_, _07034_);
  or _22460_ (_00615_, _00614_, _12129_);
  or _22461_ (_00616_, _00615_, _00612_);
  and _22462_ (_00617_, _00616_, _06821_);
  or _22463_ (_00618_, _00617_, _00609_);
  and _22464_ (_12630_, _00618_, _05141_);
  and _22465_ (_00619_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _07611_);
  and _22466_ (_00620_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22467_ (_00621_, _00620_, _00619_);
  and _22468_ (_12648_, _00621_, _05141_);
  nor _22469_ (_12656_, _12827_, rst);
  and _22470_ (_00622_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07611_);
  and _22471_ (_00623_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22472_ (_00624_, _00623_, _00622_);
  and _22473_ (_12661_, _00624_, _05141_);
  not _22474_ (_00625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _22475_ (_00626_, _06683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _22476_ (_00627_, _00626_, _00625_);
  and _22477_ (_00628_, _00627_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _22478_ (_00629_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _22479_ (_00630_, _00627_, _00629_);
  or _22480_ (_00631_, _00630_, _00628_);
  or _22481_ (_00632_, _00631_, _08280_);
  or _22482_ (_00633_, _06620_, _00629_);
  nand _22483_ (_00634_, _00633_, _08280_);
  or _22484_ (_00635_, _00634_, _10356_);
  and _22485_ (_00636_, _00635_, _00632_);
  or _22486_ (_00637_, _00636_, _08289_);
  nand _22487_ (_00638_, _08289_, _05560_);
  and _22488_ (_00639_, _00638_, _05141_);
  and _22489_ (_12722_, _00639_, _00637_);
  and _22490_ (_00640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _05141_);
  and _22491_ (_00641_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05141_);
  and _22492_ (_00642_, _00641_, _11644_);
  or _22493_ (_12734_, _00642_, _00640_);
  and _22494_ (_00643_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _22495_ (_00644_, _00643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _22496_ (_12738_, _00644_, _05141_);
  and _22497_ (_00645_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _07611_);
  and _22498_ (_00646_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22499_ (_00647_, _00646_, _00645_);
  and _22500_ (_12767_, _00647_, _05141_);
  and _22501_ (_12788_, _12409_, _05141_);
  nor _22502_ (_12791_, _12876_, rst);
  or _22503_ (_00648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _22504_ (_00649_, _00648_, _08280_);
  not _22505_ (_00650_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _22506_ (_00651_, _05288_, _00650_);
  nand _22507_ (_00652_, _00651_, _08280_);
  or _22508_ (_00653_, _00652_, _08178_);
  and _22509_ (_00654_, _00653_, _00649_);
  or _22510_ (_00655_, _00654_, _08289_);
  nand _22511_ (_00656_, _08289_, _06178_);
  and _22512_ (_00658_, _00656_, _05141_);
  and _22513_ (_12815_, _00658_, _00655_);
  and _22514_ (_12854_, _12257_, _05141_);
  and _22515_ (_12856_, _12325_, _05141_);
  nand _22516_ (_12858_, _12569_, _05141_);
  nand _22517_ (_12861_, _12515_, _05141_);
  and _22518_ (_00659_, _08280_, _10407_);
  and _22519_ (_00661_, _00659_, _05963_);
  nor _22520_ (_00662_, _00659_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _22521_ (_00663_, _00662_, _00661_);
  nand _22522_ (_00664_, _00663_, _08360_);
  or _22523_ (_00665_, _08360_, _06004_);
  and _22524_ (_00667_, _00665_, _05141_);
  and _22525_ (_12925_, _00667_, _00664_);
  or _22526_ (_00668_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  not _22527_ (_00669_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _22528_ (_00671_, pc_log_change, _00669_);
  and _22529_ (_00672_, _00671_, _05141_);
  and _22530_ (_13021_, _00672_, _00668_);
  and _22531_ (_00673_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _22532_ (_00674_, pc_log_change, _00669_);
  or _22533_ (_00675_, _00674_, _00673_);
  and _22534_ (_13030_, _00675_, _05141_);
  and _22535_ (_00676_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _22536_ (_00677_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _22537_ (_00678_, pc_log_change, _00677_);
  or _22538_ (_00679_, _00678_, _00676_);
  and _22539_ (_13067_, _00679_, _05141_);
  nand _22540_ (_00680_, _06707_, _05560_);
  or _22541_ (_00681_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _22542_ (_00682_, _00681_, _05141_);
  and _22543_ (_13174_, _00682_, _00680_);
  and _22544_ (_13205_, _12390_, _05141_);
  and _22545_ (_13207_, _10319_, _12164_);
  and _22546_ (_00683_, _05299_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _22547_ (_00685_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _22548_ (_00686_, _00685_, _05303_);
  and _22549_ (_00687_, _05605_, _05284_);
  or _22550_ (_00688_, _00687_, _00686_);
  or _22551_ (_00689_, _00688_, _00683_);
  and _22552_ (_13260_, _00689_, _05141_);
  and _22553_ (_00690_, _10342_, _06879_);
  and _22554_ (_00691_, _00690_, _06207_);
  nand _22555_ (_00692_, _00691_, _05963_);
  or _22556_ (_00693_, _00691_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _22557_ (_00694_, _00693_, _05647_);
  and _22558_ (_00695_, _00694_, _00692_);
  not _22559_ (_00696_, _05646_);
  and _22560_ (_00697_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _22561_ (_00698_, _00690_, _05210_);
  not _22562_ (_00699_, _00698_);
  or _22563_ (_00700_, _00699_, _06669_);
  or _22564_ (_00701_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _22565_ (_00702_, _00701_, _05925_);
  and _22566_ (_00703_, _00702_, _00700_);
  or _22567_ (_00704_, _00703_, _00697_);
  or _22568_ (_00705_, _00704_, _00695_);
  and _22569_ (_13332_, _00705_, _05141_);
  and _22570_ (_00707_, _00690_, _05288_);
  nand _22571_ (_00708_, _00707_, _05963_);
  or _22572_ (_00709_, _00707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _22573_ (_00710_, _00709_, _05647_);
  and _22574_ (_00711_, _00710_, _00708_);
  and _22575_ (_00712_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _22576_ (_00713_, _00699_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor _22577_ (_00714_, _00699_, _07434_);
  or _22578_ (_00715_, _00714_, _00713_);
  and _22579_ (_00716_, _00715_, _05925_);
  or _22580_ (_00717_, _00716_, _00712_);
  or _22581_ (_00718_, _00717_, _00711_);
  and _22582_ (_13352_, _00718_, _05141_);
  or _22583_ (_00719_, _00699_, _05922_);
  or _22584_ (_00720_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _22585_ (_00721_, _00720_, _05647_);
  and _22586_ (_00722_, _00721_, _00719_);
  and _22587_ (_00723_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _22588_ (_00724_, _00698_, _07496_);
  and _22589_ (_00725_, _00720_, _05925_);
  and _22590_ (_00726_, _00725_, _00724_);
  or _22591_ (_00727_, _00726_, _00723_);
  or _22592_ (_00728_, _00727_, _00722_);
  and _22593_ (_13367_, _00728_, _05141_);
  not _22594_ (_00729_, _00690_);
  or _22595_ (_00730_, _00729_, _10375_);
  and _22596_ (_00731_, _00730_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _22597_ (_00732_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _22598_ (_00733_, _00732_, _10380_);
  and _22599_ (_00734_, _00733_, _00690_);
  or _22600_ (_00735_, _00734_, _00731_);
  and _22601_ (_00736_, _00735_, _05647_);
  not _22602_ (_00737_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor _22603_ (_00738_, _05646_, _00737_);
  nand _22604_ (_00739_, _00698_, _07259_);
  or _22605_ (_00740_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _22606_ (_00741_, _00740_, _05925_);
  and _22607_ (_00742_, _00741_, _00739_);
  or _22608_ (_00743_, _00742_, _00738_);
  or _22609_ (_00744_, _00743_, _00736_);
  and _22610_ (_13380_, _00744_, _05141_);
  nand _22611_ (_00745_, _00690_, _05186_);
  and _22612_ (_00746_, _00745_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not _22613_ (_00747_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor _22614_ (_00748_, _08282_, _00747_);
  or _22615_ (_00749_, _00748_, _08281_);
  and _22616_ (_00750_, _00749_, _00690_);
  or _22617_ (_00751_, _00750_, _00746_);
  and _22618_ (_00752_, _00751_, _05647_);
  nor _22619_ (_00753_, _05646_, _00747_);
  nand _22620_ (_00754_, _00698_, _07350_);
  or _22621_ (_00755_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _22622_ (_00756_, _00755_, _05925_);
  and _22623_ (_00757_, _00756_, _00754_);
  or _22624_ (_00758_, _00757_, _00753_);
  or _22625_ (_00759_, _00758_, _00752_);
  and _22626_ (_13387_, _00759_, _05141_);
  and _22627_ (_00760_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _22628_ (_00761_, _00760_, _10380_);
  and _22629_ (_00762_, _00761_, _08280_);
  not _22630_ (_00763_, _08280_);
  or _22631_ (_00764_, _00763_, _10375_);
  and _22632_ (_00765_, _00764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _22633_ (_00766_, _00765_, _08289_);
  or _22634_ (_00767_, _00766_, _00762_);
  or _22635_ (_00768_, _08360_, _05522_);
  and _22636_ (_00769_, _00768_, _05141_);
  and _22637_ (_13390_, _00769_, _00767_);
  or _22638_ (_00770_, _12096_, _12030_);
  and _22639_ (_00771_, _00770_, _12097_);
  or _22640_ (_00772_, _00771_, _07135_);
  or _22641_ (_00773_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _22642_ (_00774_, _00773_, _12108_);
  and _22643_ (_00775_, _00774_, _00772_);
  and _22644_ (_00776_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _22645_ (_13411_, _00776_, _00775_);
  nand _22646_ (_00777_, _12099_, _12025_);
  and _22647_ (_00779_, _00777_, _12100_);
  or _22648_ (_00780_, _00779_, _07135_);
  or _22649_ (_00781_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _22650_ (_00782_, _00781_, _12108_);
  and _22651_ (_00783_, _00782_, _00780_);
  and _22652_ (_00784_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _22653_ (_13431_, _00784_, _00783_);
  nand _22654_ (_00785_, _12097_, _12027_);
  and _22655_ (_00786_, _00785_, _12099_);
  or _22656_ (_00787_, _00786_, _07135_);
  or _22657_ (_00789_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _22658_ (_00790_, _00789_, _12108_);
  and _22659_ (_00791_, _00790_, _00787_);
  and _22660_ (_00792_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _22661_ (_13436_, _00792_, _00791_);
  nor _22662_ (_00793_, _12075_, _12072_);
  nor _22663_ (_00794_, _00793_, _12077_);
  or _22664_ (_00795_, _00794_, _07135_);
  or _22665_ (_00796_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _22666_ (_00797_, _00796_, _12108_);
  and _22667_ (_00798_, _00797_, _00795_);
  and _22668_ (_00799_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _22669_ (_00147_, _00799_, _00798_);
  nor _22670_ (_00800_, _12087_, _12084_);
  nor _22671_ (_00801_, _00800_, _12088_);
  or _22672_ (_00802_, _00801_, _07135_);
  or _22673_ (_00803_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _22674_ (_00804_, _00803_, _12108_);
  and _22675_ (_00805_, _00804_, _00802_);
  and _22676_ (_00806_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _22677_ (_00158_, _00806_, _00805_);
  nor _22678_ (_00808_, _12083_, _12063_);
  nor _22679_ (_00809_, _00808_, _12084_);
  or _22680_ (_00810_, _00809_, _07135_);
  or _22681_ (_00811_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _22682_ (_00812_, _00811_, _12108_);
  and _22683_ (_00813_, _00812_, _00810_);
  and _22684_ (_00814_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _22685_ (_00172_, _00814_, _00813_);
  and _22686_ (_00815_, _11976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _22687_ (_00816_, _12081_, _12078_);
  nor _22688_ (_00817_, _00816_, _12083_);
  or _22689_ (_00818_, _00817_, _07135_);
  or _22690_ (_00819_, _07134_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _22691_ (_00820_, _00819_, _12108_);
  and _22692_ (_00821_, _00820_, _00818_);
  or _22693_ (_00209_, _00821_, _00815_);
  nand _22694_ (_00822_, _00203_, _05960_);
  and _22695_ (_00823_, _00358_, _00194_);
  nand _22696_ (_00824_, _00823_, _00193_);
  nor _22697_ (_00825_, _00824_, _00199_);
  or _22698_ (_00827_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _22699_ (_00828_, _00408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _22700_ (_00829_, _00828_, _00186_);
  nand _22701_ (_00830_, _00829_, _00196_);
  or _22702_ (_00831_, _00830_, _00199_);
  and _22703_ (_00832_, _00831_, _00827_);
  or _22704_ (_00833_, _00832_, _00203_);
  and _22705_ (_00834_, _00833_, _05141_);
  and _22706_ (_00341_, _00834_, _00822_);
  or _22707_ (_00835_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _22708_ (_00836_, _00464_, _05141_);
  and _22709_ (_00837_, _00836_, _00835_);
  not _22710_ (_00838_, _00414_);
  and _22711_ (_00839_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22712_ (_00840_, _00839_, _00838_);
  nand _22713_ (_00841_, _00840_, _00837_);
  nor _22714_ (_00842_, _00841_, _00203_);
  and _22715_ (_00343_, _00842_, _00378_);
  nand _22716_ (_00843_, _00199_, _05960_);
  and _22717_ (_00844_, _00507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _22718_ (_00845_, _00844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22719_ (_00846_, _00844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _22720_ (_00847_, _00846_, _00845_);
  and _22721_ (_00848_, _00847_, _00455_);
  not _22722_ (_00849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _22723_ (_00850_, _00414_, _00410_);
  and _22724_ (_00851_, _00850_, _00849_);
  nor _22725_ (_00852_, _00850_, _00849_);
  or _22726_ (_00854_, _00852_, _00851_);
  and _22727_ (_00856_, _00854_, _00464_);
  and _22728_ (_00857_, _00410_, _00193_);
  or _22729_ (_00858_, _00857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _22730_ (_00859_, _00858_, _00356_);
  and _22731_ (_00860_, _00839_, _00193_);
  nor _22732_ (_00861_, _00860_, _00859_);
  or _22733_ (_00862_, _00861_, _00856_);
  or _22734_ (_00864_, _00862_, _00199_);
  or _22735_ (_00865_, _00864_, _00848_);
  and _22736_ (_00866_, _00865_, _00204_);
  and _22737_ (_00867_, _00866_, _00843_);
  and _22738_ (_00868_, _00203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22739_ (_00869_, _00868_, _00867_);
  and _22740_ (_00345_, _00869_, _05141_);
  nand _22741_ (_00870_, _06707_, _06244_);
  or _22742_ (_00871_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _22743_ (_00872_, _00871_, _05141_);
  and _22744_ (_00349_, _00872_, _00870_);
  or _22745_ (_00873_, _00566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _22746_ (_00874_, _00873_, _05141_);
  nand _22747_ (_00875_, _00575_, _05960_);
  and _22748_ (_00355_, _00875_, _00874_);
  or _22749_ (_00876_, _12914_, _12773_);
  or _22750_ (_00877_, _00876_, _05739_);
  nor _22751_ (_00878_, _12772_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _22752_ (_00879_, _00878_, _12906_);
  and _22753_ (_00880_, _00879_, _00877_);
  nor _22754_ (_00881_, _00880_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _22755_ (_00882_, _00880_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _22756_ (_00883_, _00882_, _00881_);
  and _22757_ (_00884_, _00883_, _12973_);
  and _22758_ (_00885_, _12701_, _07288_);
  and _22759_ (_00886_, _11451_, _06669_);
  and _22760_ (_00887_, _12707_, _12776_);
  nand _22761_ (_00888_, _12726_, _05699_);
  and _22762_ (_00889_, _00888_, _12727_);
  and _22763_ (_00891_, _00889_, _12713_);
  or _22764_ (_00892_, _00891_, _00887_);
  and _22765_ (_00893_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _22766_ (_00894_, _00893_, _00892_);
  or _22767_ (_00895_, _00894_, _00886_);
  or _22768_ (_00896_, _00895_, _00885_);
  or _22769_ (_00897_, _00896_, _00884_);
  or _22770_ (_00898_, _00897_, _13052_);
  nor _22771_ (_00900_, _12955_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _22772_ (_00901_, _00900_, _12956_);
  or _22773_ (_00902_, _00901_, _12700_);
  and _22774_ (_00903_, _00902_, _05141_);
  and _22775_ (_00357_, _00903_, _00898_);
  and _22776_ (_00366_, t0_i, _05141_);
  and _22777_ (_00370_, t1_i, _05141_);
  and _22778_ (_00904_, _13439_, _05960_);
  and _22779_ (_00905_, _00102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _22780_ (_00906_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _22781_ (_00907_, _00906_, _00905_);
  and _22782_ (_00908_, _00907_, _00038_);
  or _22783_ (_00909_, _00908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _22784_ (_00910_, _00908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _22785_ (_00912_, _00910_, _00033_);
  and _22786_ (_00913_, _00912_, _00909_);
  and _22787_ (_00914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _22788_ (_00915_, _00907_, _00069_);
  or _22789_ (_00916_, _00915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not _22790_ (_00917_, _00048_);
  and _22791_ (_00918_, _00915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _22792_ (_00919_, _00918_, _00917_);
  and _22793_ (_00920_, _00919_, _00916_);
  or _22794_ (_00921_, _00920_, _00914_);
  nor _22795_ (_00922_, _00921_, _00913_);
  and _22796_ (_00923_, _00922_, _13375_);
  or _22797_ (_00924_, _00923_, _00904_);
  nand _22798_ (_00925_, _00924_, _00060_);
  or _22799_ (_00926_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _22800_ (_00927_, _00926_, _05141_);
  and _22801_ (_00374_, _00927_, _00925_);
  and _22802_ (_00928_, _00233_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  or _22803_ (_00929_, _00928_, _00860_);
  and _22804_ (_00930_, _00929_, _00356_);
  or _22805_ (_00931_, _00928_, _00196_);
  or _22806_ (_00932_, _00928_, _00839_);
  and _22807_ (_00933_, _00932_, _00409_);
  and _22808_ (_00934_, _00933_, _00931_);
  and _22809_ (_00935_, _00931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _22810_ (_00936_, _00935_, _00934_);
  or _22811_ (_00937_, _00936_, _00930_);
  nand _22812_ (_00938_, _00937_, _05141_);
  nor _22813_ (_00939_, _00938_, _00203_);
  and _22814_ (_00376_, _00939_, _00378_);
  not _22815_ (_00940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _22816_ (_00941_, _13389_, _00940_);
  or _22817_ (_00942_, _00941_, _00918_);
  and _22818_ (_00943_, _00942_, _00048_);
  or _22819_ (_00944_, _00941_, _00910_);
  and _22820_ (_00945_, _00944_, _13372_);
  nand _22821_ (_00946_, _13389_, _13369_);
  and _22822_ (_00947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _22823_ (_00948_, _00947_, _00946_);
  or _22824_ (_00949_, _00948_, _13443_);
  or _22825_ (_00950_, _00949_, _00945_);
  or _22826_ (_00951_, _00950_, _00943_);
  and _22827_ (_00952_, _13366_, _13375_);
  and _22828_ (_00953_, _00952_, _05141_);
  and _22829_ (_00377_, _00953_, _00951_);
  nor _22830_ (_00954_, _13400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _22831_ (_00955_, _00954_, _13401_);
  and _22832_ (_00956_, _00955_, _13374_);
  and _22833_ (_00957_, _13402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _22834_ (_00958_, _00957_, _00956_);
  and _22835_ (_00959_, _00958_, _00953_);
  and _22836_ (_00960_, _13377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _22837_ (_00961_, _00960_, _13366_);
  nor _22838_ (_00962_, _00060_, _05960_);
  or _22839_ (_00963_, _00962_, _00961_);
  and _22840_ (_00964_, _00963_, _05141_);
  or _22841_ (_00379_, _00964_, _00959_);
  nand _22842_ (_00965_, _12906_, _12773_);
  and _22843_ (_00966_, _00965_, _00876_);
  nand _22844_ (_00967_, _00966_, _05739_);
  or _22845_ (_00968_, _00966_, _05739_);
  and _22846_ (_00969_, _00968_, _12973_);
  and _22847_ (_00970_, _00969_, _00967_);
  and _22848_ (_00971_, _12701_, _07166_);
  nand _22849_ (_00972_, _12725_, _05739_);
  and _22850_ (_00973_, _00972_, _12726_);
  and _22851_ (_00974_, _00973_, _12713_);
  nor _22852_ (_00975_, _12703_, _07200_);
  or _22853_ (_00976_, _00975_, _00974_);
  and _22854_ (_00977_, _12707_, _12808_);
  and _22855_ (_00979_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _22856_ (_00981_, _00979_, _00977_);
  or _22857_ (_00982_, _00981_, _00976_);
  nor _22858_ (_00983_, _00982_, _00971_);
  nand _22859_ (_00984_, _00983_, _12700_);
  or _22860_ (_00985_, _00984_, _00970_);
  nor _22861_ (_00986_, _12954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _22862_ (_00988_, _00986_, _12955_);
  or _22863_ (_00989_, _00988_, _12700_);
  and _22864_ (_00990_, _00989_, _05141_);
  and _22865_ (_00387_, _00990_, _00985_);
  and _22866_ (_00991_, _05568_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _22867_ (_00992_, _05522_, _05291_);
  or _22868_ (_00993_, _00992_, _05572_);
  or _22869_ (_00994_, _00993_, _00991_);
  or _22870_ (_00995_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _22871_ (_00996_, _00995_, _05141_);
  and _22872_ (_00457_, _00996_, _00994_);
  and _22873_ (_00997_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _22874_ (_00998_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _22875_ (_00999_, _00998_, _06156_);
  and _22876_ (_01000_, _06180_, _05561_);
  or _22877_ (_01001_, _01000_, _00999_);
  or _22878_ (_01002_, _01001_, _00997_);
  and _22879_ (_00486_, _01002_, _05141_);
  not _22880_ (_01003_, _12827_);
  and _22881_ (_01004_, _01003_, _12707_);
  not _22882_ (_01006_, _07200_);
  and _22883_ (_01007_, _13058_, _01006_);
  and _22884_ (_01008_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _22885_ (_01009_, _12713_, _12808_);
  or _22886_ (_01010_, _01009_, _01008_);
  or _22887_ (_01011_, _01010_, _01007_);
  nand _22888_ (_01012_, _12898_, _12896_);
  nand _22889_ (_01013_, _01012_, _12835_);
  nand _22890_ (_01014_, _12837_, _01013_);
  or _22891_ (_01015_, _12837_, _01013_);
  and _22892_ (_01016_, _01015_, _12940_);
  and _22893_ (_01017_, _01016_, _01014_);
  or _22894_ (_01018_, _01017_, _01011_);
  or _22895_ (_01019_, _01018_, _01004_);
  and _22896_ (_01020_, _01019_, _12700_);
  nor _22897_ (_01021_, _00226_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _22898_ (_01022_, _01021_, _00228_);
  nor _22899_ (_01023_, _01022_, _12700_);
  or _22900_ (_01024_, _01023_, _01020_);
  and _22901_ (_00657_, _01024_, _05141_);
  not _22902_ (_01026_, _07593_);
  and _22903_ (_01028_, _12707_, _01026_);
  not _22904_ (_01029_, _07259_);
  and _22905_ (_01031_, _13058_, _01029_);
  and _22906_ (_01033_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _22907_ (_01034_, _12713_, _12831_);
  or _22908_ (_01035_, _01034_, _01033_);
  or _22909_ (_01036_, _01035_, _01031_);
  or _22910_ (_01037_, _01036_, _01028_);
  or _22911_ (_01038_, _12898_, _12896_);
  and _22912_ (_01039_, _01038_, _01012_);
  and _22913_ (_01040_, _01039_, _12940_);
  or _22914_ (_01041_, _01040_, _01037_);
  and _22915_ (_01042_, _01041_, _12700_);
  nor _22916_ (_01043_, _07622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _22917_ (_01044_, _01043_, _00226_);
  nor _22918_ (_01045_, _01044_, _12700_);
  or _22919_ (_01046_, _01045_, _01042_);
  and _22920_ (_00660_, _01046_, _05141_);
  not _22921_ (_01047_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _22922_ (_01048_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _22923_ (_01049_, _01048_, _01047_);
  nor _22924_ (_01050_, _01049_, rst);
  nand _22925_ (_01051_, _01048_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _22926_ (_01052_, _01048_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _22927_ (_01053_, _01052_, _01051_);
  and _22928_ (_00666_, _01053_, _01050_);
  or _22929_ (_01054_, _12847_, _12848_);
  not _22930_ (_01055_, _01054_);
  nand _22931_ (_01056_, _01055_, _12894_);
  or _22932_ (_01057_, _01055_, _12894_);
  and _22933_ (_01058_, _01057_, _12973_);
  and _22934_ (_01059_, _01058_, _01056_);
  not _22935_ (_01060_, _07350_);
  and _22936_ (_01061_, _13058_, _01060_);
  not _22937_ (_01062_, _07572_);
  and _22938_ (_01063_, _12707_, _01062_);
  and _22939_ (_01064_, _12713_, _12843_);
  and _22940_ (_01065_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _22941_ (_01066_, _01065_, _01064_);
  or _22942_ (_01067_, _01066_, _01063_);
  or _22943_ (_01068_, _01067_, _01061_);
  or _22944_ (_01069_, _01068_, _01059_);
  and _22945_ (_01070_, _01069_, _12700_);
  and _22946_ (_01071_, _13052_, _07623_);
  or _22947_ (_01072_, _01071_, _01070_);
  and _22948_ (_00670_, _01072_, _05141_);
  not _22949_ (_01073_, _07550_);
  and _22950_ (_01074_, _12707_, _01073_);
  not _22951_ (_01075_, _06617_);
  and _22952_ (_01076_, _13058_, _01075_);
  and _22953_ (_01077_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _22954_ (_01078_, _12713_, _12849_);
  or _22955_ (_01079_, _01078_, _01077_);
  or _22956_ (_01080_, _01079_, _01076_);
  or _22957_ (_01081_, _12892_, _12889_);
  not _22958_ (_01082_, _12893_);
  and _22959_ (_01083_, _12940_, _01082_);
  and _22960_ (_01084_, _01083_, _01081_);
  or _22961_ (_01085_, _01084_, _01080_);
  or _22962_ (_01086_, _01085_, _01074_);
  and _22963_ (_01087_, _01086_, _12700_);
  and _22964_ (_01088_, _13052_, _07636_);
  or _22965_ (_01089_, _01088_, _01087_);
  and _22966_ (_00684_, _01089_, _05141_);
  not _22967_ (_01090_, _07434_);
  and _22968_ (_01091_, _13058_, _01090_);
  not _22969_ (_01092_, _12876_);
  and _22970_ (_01093_, _01092_, _12707_);
  and _22971_ (_01094_, _12713_, _12855_);
  and _22972_ (_01095_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _22973_ (_01096_, _01095_, _01094_);
  or _22974_ (_01097_, _01096_, _01093_);
  or _22975_ (_01098_, _01097_, _01091_);
  nor _22976_ (_01099_, _12887_, _12884_);
  nor _22977_ (_01100_, _01099_, _12888_);
  and _22978_ (_01101_, _01100_, _12940_);
  or _22979_ (_01102_, _01101_, _01098_);
  or _22980_ (_01103_, _01102_, _13052_);
  or _22981_ (_01104_, _12700_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _22982_ (_01105_, _01104_, _05141_);
  and _22983_ (_00706_, _01105_, _01103_);
  and _22984_ (_01106_, _12701_, _07378_);
  and _22985_ (_01107_, _12707_, _12849_);
  nor _22986_ (_01108_, _12703_, _06617_);
  or _22987_ (_01109_, _01108_, _01107_);
  and _22988_ (_01110_, _12713_, _07014_);
  and _22989_ (_01111_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _22990_ (_01112_, _01111_, _01110_);
  or _22991_ (_01113_, _01112_, _01109_);
  or _22992_ (_01114_, _01113_, _01106_);
  nor _22993_ (_01115_, _12904_, _12772_);
  and _22994_ (_01116_, _12902_, _12910_);
  nor _22995_ (_01117_, _01116_, _12773_);
  or _22996_ (_01118_, _01117_, _01115_);
  nand _22997_ (_01119_, _01118_, _05455_);
  or _22998_ (_01120_, _01118_, _05455_);
  and _22999_ (_01121_, _01120_, _01119_);
  and _23000_ (_01122_, _01121_, _12940_);
  or _23001_ (_01123_, _01122_, _01114_);
  or _23002_ (_01124_, _01123_, _13052_);
  nor _23003_ (_01125_, _13001_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _23004_ (_01126_, _01125_, _13002_);
  or _23005_ (_01127_, _01126_, _12700_);
  and _23006_ (_01128_, _01127_, _05141_);
  and _23007_ (_00778_, _01128_, _01124_);
  and _23008_ (_01129_, _12701_, _07406_);
  and _23009_ (_01130_, _12707_, _12855_);
  and _23010_ (_01131_, _12713_, _06524_);
  or _23011_ (_01132_, _01131_, _01130_);
  and _23012_ (_01133_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _23013_ (_01134_, _11451_, _01090_);
  or _23014_ (_01135_, _01134_, _01133_);
  or _23015_ (_01136_, _01135_, _01132_);
  or _23016_ (_01137_, _01136_, _01129_);
  and _23017_ (_01138_, _12902_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _23018_ (_01139_, _01138_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _23019_ (_01140_, _01139_, _01117_);
  and _23020_ (_01141_, _12903_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _23021_ (_01142_, _01141_, _12904_);
  and _23022_ (_01143_, _01142_, _12773_);
  or _23023_ (_01144_, _01143_, _01140_);
  and _23024_ (_01145_, _01144_, _12940_);
  or _23025_ (_01146_, _01145_, _01137_);
  or _23026_ (_01147_, _01146_, _13052_);
  nor _23027_ (_01148_, _13000_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _23028_ (_01150_, _01148_, _13001_);
  or _23029_ (_01151_, _01150_, _12700_);
  and _23030_ (_01152_, _01151_, _05141_);
  and _23031_ (_00788_, _01152_, _01147_);
  and _23032_ (_01153_, _12701_, _07466_);
  and _23033_ (_01154_, _12707_, _12880_);
  and _23034_ (_01155_, _11451_, _13057_);
  or _23035_ (_01156_, _01155_, _01154_);
  and _23036_ (_01157_, _12713_, _06497_);
  and _23037_ (_01158_, _12745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _23038_ (_01159_, _01158_, _01157_);
  or _23039_ (_01160_, _01159_, _01156_);
  or _23040_ (_01161_, _01160_, _01153_);
  and _23041_ (_01162_, _12902_, _05411_);
  nor _23042_ (_01163_, _12902_, _05411_);
  nor _23043_ (_01164_, _01163_, _01162_);
  nand _23044_ (_01165_, _01164_, _12772_);
  or _23045_ (_01166_, _01164_, _12772_);
  and _23046_ (_01167_, _01166_, _01165_);
  and _23047_ (_01168_, _01167_, _12940_);
  nor _23048_ (_01169_, _01168_, _01161_);
  nand _23049_ (_01170_, _01169_, _12700_);
  nor _23050_ (_01171_, _12999_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _23051_ (_01172_, _01171_, _13000_);
  or _23052_ (_01173_, _01172_, _12700_);
  and _23053_ (_01174_, _01173_, _05141_);
  and _23054_ (_00807_, _01174_, _01170_);
  not _23055_ (_01175_, _06875_);
  and _23056_ (_01176_, _13058_, _01175_);
  not _23057_ (_01177_, _12770_);
  and _23058_ (_01178_, _01177_, _12707_);
  and _23059_ (_01179_, _12713_, _12732_);
  and _23060_ (_01180_, _11451_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _23061_ (_01181_, _01180_, _01179_);
  or _23062_ (_01182_, _01181_, _01178_);
  or _23063_ (_01184_, _01182_, _01176_);
  nor _23064_ (_01185_, _00219_, _12800_);
  nor _23065_ (_01186_, _01185_, _12802_);
  and _23066_ (_01187_, _01185_, _12802_);
  or _23067_ (_01189_, _01187_, _01186_);
  and _23068_ (_01190_, _01189_, _12940_);
  or _23069_ (_01191_, _01190_, _01184_);
  and _23070_ (_01192_, _01191_, _12700_);
  nor _23071_ (_01193_, _00227_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _23072_ (_01194_, _01193_, _12999_);
  nor _23073_ (_01195_, _01194_, _12700_);
  or _23074_ (_01196_, _01195_, _01192_);
  and _23075_ (_00826_, _01196_, _05141_);
  and _23076_ (_01197_, _11667_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _23077_ (_01198_, _01197_, _11665_);
  and _23078_ (_01199_, _01198_, _06013_);
  not _23079_ (_01200_, _06013_);
  or _23080_ (_01201_, _06209_, _01200_);
  and _23081_ (_01202_, _01201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _23082_ (_01203_, _01202_, _06020_);
  or _23083_ (_01204_, _01203_, _01199_);
  or _23084_ (_01205_, _06021_, _06004_);
  and _23085_ (_01206_, _01205_, _05141_);
  and _23086_ (_00853_, _01206_, _01204_);
  and _23087_ (_01208_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23088_ (_01209_, _01208_, _10356_);
  and _23089_ (_01210_, _01209_, _06013_);
  nand _23090_ (_01211_, _06013_, _08283_);
  and _23091_ (_01212_, _01211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23092_ (_01213_, _01212_, _06020_);
  or _23093_ (_01214_, _01213_, _01210_);
  nand _23094_ (_01215_, _06020_, _05560_);
  and _23095_ (_01216_, _01215_, _05141_);
  and _23096_ (_00863_, _01216_, _01214_);
  and _23097_ (_01217_, _11667_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _23098_ (_01218_, _01217_, _11665_);
  and _23099_ (_01219_, _01218_, _06255_);
  not _23100_ (_01220_, _06255_);
  or _23101_ (_01221_, _01220_, _06209_);
  and _23102_ (_01222_, _01221_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _23103_ (_01223_, _01222_, _06262_);
  or _23104_ (_01224_, _01223_, _01219_);
  or _23105_ (_01225_, _06263_, _06004_);
  and _23106_ (_01226_, _01225_, _05141_);
  and _23107_ (_00890_, _01226_, _01224_);
  and _23108_ (_01227_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23109_ (_01228_, _01227_, _10356_);
  and _23110_ (_01229_, _01228_, _06255_);
  nand _23111_ (_01230_, _06255_, _08283_);
  and _23112_ (_01231_, _01230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23113_ (_01232_, _01231_, _06262_);
  or _23114_ (_01233_, _01232_, _01229_);
  nand _23115_ (_01234_, _06262_, _05560_);
  and _23116_ (_01235_, _01234_, _05141_);
  and _23117_ (_00899_, _01235_, _01233_);
  or _23118_ (_01236_, \oc8051_top_1.oc8051_sfr1.prescaler [2], rst);
  nor _23119_ (_00911_, _01236_, _01051_);
  and _23120_ (_00978_, _00640_, _06065_);
  not _23121_ (_01237_, _06114_);
  nor _23122_ (_01238_, _06102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _23123_ (_01239_, _01238_, _06100_);
  or _23124_ (_01240_, _01239_, _06105_);
  and _23125_ (_01241_, _01240_, _01237_);
  or _23126_ (_01242_, _01241_, _06112_);
  and _23127_ (_01243_, _06133_, _06110_);
  and _23128_ (_01244_, _01243_, _01242_);
  not _23129_ (_01245_, _06078_);
  or _23130_ (_01246_, _06089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23131_ (_01247_, _01246_, _06085_);
  or _23132_ (_01248_, _01247_, _06093_);
  and _23133_ (_01249_, _01248_, _01245_);
  or _23134_ (_01250_, _01249_, _06076_);
  and _23135_ (_01251_, _06097_, _06074_);
  and _23136_ (_01252_, _01251_, _01250_);
  or _23137_ (_01253_, _01252_, _06065_);
  or _23138_ (_01254_, _01253_, _01244_);
  or _23139_ (_01255_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23140_ (_01256_, _01255_, _05141_);
  and _23141_ (_00980_, _01256_, _01254_);
  and _23142_ (_01257_, _06878_, _06009_);
  and _23143_ (_01258_, _01257_, _06008_);
  nand _23144_ (_01259_, _01258_, _05963_);
  or _23145_ (_01260_, _01258_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _23146_ (_01261_, _01260_, _05647_);
  and _23147_ (_01262_, _01261_, _01259_);
  and _23148_ (_01263_, _06261_, _05272_);
  not _23149_ (_01264_, _01263_);
  nor _23150_ (_01265_, _01264_, _05960_);
  and _23151_ (_01266_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _23152_ (_01267_, _01266_, _01265_);
  and _23153_ (_01268_, _01267_, _05925_);
  and _23154_ (_01269_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _23155_ (_01270_, _01269_, rst);
  or _23156_ (_01271_, _01270_, _01268_);
  or _23157_ (_00987_, _01271_, _01262_);
  and _23158_ (_01272_, _06205_, _05210_);
  nand _23159_ (_01273_, _01272_, _05963_);
  or _23160_ (_01274_, _01272_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _23161_ (_01275_, _01274_, _05928_);
  and _23162_ (_01276_, _01275_, _01273_);
  and _23163_ (_01277_, _05927_, _06703_);
  or _23164_ (_01278_, _01277_, _01276_);
  and _23165_ (_01005_, _01278_, _05141_);
  and _23166_ (_01279_, _12559_, _12502_);
  nand _23167_ (_01280_, _12397_, _12391_);
  and _23168_ (_01281_, _01280_, _12450_);
  and _23169_ (_01282_, _12261_, _12310_);
  and _23170_ (_01283_, _01282_, _01281_);
  and _23171_ (_01284_, _12608_, _12372_);
  and _23172_ (_01285_, _01284_, _01283_);
  and _23173_ (_01286_, _01285_, _01279_);
  and _23174_ (_01287_, _01286_, _06619_);
  and _23175_ (_01288_, _12557_, _12502_);
  and _23176_ (_01289_, _12610_, _12374_);
  and _23177_ (_01290_, _01289_, _01288_);
  and _23178_ (_01291_, _01280_, _12448_);
  and _23179_ (_01292_, _01291_, _01282_);
  and _23180_ (_01293_, _01292_, _01290_);
  and _23181_ (_01294_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _23182_ (_01295_, _12608_, _12374_);
  and _23183_ (_01296_, _01288_, _01295_);
  and _23184_ (_01297_, _01296_, _01292_);
  and _23185_ (_01298_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _23186_ (_01299_, _01298_, _01294_);
  and _23187_ (_01300_, _01279_, _01295_);
  and _23188_ (_01301_, _01300_, _01292_);
  and _23189_ (_01302_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _23190_ (_01303_, _12557_, _12504_);
  and _23191_ (_01304_, _01303_, _01289_);
  and _23192_ (_01305_, _01304_, _01292_);
  and _23193_ (_01306_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _23194_ (_01307_, _01306_, _01302_);
  or _23195_ (_01308_, _01307_, _01299_);
  and _23196_ (_01309_, _12559_, _12504_);
  and _23197_ (_01310_, _01295_, _01309_);
  and _23198_ (_01311_, _01292_, _01310_);
  and _23199_ (_01312_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _23200_ (_01313_, _01296_, _01283_);
  and _23201_ (_01314_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _23202_ (_01315_, _01314_, _01312_);
  not _23203_ (_01316_, _01296_);
  nand _23204_ (_01317_, _01281_, _12313_);
  or _23205_ (_01318_, _01317_, _12263_);
  nor _23206_ (_01319_, _01318_, _01316_);
  and _23207_ (_01320_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _23208_ (_01321_, _12263_, _12313_);
  and _23209_ (_01322_, _01321_, _01281_);
  and _23210_ (_01323_, _01309_, _12610_);
  and _23211_ (_01324_, _01323_, _12372_);
  and _23212_ (_01325_, _01324_, _01322_);
  and _23213_ (_01326_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _23214_ (_01327_, _01326_, _01320_);
  or _23215_ (_01328_, _01327_, _01315_);
  or _23216_ (_01329_, _01328_, _01308_);
  and _23217_ (_01330_, _01310_, _01283_);
  and _23218_ (_01331_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _23219_ (_01332_, _01303_, _01295_);
  and _23220_ (_01333_, _01332_, _01283_);
  and _23221_ (_01334_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _23222_ (_01335_, _01334_, _01331_);
  and _23223_ (_01336_, _01300_, _01283_);
  and _23224_ (_01337_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _23225_ (_01338_, _01304_, _01283_);
  and _23226_ (_01339_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _23227_ (_01340_, _01339_, _01337_);
  or _23228_ (_01341_, _01340_, _01335_);
  nand _23229_ (_01342_, _01281_, _12310_);
  nor _23230_ (_01343_, _01342_, _12261_);
  and _23231_ (_01344_, _01343_, _01296_);
  and _23232_ (_01345_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _23233_ (_01346_, _01343_, _01332_);
  and _23234_ (_01347_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _23235_ (_01348_, _01347_, _01345_);
  and _23236_ (_01349_, _01290_, _01283_);
  and _23237_ (_01350_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _23238_ (_01351_, _01324_, _01283_);
  and _23239_ (_01352_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _23240_ (_01353_, _01352_, _01350_);
  or _23241_ (_01354_, _01353_, _01348_);
  or _23242_ (_01355_, _01354_, _01341_);
  or _23243_ (_01356_, _01355_, _01329_);
  and _23244_ (_01357_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _23245_ (_01358_, _01284_, _01309_);
  and _23246_ (_01359_, _01358_, _01283_);
  and _23247_ (_01360_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _23248_ (_01361_, _01360_, _01357_);
  and _23249_ (_01362_, _01291_, _12313_);
  and _23250_ (_01363_, _01284_, _01288_);
  and _23251_ (_01364_, _01363_, _12263_);
  and _23252_ (_01365_, _01364_, _01362_);
  and _23253_ (_01366_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _23254_ (_01367_, _01303_, _01284_);
  and _23255_ (_01368_, _01367_, _01283_);
  and _23256_ (_01369_, _01368_, _12390_);
  or _23257_ (_01370_, _01369_, _01366_);
  or _23258_ (_01371_, _01370_, _01361_);
  not _23259_ (_01372_, _01363_);
  nor _23260_ (_01373_, _01318_, _01372_);
  and _23261_ (_01374_, _07053_, _06417_);
  or _23262_ (_01375_, _01374_, _06563_);
  or _23263_ (_01376_, _01375_, _06777_);
  and _23264_ (_01377_, _01376_, _06773_);
  not _23265_ (_01378_, _01377_);
  and _23266_ (_01379_, _06755_, _06564_);
  or _23267_ (_01380_, _01379_, _07073_);
  or _23268_ (_01381_, _01380_, _12130_);
  or _23269_ (_01382_, _06779_, _06772_);
  and _23270_ (_01383_, _07074_, _06574_);
  or _23271_ (_01384_, _12136_, _01383_);
  or _23272_ (_01385_, _01384_, _01382_);
  or _23273_ (_01386_, _01385_, _07056_);
  nor _23274_ (_01387_, _01386_, _01381_);
  and _23275_ (_01388_, _01387_, _01378_);
  and _23276_ (_01390_, _01388_, _12123_);
  nor _23277_ (_01391_, _01390_, _08330_);
  or _23278_ (_01393_, _01391_, p2_in[7]);
  not _23279_ (_01394_, _01391_);
  or _23280_ (_01396_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _23281_ (_01397_, _01396_, _01393_);
  and _23282_ (_01398_, _01397_, _01373_);
  and _23283_ (_01399_, _01322_, _01363_);
  or _23284_ (_01400_, _01391_, p3_in[7]);
  or _23285_ (_01401_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _23286_ (_01402_, _01401_, _01400_);
  and _23287_ (_01403_, _01402_, _01399_);
  or _23288_ (_01404_, _01403_, _01398_);
  and _23289_ (_01405_, _01363_, _01283_);
  or _23290_ (_01406_, _01391_, p0_in[7]);
  or _23291_ (_01407_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23292_ (_01408_, _01407_, _01406_);
  and _23293_ (_01409_, _01408_, _01405_);
  or _23294_ (_01410_, _01391_, p1_in[7]);
  or _23295_ (_01411_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _23296_ (_01412_, _01411_, _01410_);
  and _23297_ (_01413_, _01343_, _01363_);
  and _23298_ (_01414_, _01413_, _01412_);
  or _23299_ (_01415_, _01414_, _01409_);
  or _23300_ (_01416_, _01415_, _01404_);
  or _23301_ (_01417_, _01416_, _01371_);
  and _23302_ (_01418_, _01363_, _01280_);
  or _23303_ (_01419_, _12450_, _12313_);
  or _23304_ (_01420_, _01419_, _12261_);
  not _23305_ (_01421_, _01420_);
  and _23306_ (_01422_, _01421_, _01418_);
  and _23307_ (_01423_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _23308_ (_01424_, _01363_, _12261_);
  and _23309_ (_01425_, _01424_, _01362_);
  and _23310_ (_01426_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _23311_ (_01427_, _01426_, _01423_);
  or _23312_ (_01428_, _01427_, _01417_);
  or _23313_ (_01429_, _01428_, _01356_);
  nand _23314_ (_01430_, _01422_, _12690_);
  nand _23315_ (_01431_, _01285_, _01309_);
  or _23316_ (_01432_, _01431_, _07138_);
  and _23317_ (_01433_, _01432_, _01430_);
  or _23318_ (_01434_, _01433_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _23319_ (_01435_, _06010_);
  nor _23320_ (_01436_, _01323_, _01435_);
  nand _23321_ (_01437_, _01436_, _12455_);
  nand _23322_ (_01438_, _01425_, _08161_);
  and _23323_ (_01439_, _01438_, _01437_);
  and _23324_ (_01440_, _01439_, _12617_);
  and _23325_ (_01441_, _01440_, _01434_);
  and _23326_ (_01442_, _01441_, _01429_);
  not _23327_ (_01443_, _01441_);
  nor _23328_ (_01444_, _01297_, _01293_);
  nor _23329_ (_01445_, _01305_, _01301_);
  and _23330_ (_01446_, _01445_, _01444_);
  nor _23331_ (_01447_, _01313_, _01311_);
  nor _23332_ (_01448_, _01325_, _01319_);
  and _23333_ (_01449_, _01448_, _01447_);
  and _23334_ (_01450_, _01449_, _01446_);
  nor _23335_ (_01452_, _01346_, _01344_);
  nor _23336_ (_01453_, _01351_, _01349_);
  and _23337_ (_01454_, _01453_, _01452_);
  nor _23338_ (_01455_, _01333_, _01330_);
  nor _23339_ (_01456_, _01338_, _01336_);
  and _23340_ (_01457_, _01456_, _01455_);
  and _23341_ (_01458_, _01457_, _01454_);
  and _23342_ (_01460_, _01458_, _01450_);
  nor _23343_ (_01461_, _01425_, _01422_);
  nor _23344_ (_01462_, _01359_, _01286_);
  nor _23345_ (_01463_, _01368_, _01365_);
  and _23346_ (_01464_, _01463_, _01462_);
  nor _23347_ (_01466_, _01399_, _01373_);
  nor _23348_ (_01468_, _01413_, _01405_);
  and _23349_ (_01469_, _01468_, _01466_);
  and _23350_ (_01470_, _01469_, _01464_);
  and _23351_ (_01471_, _01470_, _01461_);
  and _23352_ (_01472_, _01471_, _01460_);
  or _23353_ (_01474_, _01472_, _01443_);
  and _23354_ (_01475_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _23355_ (_01476_, _01475_, _01442_);
  or _23356_ (_01477_, _01476_, _01287_);
  nand _23357_ (_01478_, _01287_, _06875_);
  and _23358_ (_01480_, _01478_, _05141_);
  and _23359_ (_01025_, _01480_, _01477_);
  and _23360_ (_01481_, _06004_, _05277_);
  and _23361_ (_01482_, _08484_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _23362_ (_01483_, _01482_, _05572_);
  or _23363_ (_01485_, _01483_, _01481_);
  or _23364_ (_01486_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _23365_ (_01487_, _01486_, _05141_);
  and _23366_ (_01027_, _01487_, _01485_);
  and _23367_ (_01488_, _06013_, _06207_);
  nand _23368_ (_01489_, _01488_, _05963_);
  or _23369_ (_01490_, _01488_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _23370_ (_01491_, _01490_, _01489_);
  or _23371_ (_01492_, _01491_, _06020_);
  nand _23372_ (_01493_, _06244_, _06020_);
  and _23373_ (_01494_, _01493_, _05141_);
  and _23374_ (_01030_, _01494_, _01492_);
  and _23375_ (_01495_, _06255_, _06207_);
  nand _23376_ (_01496_, _01495_, _05963_);
  or _23377_ (_01497_, _01495_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _23378_ (_01498_, _01497_, _06263_);
  and _23379_ (_01499_, _01498_, _01496_);
  nor _23380_ (_01501_, _06263_, _06244_);
  or _23381_ (_01502_, _01501_, _01499_);
  and _23382_ (_01032_, _01502_, _05141_);
  and _23383_ (_01504_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _23384_ (_01505_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _23385_ (_01506_, _01505_, _01504_);
  and _23386_ (_01507_, _01506_, _08355_);
  and _23387_ (_01508_, _08348_, _05522_);
  or _23388_ (_01509_, _01508_, _01507_);
  and _23389_ (_01149_, _01509_, _05141_);
  and _23390_ (_01510_, _06281_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _23391_ (_01512_, _06275_, _06179_);
  or _23392_ (_01513_, _01512_, _01510_);
  and _23393_ (_01183_, _01513_, _05141_);
  nor _23394_ (_01514_, _06121_, _06065_);
  and _23395_ (_01515_, _06065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _23396_ (_01517_, _01515_, _01514_);
  and _23397_ (_01389_, _01517_, _05141_);
  not _23398_ (_01518_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _23399_ (_01519_, _06089_, _05630_);
  or _23400_ (_01520_, _01519_, _01518_);
  nor _23401_ (_01521_, _06085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23402_ (_01522_, _01521_, _06093_);
  nand _23403_ (_01524_, _01522_, _01520_);
  or _23404_ (_01525_, _06094_, _05629_);
  and _23405_ (_01526_, _01525_, _01524_);
  or _23406_ (_01527_, _01526_, _06078_);
  not _23407_ (_01528_, _06076_);
  or _23408_ (_01529_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _05630_);
  or _23409_ (_01530_, _01529_, _01245_);
  and _23410_ (_01531_, _01530_, _01528_);
  and _23411_ (_01532_, _01531_, _01527_);
  and _23412_ (_01533_, _06076_, _05629_);
  or _23413_ (_01534_, _01533_, _06073_);
  or _23414_ (_01535_, _01534_, _01532_);
  or _23415_ (_01536_, _01529_, _06074_);
  and _23416_ (_01537_, _01536_, _01535_);
  or _23417_ (_01538_, _01537_, _06123_);
  and _23418_ (_01539_, _06102_, _05630_);
  or _23419_ (_01541_, _01539_, _01518_);
  and _23420_ (_01542_, _06100_, _05630_);
  nor _23421_ (_01544_, _01542_, _06105_);
  nand _23422_ (_01546_, _01544_, _01541_);
  or _23423_ (_01547_, _06106_, _05629_);
  and _23424_ (_01549_, _01547_, _01546_);
  or _23425_ (_01550_, _01549_, _06114_);
  not _23426_ (_01551_, _06112_);
  or _23427_ (_01552_, _01529_, _01237_);
  and _23428_ (_01554_, _01552_, _01551_);
  and _23429_ (_01555_, _01554_, _01550_);
  and _23430_ (_01556_, _06112_, _05629_);
  or _23431_ (_01557_, _01556_, _06109_);
  or _23432_ (_01558_, _01557_, _01555_);
  or _23433_ (_01559_, _01529_, _06110_);
  and _23434_ (_01560_, _01559_, _01558_);
  or _23435_ (_01561_, _01560_, _06134_);
  and _23436_ (_01562_, _01561_, _01538_);
  or _23437_ (_01563_, _01562_, _06065_);
  or _23438_ (_01565_, _01514_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _23439_ (_01566_, _01565_, _05141_);
  and _23440_ (_01392_, _01566_, _01563_);
  and _23441_ (_01567_, _06205_, _06620_);
  nand _23442_ (_01568_, _01567_, _05963_);
  or _23443_ (_01569_, _01567_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _23444_ (_01570_, _01569_, _05928_);
  and _23445_ (_01571_, _01570_, _01568_);
  nor _23446_ (_01572_, _05928_, _05560_);
  or _23447_ (_01573_, _01572_, _01571_);
  and _23448_ (_01395_, _01573_, _05141_);
  and _23449_ (_01451_, _11861_, _05141_);
  or _23450_ (_01574_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _05630_);
  and _23451_ (_01575_, _01574_, _06110_);
  or _23452_ (_01576_, _01575_, _06116_);
  and _23453_ (_01577_, _06105_, _05639_);
  not _23454_ (_01579_, _06115_);
  or _23455_ (_01580_, _01539_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23456_ (_01581_, _01580_, _01544_);
  or _23457_ (_01583_, _01581_, _01579_);
  or _23458_ (_01584_, _01583_, _01577_);
  and _23459_ (_01586_, _01584_, _01576_);
  and _23460_ (_01587_, _06109_, _05639_);
  or _23461_ (_01588_, _01587_, _06119_);
  or _23462_ (_01589_, _01588_, _01586_);
  or _23463_ (_01590_, _06120_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23464_ (_01591_, _01590_, _01589_);
  and _23465_ (_01592_, _01591_, _06123_);
  and _23466_ (_01593_, _01574_, _06074_);
  or _23467_ (_01594_, _01593_, _06081_);
  and _23468_ (_01595_, _06093_, _05639_);
  or _23469_ (_01596_, _01519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nand _23470_ (_01597_, _01596_, _01522_);
  nand _23471_ (_01598_, _01597_, _06080_);
  or _23472_ (_01599_, _01598_, _01595_);
  and _23473_ (_01600_, _01599_, _01594_);
  and _23474_ (_01601_, _06073_, _05639_);
  or _23475_ (_01602_, _01601_, _01600_);
  and _23476_ (_01603_, _01602_, _06097_);
  or _23477_ (_01604_, _01603_, _06065_);
  or _23478_ (_01605_, _01604_, _01592_);
  or _23479_ (_01606_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23480_ (_01607_, _01606_, _05141_);
  and _23481_ (_01459_, _01607_, _01605_);
  and _23482_ (_01608_, _06205_, _08469_);
  or _23483_ (_01609_, _01608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _23484_ (_01610_, _01609_, _05928_);
  nand _23485_ (_01611_, _01608_, _05963_);
  and _23486_ (_01612_, _01611_, _01610_);
  and _23487_ (_01613_, _05927_, _05522_);
  or _23488_ (_01614_, _01613_, _01612_);
  and _23489_ (_01465_, _01614_, _05141_);
  and _23490_ (_01467_, _06391_, _05141_);
  and _23491_ (_01473_, _13350_, _06065_);
  and _23492_ (_01615_, _06065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _23493_ (_01616_, _01615_, _01514_);
  and _23494_ (_01479_, _01616_, _05141_);
  nand _23495_ (_01617_, _06117_, _06141_);
  nor _23496_ (_01618_, _01617_, _06097_);
  and _23497_ (_01619_, _06065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor _23498_ (_01620_, _06093_, _06071_);
  not _23499_ (_01621_, _06081_);
  nor _23500_ (_01622_, _06091_, _01621_);
  and _23501_ (_01623_, _01622_, _01620_);
  and _23502_ (_01624_, _01623_, _06066_);
  or _23503_ (_01625_, _01624_, _01619_);
  or _23504_ (_01627_, _01625_, _01618_);
  and _23505_ (_01484_, _01627_, _05141_);
  or _23506_ (_01628_, _06093_, _06078_);
  and _23507_ (_01629_, _06091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23508_ (_01630_, _01629_, _01628_);
  and _23509_ (_01631_, _01630_, _01528_);
  and _23510_ (_01632_, _01631_, _01251_);
  nor _23511_ (_01633_, _06112_, _06109_);
  or _23512_ (_01634_, _06114_, _06105_);
  and _23513_ (_01635_, _06103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23514_ (_01636_, _01635_, _01634_);
  and _23515_ (_01637_, _01636_, _01633_);
  and _23516_ (_01638_, _01637_, _06133_);
  or _23517_ (_01639_, _01638_, _06065_);
  or _23518_ (_01640_, _01639_, _01632_);
  or _23519_ (_01641_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _23520_ (_01642_, _01641_, _05141_);
  and _23521_ (_01500_, _01642_, _01640_);
  nor _23522_ (_01643_, _06097_, _06065_);
  or _23523_ (_01644_, _01643_, _05630_);
  nand _23524_ (_01645_, _06247_, _06121_);
  and _23525_ (_01646_, _01645_, _05141_);
  and _23526_ (_01503_, _01646_, _01644_);
  or _23527_ (_01647_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23528_ (_01648_, _01647_, _05141_);
  or _23529_ (_01649_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23530_ (_01650_, _01649_, _06074_);
  or _23531_ (_01652_, _01650_, _06081_);
  and _23532_ (_01653_, _06089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23533_ (_01654_, _01653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor _23534_ (_01655_, _06085_, _05630_);
  nor _23535_ (_01656_, _01655_, _06093_);
  and _23536_ (_01657_, _01656_, _01654_);
  nand _23537_ (_01658_, _06093_, _05640_);
  nand _23538_ (_01659_, _01658_, _06080_);
  or _23539_ (_01660_, _01659_, _01657_);
  and _23540_ (_01661_, _01660_, _01652_);
  and _23541_ (_01662_, _06073_, _05640_);
  or _23542_ (_01663_, _01662_, _01661_);
  and _23543_ (_01664_, _01663_, _06097_);
  and _23544_ (_01665_, _01649_, _06110_);
  or _23545_ (_01666_, _01665_, _06116_);
  and _23546_ (_01667_, _06105_, _05640_);
  and _23547_ (_01668_, _06100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23548_ (_01669_, _01668_, _06105_);
  and _23549_ (_01670_, _06102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23550_ (_01671_, _01670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23551_ (_01672_, _01671_, _01669_);
  or _23552_ (_01673_, _01672_, _01579_);
  or _23553_ (_01674_, _01673_, _01667_);
  and _23554_ (_01675_, _01674_, _01666_);
  and _23555_ (_01676_, _06109_, _05640_);
  or _23556_ (_01677_, _01676_, _06119_);
  or _23557_ (_01678_, _01677_, _01675_);
  or _23558_ (_01679_, _06120_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23559_ (_01680_, _01679_, _01678_);
  and _23560_ (_01682_, _01680_, _06123_);
  or _23561_ (_01683_, _01682_, _01664_);
  or _23562_ (_01684_, _01683_, _06065_);
  and _23563_ (_01511_, _01684_, _01648_);
  not _23564_ (_01685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor _23565_ (_01686_, _01514_, _01685_);
  or _23566_ (_01687_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23567_ (_01688_, _01687_, _06074_);
  and _23568_ (_01689_, _01688_, _06097_);
  or _23569_ (_01690_, _01653_, _01685_);
  nand _23570_ (_01691_, _01690_, _01656_);
  or _23571_ (_01692_, _06094_, _05631_);
  and _23572_ (_01693_, _01692_, _01691_);
  or _23573_ (_01694_, _01693_, _06078_);
  or _23574_ (_01695_, _01687_, _01245_);
  and _23575_ (_01696_, _01695_, _01528_);
  and _23576_ (_01697_, _01696_, _01694_);
  and _23577_ (_01698_, _06076_, _05631_);
  or _23578_ (_01699_, _01698_, _06073_);
  or _23579_ (_01700_, _01699_, _01697_);
  and _23580_ (_01701_, _01700_, _01689_);
  or _23581_ (_01702_, _01670_, _01685_);
  nand _23582_ (_01703_, _01702_, _01669_);
  or _23583_ (_01704_, _06106_, _05631_);
  and _23584_ (_01705_, _01704_, _01703_);
  or _23585_ (_01706_, _01705_, _06114_);
  or _23586_ (_01707_, _01687_, _01237_);
  and _23587_ (_01708_, _01707_, _01551_);
  and _23588_ (_01709_, _01708_, _01706_);
  and _23589_ (_01710_, _06112_, _05631_);
  or _23590_ (_01711_, _01710_, _06109_);
  or _23591_ (_01712_, _01711_, _01709_);
  or _23592_ (_01713_, _01687_, _06110_);
  and _23593_ (_01714_, _01713_, _06133_);
  and _23594_ (_01715_, _01714_, _01712_);
  or _23595_ (_01716_, _01715_, _01701_);
  and _23596_ (_01717_, _01716_, _06066_);
  or _23597_ (_01718_, _01717_, _01686_);
  and _23598_ (_01516_, _01718_, _05141_);
  nand _23599_ (_01719_, _06247_, _06133_);
  and _23600_ (_01720_, _06247_, _06097_);
  or _23601_ (_01721_, _01720_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _23602_ (_01722_, _01721_, _05141_);
  and _23603_ (_01523_, _01722_, _01719_);
  nand _23604_ (_01723_, _06137_, _06133_);
  and _23605_ (_01724_, _06137_, _06097_);
  or _23606_ (_01725_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and _23607_ (_01726_, _01725_, _05141_);
  and _23608_ (_01540_, _01726_, _01723_);
  and _23609_ (_01727_, _06255_, _05288_);
  nand _23610_ (_01728_, _01727_, _05963_);
  or _23611_ (_01729_, _01727_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _23612_ (_01730_, _01729_, _06263_);
  and _23613_ (_01731_, _01730_, _01728_);
  nor _23614_ (_01732_, _06263_, _06178_);
  or _23615_ (_01734_, _01732_, _01731_);
  and _23616_ (_01543_, _01734_, _05141_);
  and _23617_ (_01735_, _06255_, _05210_);
  and _23618_ (_01736_, _01735_, _05963_);
  nor _23619_ (_01737_, _01735_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _23620_ (_01738_, _01737_, _01736_);
  nand _23621_ (_01739_, _01738_, _06263_);
  nand _23622_ (_01740_, _06262_, _05604_);
  and _23623_ (_01741_, _01740_, _05141_);
  and _23624_ (_01545_, _01741_, _01739_);
  and _23625_ (_01742_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _23626_ (_01743_, _01742_, _10380_);
  and _23627_ (_01744_, _01743_, _06255_);
  or _23628_ (_01745_, _01220_, _10375_);
  and _23629_ (_01746_, _01745_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _23630_ (_01747_, _01746_, _06262_);
  or _23631_ (_01748_, _01747_, _01744_);
  or _23632_ (_01749_, _06263_, _05522_);
  and _23633_ (_01750_, _01749_, _05141_);
  and _23634_ (_01548_, _01750_, _01748_);
  and _23635_ (_01751_, _08283_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _23636_ (_01752_, _01751_, _08281_);
  and _23637_ (_01753_, _01752_, _06255_);
  nand _23638_ (_01754_, _06255_, _05186_);
  and _23639_ (_01755_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _23640_ (_01757_, _01755_, _06262_);
  or _23641_ (_01759_, _01757_, _01753_);
  nand _23642_ (_01760_, _06262_, _06062_);
  and _23643_ (_01761_, _01760_, _05141_);
  and _23644_ (_01553_, _01761_, _01759_);
  and _23645_ (_01564_, _06532_, _05141_);
  and _23646_ (_01763_, _06283_, _06180_);
  and _23647_ (_01765_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _23648_ (_01766_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _23649_ (_01767_, _01766_, _06156_);
  or _23650_ (_01768_, _01767_, _01765_);
  or _23651_ (_01769_, _01768_, _01763_);
  and _23652_ (_01578_, _01769_, _05141_);
  or _23653_ (_01770_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _23654_ (_01771_, pc_log_change, _05411_);
  and _23655_ (_01772_, _01771_, _05141_);
  and _23656_ (_01582_, _01772_, _01770_);
  and _23657_ (_01773_, _06013_, _05288_);
  nand _23658_ (_01774_, _01773_, _05963_);
  or _23659_ (_01775_, _01773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _23660_ (_01776_, _01775_, _06021_);
  and _23661_ (_01777_, _01776_, _01774_);
  nor _23662_ (_01778_, _06178_, _06021_);
  or _23663_ (_01780_, _01778_, _01777_);
  and _23664_ (_01585_, _01780_, _05141_);
  or _23665_ (_01781_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand _23666_ (_01782_, _07619_, _06379_);
  and _23667_ (_01784_, _01782_, _05141_);
  and _23668_ (_01626_, _01784_, _01781_);
  nand _23669_ (_01785_, _06875_, _06624_);
  or _23670_ (_01786_, _06624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _23671_ (_01787_, _01786_, _05141_);
  and _23672_ (_01651_, _01787_, _01785_);
  and _23673_ (_01788_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _23674_ (_01789_, _01788_, _06683_);
  not _23675_ (_01790_, _01789_);
  and _23676_ (_01791_, _00626_, _08295_);
  nor _23677_ (_01792_, _01791_, _06685_);
  nor _23678_ (_01793_, _09785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  not _23679_ (_01794_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _23680_ (_01795_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01794_);
  and _23681_ (_01796_, _01795_, _01793_);
  nor _23682_ (_01797_, _01796_, _06686_);
  and _23683_ (_01798_, _01797_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _23684_ (_01799_, _01798_, _01792_);
  and _23685_ (_01800_, _01799_, _01790_);
  and _23686_ (_01801_, _01796_, _06685_);
  nor _23687_ (_01802_, _01801_, _01789_);
  not _23688_ (_01803_, _01802_);
  nand _23689_ (_01804_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _23690_ (_01805_, _01804_, _06715_);
  or _23691_ (_01681_, _01805_, _01800_);
  or _23692_ (_01806_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand _23693_ (_01807_, _07619_, _06403_);
  and _23694_ (_01808_, _01807_, _05141_);
  and _23695_ (_01733_, _01808_, _01806_);
  and _23696_ (_01809_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _23697_ (_01810_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _23698_ (_01811_, pc_log_change, _01810_);
  or _23699_ (_01812_, _01811_, _01809_);
  and _23700_ (_01756_, _01812_, _05141_);
  and _23701_ (_01813_, _06013_, _05210_);
  nand _23702_ (_01814_, _01813_, _05963_);
  or _23703_ (_01815_, _01813_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _23704_ (_01816_, _01815_, _01814_);
  or _23705_ (_01817_, _01816_, _06020_);
  nand _23706_ (_01818_, _06020_, _05604_);
  and _23707_ (_01819_, _01818_, _05141_);
  and _23708_ (_01758_, _01819_, _01817_);
  and _23709_ (_01820_, _10374_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _23710_ (_01821_, _01820_, _10380_);
  and _23711_ (_01822_, _01821_, _06013_);
  or _23712_ (_01823_, _10375_, _01200_);
  and _23713_ (_01825_, _01823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _23714_ (_01826_, _01825_, _06020_);
  or _23715_ (_01827_, _01826_, _01822_);
  or _23716_ (_01828_, _06021_, _05522_);
  and _23717_ (_01829_, _01828_, _05141_);
  and _23718_ (_01762_, _01829_, _01827_);
  nor _23719_ (_01830_, _08282_, _06104_);
  or _23720_ (_01831_, _01830_, _08281_);
  and _23721_ (_01832_, _01831_, _06013_);
  nand _23722_ (_01833_, _06013_, _05186_);
  and _23723_ (_01834_, _01833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _23724_ (_01835_, _01834_, _06020_);
  or _23725_ (_01836_, _01835_, _01832_);
  nand _23726_ (_01837_, _06062_, _06020_);
  and _23727_ (_01838_, _01837_, _05141_);
  and _23728_ (_01764_, _01838_, _01836_);
  and _23729_ (_01839_, _10346_, _06032_);
  nand _23730_ (_01840_, _01839_, _05963_);
  or _23731_ (_01841_, _01839_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _23732_ (_01843_, _01841_, _10355_);
  nand _23733_ (_01844_, _01843_, _01840_);
  nand _23734_ (_01845_, _01844_, _11860_);
  and _23735_ (_01779_, _01845_, _05141_);
  and _23736_ (_01846_, _06293_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _23737_ (_01847_, _06766_, _06550_);
  or _23738_ (_01848_, _13288_, _12117_);
  or _23739_ (_01849_, _01848_, _01847_);
  or _23740_ (_01850_, _01374_, _06996_);
  not _23741_ (_01851_, _07054_);
  or _23742_ (_01852_, _01851_, _06772_);
  or _23743_ (_01854_, _01852_, _01850_);
  or _23744_ (_01855_, _01854_, _01849_);
  or _23745_ (_01856_, _01855_, _06780_);
  and _23746_ (_01857_, _07069_, _06546_);
  or _23747_ (_01858_, _01383_, _01857_);
  or _23748_ (_01859_, _11431_, _06980_);
  or _23749_ (_01861_, _01859_, _01858_);
  or _23750_ (_01862_, _01861_, _06764_);
  and _23751_ (_01864_, _06565_, _06420_);
  or _23752_ (_01865_, _12114_, _07037_);
  or _23753_ (_01866_, _01865_, _01864_);
  and _23754_ (_01867_, _06556_, _06536_);
  and _23755_ (_01869_, _06552_, _06536_);
  or _23756_ (_01870_, _01869_, _01867_);
  and _23757_ (_01872_, _06755_, _07053_);
  or _23758_ (_01873_, _01872_, _01870_);
  or _23759_ (_01875_, _01873_, _01866_);
  or _23760_ (_01876_, _01875_, _01862_);
  or _23761_ (_01877_, _01876_, _01856_);
  and _23762_ (_01878_, _01877_, _06296_);
  or _23763_ (_01783_, _01878_, _01846_);
  or _23764_ (_01879_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand _23765_ (_01880_, _07619_, _06514_);
  and _23766_ (_01881_, _01880_, _05141_);
  and _23767_ (_01824_, _01881_, _01879_);
  and _23768_ (_01882_, _05563_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _23769_ (_01884_, _06290_, _05523_);
  or _23770_ (_01885_, _01884_, _01882_);
  and _23771_ (_01842_, _01885_, _05141_);
  nand _23772_ (_01887_, _06743_, _05960_);
  and _23773_ (_01889_, _08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _23774_ (_01891_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _23775_ (_01892_, _01891_, _01889_);
  or _23776_ (_01893_, _01892_, _06743_);
  and _23777_ (_01894_, _01893_, _05141_);
  and _23778_ (_01853_, _01894_, _01887_);
  or _23779_ (_01895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _23780_ (_01896_, _01895_, _11458_);
  and _23781_ (_01897_, _05922_, _06008_);
  not _23782_ (_01898_, _06008_);
  nand _23783_ (_01899_, _01898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _23784_ (_01900_, _01899_, _11458_);
  or _23785_ (_01901_, _01900_, _01897_);
  and _23786_ (_01902_, _01901_, _01896_);
  or _23787_ (_01903_, _01902_, _11462_);
  nand _23788_ (_01904_, _11462_, _05960_);
  and _23789_ (_01905_, _01904_, _05141_);
  and _23790_ (_01860_, _01905_, _01903_);
  nor _23791_ (_01906_, _11727_, _11651_);
  and _23792_ (_01907_, _11727_, _08439_);
  and _23793_ (_01908_, _08462_, _06726_);
  and _23794_ (_01909_, _01908_, _08457_);
  and _23795_ (_01910_, _01909_, _01907_);
  or _23796_ (_01911_, _01910_, _01906_);
  and _23797_ (_01863_, _01911_, _05141_);
  nand _23798_ (_01912_, _11726_, _05960_);
  or _23799_ (_01913_, _11830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _23800_ (_01914_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _23801_ (_01915_, _01914_, _08439_);
  nand _23802_ (_01916_, _01915_, _08457_);
  and _23803_ (_01918_, _01916_, _01913_);
  or _23804_ (_01919_, _01918_, _08463_);
  nor _23805_ (_01920_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor _23806_ (_01922_, _01920_, _08471_);
  and _23807_ (_01923_, _01922_, _01919_);
  nor _23808_ (_01924_, _11726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor _23809_ (_01925_, _01924_, _11727_);
  or _23810_ (_01926_, _01925_, _01923_);
  and _23811_ (_01928_, _01926_, _05141_);
  and _23812_ (_01868_, _01928_, _01912_);
  nor _23813_ (_01929_, _11902_, _05960_);
  and _23814_ (_01930_, _11753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _23815_ (_01931_, _01930_, _08457_);
  nor _23816_ (_01932_, _08452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor _23817_ (_01933_, _01932_, _08453_);
  or _23818_ (_01934_, _01933_, _13159_);
  or _23819_ (_01935_, _01934_, _01931_);
  or _23820_ (_01936_, _08439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _23821_ (_01937_, _01936_, _01935_);
  or _23822_ (_01938_, _01937_, _08463_);
  nor _23823_ (_01939_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor _23824_ (_01940_, _01939_, _08471_);
  and _23825_ (_01941_, _01940_, _01938_);
  or _23826_ (_01942_, _01941_, _08478_);
  or _23827_ (_01943_, _01942_, _01929_);
  or _23828_ (_01944_, _08479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _23829_ (_01945_, _01944_, _05141_);
  and _23830_ (_01871_, _01945_, _01943_);
  not _23831_ (_01946_, _08457_);
  and _23832_ (_01947_, _01907_, _08460_);
  nand _23833_ (_01948_, _01947_, _01946_);
  or _23834_ (_01949_, _01947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _23835_ (_01950_, _01949_, _05141_);
  and _23836_ (_01874_, _01950_, _01948_);
  and _23837_ (_01883_, t2_i, _05141_);
  nand _23838_ (_01951_, _06738_, _05960_);
  and _23839_ (_01952_, _06730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _23840_ (_01953_, _06728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _23841_ (_01954_, _01953_, _01952_);
  or _23842_ (_01955_, _01954_, _06738_);
  and _23843_ (_01956_, _01955_, _06745_);
  and _23844_ (_01957_, _01956_, _01951_);
  and _23845_ (_01958_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _23846_ (_01959_, _01958_, _01957_);
  and _23847_ (_01886_, _01959_, _05141_);
  and _23848_ (_01888_, t2ex_i, _05141_);
  and _23849_ (_01890_, _06531_, _05141_);
  nor _23850_ (_01960_, t2ex_i, rst);
  and _23851_ (_01917_, _01960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor _23852_ (_01961_, t2_i, rst);
  and _23853_ (_01921_, _01961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and _23854_ (_01962_, _06283_, _05523_);
  and _23855_ (_01963_, _05303_, _05297_);
  or _23856_ (_01964_, _01963_, _05299_);
  and _23857_ (_01965_, _01964_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _23858_ (_01966_, _01965_, _01962_);
  and _23859_ (_01927_, _01966_, _05141_);
  and _23860_ (_01967_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _23861_ (_01968_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _23862_ (_01969_, pc_log_change, _01968_);
  or _23863_ (_01970_, _01969_, _01967_);
  and _23864_ (_02067_, _01970_, _05141_);
  or _23865_ (_01971_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _23866_ (_01972_, pc_log_change, _05436_);
  and _23867_ (_01973_, _01972_, _05141_);
  and _23868_ (_02103_, _01973_, _01971_);
  nor _23869_ (_01974_, _05560_, _08484_);
  and _23870_ (_01975_, _08484_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _23871_ (_01976_, _01975_, _01974_);
  or _23872_ (_01977_, _01976_, _05572_);
  or _23873_ (_01978_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _23874_ (_01979_, _01978_, _05141_);
  and _23875_ (_02137_, _01979_, _01977_);
  nand _23876_ (_01980_, _06678_, _06244_);
  or _23877_ (_01981_, _06678_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _23878_ (_01982_, _01981_, _05141_);
  and _23879_ (_02194_, _01982_, _01980_);
  or _23880_ (_01983_, _06975_, _07138_);
  nor _23881_ (_01984_, _07169_, _06875_);
  and _23882_ (_01985_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _23883_ (_01986_, _01985_, _06619_);
  or _23884_ (_01987_, _01986_, _01984_);
  and _23885_ (_01988_, _01987_, _05141_);
  and _23886_ (_02221_, _01988_, _01983_);
  and _23887_ (_01989_, _00690_, _10407_);
  nand _23888_ (_01990_, _01989_, _05963_);
  or _23889_ (_01991_, _01989_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _23890_ (_01992_, _01991_, _05647_);
  and _23891_ (_01993_, _01992_, _01990_);
  not _23892_ (_01994_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor _23893_ (_01995_, _05646_, _01994_);
  nand _23894_ (_01996_, _00698_, _07200_);
  or _23895_ (_01997_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _23896_ (_01998_, _01997_, _05925_);
  and _23897_ (_01999_, _01998_, _01996_);
  or _23898_ (_02000_, _01999_, _01995_);
  or _23899_ (_02001_, _02000_, _01993_);
  and _23900_ (_02394_, _02001_, _05141_);
  nand _23901_ (_02002_, _00690_, _08283_);
  and _23902_ (_02003_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _23903_ (_02004_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _23904_ (_02005_, _02004_, _10356_);
  and _23905_ (_02006_, _02005_, _00690_);
  or _23906_ (_02007_, _02006_, _02003_);
  and _23907_ (_02008_, _02007_, _05647_);
  and _23908_ (_02009_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _23909_ (_02010_, _00698_, _06617_);
  or _23910_ (_02011_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _23911_ (_02012_, _02011_, _05925_);
  and _23912_ (_02013_, _02012_, _02010_);
  or _23913_ (_02014_, _02013_, _02009_);
  or _23914_ (_02015_, _02014_, _02008_);
  and _23915_ (_02397_, _02015_, _05141_);
  nor _23916_ (_02429_, _12304_, rst);
  nand _23917_ (_02431_, _12463_, _05141_);
  and _23918_ (_02016_, _10342_, _06009_);
  and _23919_ (_02017_, _02016_, _05210_);
  nand _23920_ (_02018_, _02017_, _05963_);
  or _23921_ (_02019_, _02017_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _23922_ (_02020_, _02019_, _05647_);
  and _23923_ (_02021_, _02020_, _02018_);
  and _23924_ (_02022_, _06017_, _05272_);
  and _23925_ (_02023_, _02022_, _06703_);
  not _23926_ (_02024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _23927_ (_02025_, _02022_, _02024_);
  or _23928_ (_02026_, _02025_, _02023_);
  and _23929_ (_02027_, _02026_, _05925_);
  nor _23930_ (_02028_, _05646_, _02024_);
  or _23931_ (_02029_, _02028_, rst);
  or _23932_ (_02030_, _02029_, _02027_);
  or _23933_ (_02493_, _02030_, _02021_);
  and _23934_ (_02031_, _01257_, _06207_);
  nand _23935_ (_02032_, _02031_, _05963_);
  or _23936_ (_02033_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _23937_ (_02034_, _02033_, _05647_);
  and _23938_ (_02035_, _02034_, _02032_);
  nor _23939_ (_02036_, _01264_, _06244_);
  and _23940_ (_02037_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _23941_ (_02038_, _02037_, _02036_);
  and _23942_ (_02039_, _02038_, _05925_);
  and _23943_ (_02040_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _23944_ (_02041_, _02040_, rst);
  or _23945_ (_02042_, _02041_, _02039_);
  or _23946_ (_02495_, _02042_, _02035_);
  and _23947_ (_02043_, _10342_, _06202_);
  and _23948_ (_02044_, _02043_, _06620_);
  nand _23949_ (_02045_, _02044_, _05963_);
  or _23950_ (_02046_, _02044_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _23951_ (_02047_, _02046_, _05647_);
  and _23952_ (_02048_, _02047_, _02045_);
  and _23953_ (_02049_, _08241_, _05272_);
  nand _23954_ (_02050_, _02049_, _05560_);
  or _23955_ (_02051_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _23956_ (_02052_, _02051_, _05925_);
  and _23957_ (_02053_, _02052_, _02050_);
  and _23958_ (_02054_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _23959_ (_02055_, _02054_, rst);
  or _23960_ (_02056_, _02055_, _02053_);
  or _23961_ (_02499_, _02056_, _02048_);
  or _23962_ (_02057_, _01264_, _05922_);
  or _23963_ (_02058_, _01263_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _23964_ (_02059_, _02058_, _05647_);
  and _23965_ (_02060_, _02059_, _02057_);
  and _23966_ (_02061_, _01263_, _06703_);
  not _23967_ (_02062_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _23968_ (_02063_, _01263_, _02062_);
  or _23969_ (_02064_, _02063_, _02061_);
  and _23970_ (_02065_, _02064_, _05925_);
  nor _23971_ (_02066_, _05646_, _02062_);
  or _23972_ (_02068_, _02066_, rst);
  or _23973_ (_02069_, _02068_, _02065_);
  or _23974_ (_02501_, _02069_, _02060_);
  and _23975_ (_02070_, _06878_, _06202_);
  nand _23976_ (_02071_, _02070_, _05186_);
  and _23977_ (_02072_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _23978_ (_02073_, _08283_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _23979_ (_02074_, _02073_, _08281_);
  and _23980_ (_02075_, _02074_, _02070_);
  or _23981_ (_02076_, _02075_, _02072_);
  and _23982_ (_02077_, _02076_, _05647_);
  and _23983_ (_02078_, _05649_, _05272_);
  nand _23984_ (_02079_, _02078_, _06062_);
  or _23985_ (_02080_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _23986_ (_02081_, _02080_, _05925_);
  and _23987_ (_02082_, _02081_, _02079_);
  and _23988_ (_02083_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _23989_ (_02084_, _02083_, rst);
  or _23990_ (_02085_, _02084_, _02082_);
  or _23991_ (_02502_, _02085_, _02077_);
  not _23992_ (_02086_, _02078_);
  or _23993_ (_02087_, _02086_, _05922_);
  or _23994_ (_02088_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _23995_ (_02089_, _02088_, _05647_);
  and _23996_ (_02090_, _02089_, _02087_);
  nand _23997_ (_02091_, _02078_, _05604_);
  and _23998_ (_02092_, _02088_, _05925_);
  and _23999_ (_02093_, _02092_, _02091_);
  not _24000_ (_02094_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _24001_ (_02095_, _05646_, _02094_);
  or _24002_ (_02096_, _02095_, rst);
  or _24003_ (_02097_, _02096_, _02093_);
  or _24004_ (_02504_, _02097_, _02090_);
  and _24005_ (_02098_, _02016_, _10407_);
  nand _24006_ (_02099_, _02098_, _05963_);
  or _24007_ (_02100_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _24008_ (_02101_, _02100_, _05647_);
  and _24009_ (_02102_, _02101_, _02099_);
  and _24010_ (_02104_, _02022_, _06004_);
  not _24011_ (_02105_, _02022_);
  and _24012_ (_02106_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _24013_ (_02107_, _02106_, _02104_);
  and _24014_ (_02108_, _02107_, _05925_);
  and _24015_ (_02109_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _24016_ (_02110_, _02109_, rst);
  or _24017_ (_02111_, _02110_, _02108_);
  or _24018_ (_02517_, _02111_, _02102_);
  and _24019_ (_02112_, _01257_, _10407_);
  nand _24020_ (_02113_, _02112_, _05963_);
  or _24021_ (_02114_, _02112_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _24022_ (_02115_, _02114_, _05647_);
  and _24023_ (_02116_, _02115_, _02113_);
  and _24024_ (_02117_, _01263_, _06004_);
  and _24025_ (_02118_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _24026_ (_02119_, _02118_, _02117_);
  and _24027_ (_02120_, _02119_, _05925_);
  and _24028_ (_02121_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _24029_ (_02122_, _02121_, rst);
  or _24030_ (_02123_, _02122_, _02120_);
  or _24031_ (_02519_, _02123_, _02116_);
  and _24032_ (_02124_, _02043_, _06207_);
  nand _24033_ (_02125_, _02124_, _05963_);
  or _24034_ (_02126_, _02124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _24035_ (_02127_, _02126_, _05647_);
  and _24036_ (_02128_, _02127_, _02125_);
  nand _24037_ (_02129_, _02049_, _06244_);
  or _24038_ (_02130_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _24039_ (_02131_, _02130_, _05925_);
  and _24040_ (_02132_, _02131_, _02129_);
  and _24041_ (_02133_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _24042_ (_02134_, _02133_, rst);
  or _24043_ (_02135_, _02134_, _02132_);
  or _24044_ (_02522_, _02135_, _02128_);
  and _24045_ (_02136_, _02043_, _05288_);
  nand _24046_ (_02138_, _02136_, _05963_);
  or _24047_ (_02139_, _02136_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _24048_ (_02140_, _02139_, _05647_);
  and _24049_ (_02141_, _02140_, _02138_);
  nand _24050_ (_02142_, _02049_, _06178_);
  or _24051_ (_02143_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _24052_ (_02144_, _02143_, _05925_);
  and _24053_ (_02145_, _02144_, _02142_);
  and _24054_ (_02146_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _24055_ (_02147_, _02146_, rst);
  or _24056_ (_02148_, _02147_, _02145_);
  or _24057_ (_02523_, _02148_, _02141_);
  and _24058_ (_02149_, _02043_, _08469_);
  nand _24059_ (_02150_, _02149_, _05963_);
  or _24060_ (_02151_, _02149_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24061_ (_02152_, _02151_, _05647_);
  and _24062_ (_02153_, _02152_, _02150_);
  not _24063_ (_02154_, _02049_);
  or _24064_ (_02155_, _02154_, _05522_);
  or _24065_ (_02156_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24066_ (_02157_, _02156_, _05925_);
  and _24067_ (_02158_, _02157_, _02155_);
  and _24068_ (_02159_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _24069_ (_02160_, _02159_, rst);
  or _24070_ (_02161_, _02160_, _02158_);
  or _24071_ (_02525_, _02161_, _02153_);
  nand _24072_ (_02162_, _02070_, _08283_);
  and _24073_ (_02163_, _02162_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _24074_ (_02164_, _05287_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _24075_ (_02165_, _02164_, _10356_);
  and _24076_ (_02166_, _02165_, _02070_);
  or _24077_ (_02167_, _02166_, _02163_);
  and _24078_ (_02168_, _02167_, _05647_);
  nand _24079_ (_02169_, _02078_, _05560_);
  or _24080_ (_02170_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _24081_ (_02171_, _02170_, _05925_);
  and _24082_ (_02172_, _02171_, _02169_);
  and _24083_ (_02173_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _24084_ (_02174_, _02173_, rst);
  or _24085_ (_02175_, _02174_, _02172_);
  or _24086_ (_02526_, _02175_, _02168_);
  and _24087_ (_02176_, _02070_, _10407_);
  nand _24088_ (_02177_, _02176_, _05963_);
  or _24089_ (_02178_, _02176_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24090_ (_02179_, _02178_, _05647_);
  and _24091_ (_02180_, _02179_, _02177_);
  or _24092_ (_02181_, _02086_, _06004_);
  or _24093_ (_02182_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24094_ (_02183_, _02182_, _05925_);
  and _24095_ (_02184_, _02183_, _02181_);
  and _24096_ (_02185_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _24097_ (_02186_, _02185_, rst);
  or _24098_ (_02187_, _02186_, _02184_);
  or _24099_ (_02529_, _02187_, _02180_);
  and _24100_ (_02188_, _01257_, _08469_);
  nand _24101_ (_02189_, _02188_, _05963_);
  or _24102_ (_02190_, _02188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _24103_ (_02191_, _02190_, _05647_);
  and _24104_ (_02192_, _02191_, _02189_);
  and _24105_ (_02193_, _01263_, _05522_);
  and _24106_ (_02195_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _24107_ (_02196_, _02195_, _02193_);
  and _24108_ (_02197_, _02196_, _05925_);
  and _24109_ (_02198_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _24110_ (_02199_, _02198_, rst);
  or _24111_ (_02200_, _02199_, _02197_);
  or _24112_ (_02613_, _02200_, _02192_);
  and _24113_ (_02201_, _01257_, _06032_);
  nand _24114_ (_02202_, _02201_, _05963_);
  or _24115_ (_02203_, _02201_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _24116_ (_02204_, _02203_, _05647_);
  and _24117_ (_02205_, _02204_, _02202_);
  nor _24118_ (_02206_, _01264_, _06062_);
  and _24119_ (_02207_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _24120_ (_02208_, _02207_, _02206_);
  and _24121_ (_02209_, _02208_, _05925_);
  and _24122_ (_02210_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _24123_ (_02211_, _02210_, rst);
  or _24124_ (_02212_, _02211_, _02209_);
  or _24125_ (_02615_, _02212_, _02205_);
  and _24126_ (_02213_, _01257_, _06620_);
  nand _24127_ (_02214_, _02213_, _05963_);
  or _24128_ (_02215_, _02213_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _24129_ (_02216_, _02215_, _05647_);
  and _24130_ (_02217_, _02216_, _02214_);
  nor _24131_ (_02218_, _01264_, _05560_);
  and _24132_ (_02219_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _24133_ (_02220_, _02219_, _02218_);
  and _24134_ (_02222_, _02220_, _05925_);
  and _24135_ (_02223_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _24136_ (_02224_, _02223_, rst);
  or _24137_ (_02225_, _02224_, _02222_);
  or _24138_ (_02634_, _02225_, _02217_);
  or _24139_ (_02226_, _02154_, _05922_);
  or _24140_ (_02227_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _24141_ (_02228_, _02227_, _05647_);
  and _24142_ (_02229_, _02228_, _02226_);
  nand _24143_ (_02230_, _02049_, _05604_);
  and _24144_ (_02231_, _02227_, _05925_);
  and _24145_ (_02232_, _02231_, _02230_);
  not _24146_ (_02233_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _24147_ (_02234_, _05646_, _02233_);
  or _24148_ (_02235_, _02234_, rst);
  or _24149_ (_02236_, _02235_, _02232_);
  or _24150_ (_02635_, _02236_, _02229_);
  and _24151_ (_02237_, _02016_, _06032_);
  nand _24152_ (_02238_, _02237_, _05963_);
  or _24153_ (_02239_, _02237_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _24154_ (_02240_, _02239_, _05647_);
  and _24155_ (_02241_, _02240_, _02238_);
  nor _24156_ (_02242_, _02105_, _06062_);
  and _24157_ (_02243_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _24158_ (_02244_, _02243_, _02242_);
  and _24159_ (_02245_, _02244_, _05925_);
  and _24160_ (_02246_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _24161_ (_02247_, _02246_, rst);
  or _24162_ (_02248_, _02247_, _02245_);
  or _24163_ (_02638_, _02248_, _02241_);
  and _24164_ (_02249_, _02016_, _06620_);
  nand _24165_ (_02250_, _02249_, _05963_);
  or _24166_ (_02251_, _02249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _24167_ (_02252_, _02251_, _05647_);
  and _24168_ (_02253_, _02252_, _02250_);
  nor _24169_ (_02254_, _02105_, _05560_);
  and _24170_ (_02255_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _24171_ (_02256_, _02255_, _02254_);
  and _24172_ (_02257_, _02256_, _05925_);
  and _24173_ (_02258_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _24174_ (_02259_, _02258_, rst);
  or _24175_ (_02260_, _02259_, _02257_);
  or _24176_ (_02640_, _02260_, _02253_);
  and _24177_ (_02261_, _05649_, _05276_);
  nand _24178_ (_02262_, _02261_, _05963_);
  or _24179_ (_02263_, _02261_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _24180_ (_02264_, _02263_, _05647_);
  and _24181_ (_02265_, _02264_, _02262_);
  nand _24182_ (_02266_, _02078_, _06178_);
  or _24183_ (_02267_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _24184_ (_02268_, _02267_, _05925_);
  and _24185_ (_02269_, _02268_, _02266_);
  and _24186_ (_02270_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _24187_ (_02271_, _02270_, rst);
  or _24188_ (_02272_, _02271_, _02269_);
  or _24189_ (_02658_, _02272_, _02265_);
  and _24190_ (_02273_, _02070_, _06207_);
  nand _24191_ (_02274_, _02273_, _05963_);
  or _24192_ (_02275_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _24193_ (_02276_, _02275_, _05647_);
  and _24194_ (_02277_, _02276_, _02274_);
  nand _24195_ (_02278_, _02078_, _06244_);
  or _24196_ (_02279_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _24197_ (_02280_, _02279_, _05925_);
  and _24198_ (_02281_, _02280_, _02278_);
  and _24199_ (_02282_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _24200_ (_02283_, _02282_, rst);
  or _24201_ (_02284_, _02283_, _02281_);
  or _24202_ (_02661_, _02284_, _02277_);
  and _24203_ (_02285_, _02070_, _08469_);
  nand _24204_ (_02286_, _02285_, _05963_);
  or _24205_ (_02287_, _02285_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _24206_ (_02288_, _02287_, _05647_);
  and _24207_ (_02289_, _02288_, _02286_);
  or _24208_ (_02290_, _02086_, _05522_);
  or _24209_ (_02291_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _24210_ (_02292_, _02291_, _05925_);
  and _24211_ (_02293_, _02292_, _02290_);
  and _24212_ (_02294_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _24213_ (_02295_, _02294_, rst);
  or _24214_ (_02296_, _02295_, _02293_);
  or _24215_ (_02664_, _02296_, _02289_);
  and _24216_ (_02297_, _01257_, _05288_);
  nand _24217_ (_02298_, _02297_, _05963_);
  or _24218_ (_02299_, _02297_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _24219_ (_02300_, _02299_, _05647_);
  and _24220_ (_02301_, _02300_, _02298_);
  nor _24221_ (_02302_, _01264_, _06178_);
  and _24222_ (_02303_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _24223_ (_02304_, _02303_, _02302_);
  and _24224_ (_02305_, _02304_, _05925_);
  and _24225_ (_02306_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _24226_ (_02307_, _02306_, rst);
  or _24227_ (_02308_, _02307_, _02305_);
  or _24228_ (_02666_, _02308_, _02301_);
  and _24229_ (_02309_, _02043_, _10407_);
  nand _24230_ (_02310_, _02309_, _05963_);
  or _24231_ (_02311_, _02309_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _24232_ (_02312_, _02311_, _05647_);
  and _24233_ (_02313_, _02312_, _02310_);
  or _24234_ (_02314_, _02154_, _06004_);
  or _24235_ (_02315_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _24236_ (_02316_, _02315_, _05925_);
  and _24237_ (_02317_, _02316_, _02314_);
  and _24238_ (_02318_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _24239_ (_02319_, _02318_, rst);
  or _24240_ (_02320_, _02319_, _02317_);
  or _24241_ (_02668_, _02320_, _02313_);
  and _24242_ (_02321_, _02043_, _06032_);
  nand _24243_ (_02322_, _02321_, _05963_);
  or _24244_ (_02323_, _02321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _24245_ (_02324_, _02323_, _05647_);
  and _24246_ (_02325_, _02324_, _02322_);
  nand _24247_ (_02326_, _02049_, _06062_);
  or _24248_ (_02327_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _24249_ (_02328_, _02327_, _05925_);
  and _24250_ (_02329_, _02328_, _02326_);
  and _24251_ (_02330_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _24252_ (_02331_, _02330_, rst);
  or _24253_ (_02332_, _02331_, _02329_);
  or _24254_ (_02670_, _02332_, _02325_);
  and _24255_ (_02333_, _02016_, _05288_);
  nand _24256_ (_02334_, _02333_, _05963_);
  or _24257_ (_02335_, _02333_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _24258_ (_02336_, _02335_, _05647_);
  and _24259_ (_02337_, _02336_, _02334_);
  nor _24260_ (_02338_, _02105_, _06178_);
  and _24261_ (_02339_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _24262_ (_02340_, _02339_, _02338_);
  and _24263_ (_02341_, _02340_, _05925_);
  and _24264_ (_02342_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _24265_ (_02343_, _02342_, rst);
  or _24266_ (_02344_, _02343_, _02341_);
  or _24267_ (_02672_, _02344_, _02337_);
  and _24268_ (_02345_, _02016_, _06207_);
  nand _24269_ (_02346_, _02345_, _05963_);
  or _24270_ (_02347_, _02345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _24271_ (_02348_, _02347_, _05647_);
  and _24272_ (_02349_, _02348_, _02346_);
  nor _24273_ (_02350_, _02105_, _06244_);
  and _24274_ (_02351_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _24275_ (_02352_, _02351_, _02350_);
  and _24276_ (_02353_, _02352_, _05925_);
  and _24277_ (_02354_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _24278_ (_02355_, _02354_, rst);
  or _24279_ (_02356_, _02355_, _02353_);
  or _24280_ (_02677_, _02356_, _02349_);
  and _24281_ (_02357_, _02016_, _08469_);
  nand _24282_ (_02358_, _02357_, _05963_);
  or _24283_ (_02359_, _02357_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _24284_ (_02360_, _02359_, _05647_);
  and _24285_ (_02361_, _02360_, _02358_);
  and _24286_ (_02362_, _02022_, _05522_);
  and _24287_ (_02363_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _24288_ (_02364_, _02363_, _02362_);
  and _24289_ (_02365_, _02364_, _05925_);
  and _24290_ (_02366_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _24291_ (_02367_, _02366_, rst);
  or _24292_ (_02368_, _02367_, _02365_);
  or _24293_ (_02679_, _02368_, _02361_);
  or _24294_ (_02369_, _05277_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nand _24295_ (_02370_, _06178_, _05277_);
  and _24296_ (_02371_, _02370_, _02369_);
  or _24297_ (_02372_, _02371_, _05572_);
  or _24298_ (_02373_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _24299_ (_02374_, _02373_, _05141_);
  and _24300_ (_02698_, _02374_, _02372_);
  and _24301_ (_02375_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _24302_ (_02376_, pc_log_change, _13154_);
  or _24303_ (_02377_, _02376_, _02375_);
  and _24304_ (_02701_, _02377_, _05141_);
  or _24305_ (_02378_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not _24306_ (_02379_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _24307_ (_02380_, pc_log_change, _02379_);
  and _24308_ (_02381_, _02380_, _05141_);
  and _24309_ (_02705_, _02381_, _02378_);
  and _24310_ (_02382_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not _24311_ (_02383_, pc_log_change);
  and _24312_ (_02384_, _02383_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or _24313_ (_02385_, _02384_, _02382_);
  and _24314_ (_02710_, _02385_, _05141_);
  or _24315_ (_02386_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nand _24316_ (_02387_, pc_log_change, _01968_);
  and _24317_ (_02388_, _02387_, _05141_);
  and _24318_ (_02713_, _02388_, _02386_);
  and _24319_ (_02389_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _24320_ (_02390_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _24321_ (_02391_, pc_log_change, _02390_);
  or _24322_ (_02392_, _02391_, _02389_);
  and _24323_ (_02715_, _02392_, _05141_);
  and _24324_ (_02393_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _24325_ (_02395_, pc_log_change, _02379_);
  or _24326_ (_02396_, _02395_, _02393_);
  and _24327_ (_02723_, _02396_, _05141_);
  and _24328_ (_02398_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not _24329_ (_02399_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _24330_ (_02400_, pc_log_change, _02399_);
  or _24331_ (_02401_, _02400_, _02398_);
  and _24332_ (_02726_, _02401_, _05141_);
  and _24333_ (_02402_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _24334_ (_02403_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _24335_ (_02404_, pc_log_change, _02403_);
  or _24336_ (_02405_, _02404_, _02402_);
  and _24337_ (_02730_, _02405_, _05141_);
  and _24338_ (_02406_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _24339_ (_02407_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _24340_ (_02408_, pc_log_change, _02407_);
  or _24341_ (_02409_, _02408_, _02406_);
  and _24342_ (_02734_, _02409_, _05141_);
  and _24343_ (_02410_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _24344_ (_02411_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _24345_ (_02412_, pc_log_change, _02411_);
  or _24346_ (_02413_, _02412_, _02410_);
  and _24347_ (_02738_, _02413_, _05141_);
  and _24348_ (_02414_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _24349_ (_02415_, _02383_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or _24350_ (_02416_, _02415_, _02414_);
  and _24351_ (_02759_, _02416_, _05141_);
  and _24352_ (_02417_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _24353_ (_02418_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _24354_ (_02419_, pc_log_change, _02418_);
  or _24355_ (_02420_, _02419_, _02417_);
  and _24356_ (_02760_, _02420_, _05141_);
  or _24357_ (_02421_, _06363_, _07117_);
  or _24358_ (_02422_, _06270_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _24359_ (_02423_, _02422_, _05141_);
  and _24360_ (_02768_, _02423_, _02421_);
  and _24361_ (_02424_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _24362_ (_02425_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _24363_ (_02426_, pc_log_change, _02425_);
  or _24364_ (_02427_, _02426_, _02424_);
  and _24365_ (_02771_, _02427_, _05141_);
  or _24366_ (_02428_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nand _24367_ (_02430_, pc_log_change, _02399_);
  and _24368_ (_02432_, _02430_, _05141_);
  and _24369_ (_02797_, _02432_, _02428_);
  or _24370_ (_02433_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  not _24371_ (_02434_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _24372_ (_02435_, pc_log_change, _02434_);
  and _24373_ (_02436_, _02435_, _05141_);
  and _24374_ (_02804_, _02436_, _02433_);
  and _24375_ (_02437_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _24376_ (_02438_, pc_log_change, _02434_);
  or _24377_ (_02439_, _02438_, _02437_);
  and _24378_ (_02806_, _02439_, _05141_);
  and _24379_ (_02440_, _02070_, _06008_);
  nand _24380_ (_02441_, _02440_, _05963_);
  or _24381_ (_02442_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _24382_ (_02443_, _02442_, _05647_);
  and _24383_ (_02444_, _02443_, _02441_);
  nand _24384_ (_02445_, _02078_, _05960_);
  or _24385_ (_02446_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _24386_ (_02447_, _02446_, _05925_);
  and _24387_ (_02448_, _02447_, _02445_);
  and _24388_ (_02449_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _24389_ (_02450_, _02449_, rst);
  or _24390_ (_02451_, _02450_, _02448_);
  or _24391_ (_02824_, _02451_, _02444_);
  or _24392_ (_02452_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand _24393_ (_02453_, _07619_, _06462_);
  and _24394_ (_02454_, _02453_, _05141_);
  and _24395_ (_02828_, _02454_, _02452_);
  nor _24396_ (_02455_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _24397_ (_02830_, _02455_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _24398_ (_02832_, _01280_, _05141_);
  and _24399_ (_02456_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _24400_ (_02457_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  or _24401_ (_02458_, _02457_, _02456_);
  and _24402_ (_02840_, _02458_, _05141_);
  not _24403_ (_02459_, _06678_);
  nor _24404_ (_02460_, _02459_, _05960_);
  and _24405_ (_02461_, _02459_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or _24406_ (_02462_, _02461_, _02460_);
  and _24407_ (_02863_, _02462_, _05141_);
  nor _24408_ (_02463_, _05960_, _08484_);
  and _24409_ (_02464_, _08484_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _24410_ (_02465_, _02464_, _05572_);
  or _24411_ (_02466_, _02465_, _02463_);
  or _24412_ (_02467_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _24413_ (_02468_, _02467_, _05141_);
  and _24414_ (_02871_, _02468_, _02466_);
  nand _24415_ (_02469_, _06707_, _05960_);
  or _24416_ (_02470_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _24417_ (_02471_, _02470_, _05141_);
  and _24418_ (_02876_, _02471_, _02469_);
  or _24419_ (_02472_, _02459_, _05522_);
  or _24420_ (_02473_, _06678_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _24421_ (_02474_, _02473_, _05141_);
  and _24422_ (_02888_, _02474_, _02472_);
  and _24423_ (_02475_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _24424_ (_02476_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or _24425_ (_02897_, _02476_, _02475_);
  and _24426_ (_02477_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _24427_ (_02478_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _24428_ (_02479_, _02478_, _06156_);
  and _24429_ (_02480_, _06180_, _06290_);
  or _24430_ (_02481_, _02480_, _02479_);
  or _24431_ (_02482_, _02481_, _02477_);
  and _24432_ (_02915_, _02482_, _05141_);
  and _24433_ (_02483_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _24434_ (_02484_, _13031_, _05617_);
  or _24435_ (_02485_, _02484_, _02483_);
  and _24436_ (_02925_, _02485_, _05141_);
  nor _24437_ (_02486_, _06180_, _11869_);
  and _24438_ (_02487_, _06180_, _13031_);
  or _24439_ (_02488_, _02487_, _02486_);
  and _24440_ (_02935_, _02488_, _05141_);
  nor _24441_ (_02489_, _08294_, rxd_i);
  and _24442_ (_02490_, _02489_, _06693_);
  nor _24443_ (_02491_, _06693_, _06682_);
  not _24444_ (_02492_, _06684_);
  and _24445_ (_02494_, _08374_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand _24446_ (_02496_, _02494_, _06683_);
  nand _24447_ (_02497_, _02496_, _02492_);
  or _24448_ (_02498_, _02497_, _02491_);
  or _24449_ (_02500_, _02498_, _02490_);
  and _24450_ (_02973_, _02500_, _06715_);
  and _24451_ (_02503_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _24452_ (_02505_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _24453_ (_02987_, _02505_, _02503_);
  and _24454_ (_02999_, _12483_, _05141_);
  and _24455_ (_03006_, _12220_, _05141_);
  and _24456_ (_03011_, _12351_, _05141_);
  or _24457_ (_02506_, _08464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _24458_ (_02507_, _08447_, _08439_);
  or _24459_ (_02508_, _02507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _24460_ (_02509_, _02508_, _11907_);
  or _24461_ (_02510_, _02509_, _08463_);
  and _24462_ (_02511_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _24463_ (_02512_, _02511_, _08457_);
  or _24464_ (_02513_, _02512_, _02510_);
  nand _24465_ (_02514_, _02513_, _02506_);
  nand _24466_ (_02515_, _02514_, _11727_);
  nand _24467_ (_02516_, _08471_, _05560_);
  or _24468_ (_02518_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _24469_ (_02520_, _02518_, _05141_);
  and _24470_ (_02521_, _02520_, _02516_);
  and _24471_ (_03017_, _02521_, _02515_);
  and _24472_ (_03021_, _12588_, _05141_);
  nor _24473_ (_02524_, _11451_, rst);
  and _24474_ (_03031_, _02524_, _12700_);
  and _24475_ (_02527_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _24476_ (_02528_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or _24477_ (_02530_, _02528_, _02527_);
  and _24478_ (_03033_, _02530_, _05141_);
  nor _24479_ (_03035_, _12770_, rst);
  or _24480_ (_02531_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05143_);
  and _24481_ (_02532_, _02531_, _06814_);
  or _24482_ (_02533_, _11443_, _07105_);
  and _24483_ (_02534_, _06995_, _06528_);
  and _24484_ (_02535_, _06995_, _08339_);
  or _24485_ (_02536_, _02535_, _02534_);
  or _24486_ (_02537_, _02536_, _06530_);
  or _24487_ (_02538_, _02537_, _02533_);
  and _24488_ (_02539_, _06778_, _06540_);
  and _24489_ (_02540_, _06771_, _06556_);
  nor _24490_ (_02541_, _02540_, _02539_);
  nand _24491_ (_02542_, _11434_, _02541_);
  or _24492_ (_02543_, _02542_, _02538_);
  or _24493_ (_02544_, _07110_, _06784_);
  or _24494_ (_02545_, _12144_, _11430_);
  and _24495_ (_02546_, _07041_, _06420_);
  or _24496_ (_02547_, _02546_, _01379_);
  or _24497_ (_02548_, _02547_, _02545_);
  or _24498_ (_02549_, _02548_, _02544_);
  or _24499_ (_02550_, _02549_, _02543_);
  and _24500_ (_02551_, _06755_, _06565_);
  or _24501_ (_02552_, _02551_, _06781_);
  and _24502_ (_02553_, _11428_, _06417_);
  or _24503_ (_02554_, _06570_, _06552_);
  and _24504_ (_02555_, _02554_, _06420_);
  or _24505_ (_02556_, _02555_, _02553_);
  or _24506_ (_02557_, _02556_, _02552_);
  or _24507_ (_02558_, _02557_, _01873_);
  or _24508_ (_02559_, _02558_, _02550_);
  and _24509_ (_02560_, _02559_, _06271_);
  or _24510_ (_02561_, _02560_, _02532_);
  and _24511_ (_03039_, _02561_, _05141_);
  and _24512_ (_03045_, _12534_, _05141_);
  nor _24513_ (_02562_, _06244_, _08484_);
  and _24514_ (_02563_, _08484_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _24515_ (_02564_, _02563_, _05572_);
  or _24516_ (_02565_, _02564_, _02562_);
  or _24517_ (_02566_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _24518_ (_02567_, _02566_, _05141_);
  and _24519_ (_03049_, _02567_, _02565_);
  and _24520_ (_02568_, _08280_, _06008_);
  nand _24521_ (_02569_, _02568_, _05963_);
  or _24522_ (_02570_, _02568_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _24523_ (_02571_, _02570_, _08360_);
  and _24524_ (_02572_, _02571_, _02569_);
  nor _24525_ (_02573_, _08360_, _05960_);
  or _24526_ (_02574_, _02573_, _02572_);
  and _24527_ (_03067_, _02574_, _05141_);
  and _24528_ (_02575_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _24529_ (_02576_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _24530_ (_03074_, _02576_, _02575_);
  and _24531_ (_02577_, _06293_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _24532_ (_02578_, _07053_, _06565_);
  and _24533_ (_02579_, _02578_, _06544_);
  or _24534_ (_02580_, _02579_, _02552_);
  and _24535_ (_02581_, _11428_, _06420_);
  and _24536_ (_02582_, _06574_, _06420_);
  and _24537_ (_02583_, _02582_, _06450_);
  or _24538_ (_02584_, _02583_, _02581_);
  or _24539_ (_02585_, _02584_, _02580_);
  or _24540_ (_02586_, _06774_, _06769_);
  or _24541_ (_02587_, _01850_, _12138_);
  or _24542_ (_02588_, _02587_, _02586_);
  or _24543_ (_02589_, _02588_, _02585_);
  or _24544_ (_02590_, _01861_, _06543_);
  or _24545_ (_02591_, _02590_, _02589_);
  and _24546_ (_02592_, _02591_, _06296_);
  or _24547_ (_03080_, _02592_, _02577_);
  and _24548_ (_03087_, _11633_, _06065_);
  and _24549_ (_02593_, _06688_, _01794_);
  and _24550_ (_02594_, _02593_, _06697_);
  or _24551_ (_02595_, _02594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not _24552_ (_02596_, rxd_i);
  nand _24553_ (_02597_, _02594_, _02596_);
  and _24554_ (_02598_, _02597_, _05141_);
  and _24555_ (_03090_, _02598_, _02595_);
  and _24556_ (_02599_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _24557_ (_02600_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _24558_ (_03098_, _02600_, _02599_);
  and _24559_ (_02601_, _02016_, _06008_);
  nand _24560_ (_02602_, _02601_, _05963_);
  or _24561_ (_02603_, _02601_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _24562_ (_02604_, _02603_, _05647_);
  and _24563_ (_02605_, _02604_, _02602_);
  nor _24564_ (_02606_, _02105_, _05960_);
  and _24565_ (_02607_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _24566_ (_02608_, _02607_, _02606_);
  and _24567_ (_02609_, _02608_, _05925_);
  and _24568_ (_02610_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _24569_ (_02611_, _02610_, rst);
  or _24570_ (_02612_, _02611_, _02609_);
  or _24571_ (_03119_, _02612_, _02605_);
  and _24572_ (_02614_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor _24573_ (_02616_, _01802_, _08366_);
  not _24574_ (_02617_, _06693_);
  or _24575_ (_02618_, _02496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _24576_ (_02619_, _02618_, _06686_);
  and _24577_ (_02620_, _02619_, _02617_);
  nor _24578_ (_02621_, _02620_, _01797_);
  nand _24579_ (_02622_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor _24580_ (_02623_, _02622_, _02621_);
  or _24581_ (_02624_, _02623_, _02616_);
  and _24582_ (_02625_, _02624_, _06715_);
  or _24583_ (_03123_, _02625_, _02614_);
  nand _24584_ (_02626_, _08305_, _05960_);
  or _24585_ (_02627_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _24586_ (_02628_, _02627_, _05141_);
  and _24587_ (_03126_, _02628_, _02626_);
  and _24588_ (_02629_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand _24589_ (_02630_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor _24590_ (_02631_, _02630_, _02621_);
  or _24591_ (_02632_, _02631_, _02629_);
  and _24592_ (_02633_, _02632_, _06715_);
  or _24593_ (_03132_, _02633_, _02475_);
  and _24594_ (_02636_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _24595_ (_02637_, _01797_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _24596_ (_02639_, _02637_, _02619_);
  or _24597_ (_02641_, _06693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _24598_ (_02642_, _02641_, _01790_);
  and _24599_ (_02643_, _02642_, _02639_);
  or _24600_ (_02644_, _02643_, _02636_);
  and _24601_ (_02645_, _02644_, _06715_);
  or _24602_ (_03134_, _02645_, _02503_);
  or _24603_ (_02646_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _24604_ (_02647_, _02646_, _02621_);
  or _24605_ (_02648_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _24606_ (_02649_, _02648_, _06715_);
  and _24607_ (_02650_, _02649_, _02647_);
  or _24608_ (_03136_, _02650_, _02575_);
  and _24609_ (_02651_, _01898_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _24610_ (_02652_, _02651_, _01897_);
  and _24611_ (_02653_, _02652_, _10346_);
  or _24612_ (_02654_, _12689_, _05922_);
  nor _24613_ (_02655_, _12690_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _24614_ (_02656_, _02655_, _10346_);
  and _24615_ (_02657_, _02656_, _02654_);
  or _24616_ (_02659_, _02657_, _10354_);
  or _24617_ (_02662_, _02659_, _02653_);
  nand _24618_ (_02663_, _10354_, _05960_);
  and _24619_ (_02665_, _02663_, _05141_);
  and _24620_ (_03139_, _02665_, _02662_);
  or _24621_ (_02667_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _24622_ (_02669_, _02667_, _02621_);
  or _24623_ (_02671_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _24624_ (_02673_, _02671_, _06715_);
  and _24625_ (_02674_, _02673_, _02669_);
  or _24626_ (_03141_, _02674_, _02599_);
  and _24627_ (_02675_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _24628_ (_02676_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _24629_ (_02678_, _02676_, _02621_);
  or _24630_ (_02680_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _24631_ (_02681_, _02680_, _06715_);
  and _24632_ (_02682_, _02681_, _02678_);
  or _24633_ (_03143_, _02682_, _02675_);
  or _24634_ (_02683_, _07080_, _07059_);
  and _24635_ (_02684_, _02683_, _06271_);
  and _24636_ (_02685_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _24637_ (_02686_, _02685_, _07092_);
  or _24638_ (_02687_, _02686_, _02684_);
  and _24639_ (_03150_, _02687_, _05141_);
  and _24640_ (_02688_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _24641_ (_02689_, _07044_, _06450_);
  or _24642_ (_02690_, _02689_, _06979_);
  or _24643_ (_02691_, _02690_, _07072_);
  or _24644_ (_02692_, _02691_, _06820_);
  and _24645_ (_02693_, _02692_, _06271_);
  or _24646_ (_02694_, _02693_, _02688_);
  or _24647_ (_02695_, _02694_, _07090_);
  and _24648_ (_03152_, _02695_, _05141_);
  nand _24649_ (_02696_, _08390_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _24650_ (_02697_, _02696_, _08243_);
  and _24651_ (_02699_, _08243_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _24652_ (_02700_, _02699_, _02697_);
  and _24653_ (_03160_, _02700_, _05141_);
  or _24654_ (_02702_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _24655_ (_02703_, _02702_, _02621_);
  or _24656_ (_02704_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _24657_ (_02706_, _02704_, _06715_);
  and _24658_ (_02707_, _02706_, _02703_);
  or _24659_ (_03168_, _02707_, _06714_);
  or _24660_ (_02708_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _24661_ (_02709_, _02708_, _02621_);
  or _24662_ (_02711_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _24663_ (_02712_, _02711_, _06715_);
  and _24664_ (_02714_, _02712_, _02709_);
  or _24665_ (_03170_, _02714_, _10324_);
  or _24666_ (_02716_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _24667_ (_02717_, _02716_, _02621_);
  and _24668_ (_02718_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _24669_ (_02719_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _24670_ (_02720_, _02719_, _06715_);
  or _24671_ (_02721_, _02720_, _02718_);
  and _24672_ (_03172_, _02721_, _02717_);
  or _24673_ (_02722_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _24674_ (_02724_, _02722_, _02621_);
  and _24675_ (_02725_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _24676_ (_02727_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  and _24677_ (_02728_, _02727_, _06715_);
  or _24678_ (_02729_, _02728_, _02725_);
  and _24679_ (_03175_, _02729_, _02724_);
  or _24680_ (_02731_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _24681_ (_02732_, _02731_, _02621_);
  and _24682_ (_02733_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _24683_ (_02735_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  and _24684_ (_02736_, _02735_, _06715_);
  or _24685_ (_02737_, _02736_, _02733_);
  and _24686_ (_03178_, _02737_, _02732_);
  nor _24687_ (_02739_, _10407_, _05751_);
  or _24688_ (_02740_, _02739_, _11665_);
  nand _24689_ (_02741_, _02740_, _08163_);
  nor _24690_ (_02742_, _07200_, _06842_);
  and _24691_ (_02743_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _24692_ (_02744_, _02743_, _02742_);
  nand _24693_ (_02745_, _02744_, _02741_);
  nand _24694_ (_02746_, _02745_, _08158_);
  nand _24695_ (_02747_, _07166_, _06836_);
  nand _24696_ (_02748_, _02747_, _02746_);
  and _24697_ (_03180_, _02748_, _05141_);
  and _24698_ (_03183_, _12444_, _05141_);
  nor _24699_ (_02749_, _06620_, _05464_);
  or _24700_ (_02750_, _02749_, _10356_);
  nand _24701_ (_02751_, _02750_, _08163_);
  nor _24702_ (_02752_, _06842_, _06617_);
  and _24703_ (_02753_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _24704_ (_02754_, _02753_, _02752_);
  and _24705_ (_02755_, _02754_, _08158_);
  nand _24706_ (_02756_, _02755_, _02751_);
  or _24707_ (_02757_, _07378_, _08158_);
  and _24708_ (_02758_, _02757_, _02756_);
  and _24709_ (_03193_, _02758_, _05141_);
  or _24710_ (_02761_, _11443_, _07070_);
  and _24711_ (_02762_, _06755_, _06557_);
  or _24712_ (_02763_, _02762_, _02582_);
  or _24713_ (_02764_, _02763_, _02761_);
  or _24714_ (_02765_, _07062_, _06818_);
  or _24715_ (_02766_, _08334_, _02765_);
  or _24716_ (_02767_, _02766_, _02764_);
  or _24717_ (_02769_, _11429_, _02539_);
  or _24718_ (_02770_, _02769_, _06819_);
  or _24719_ (_02772_, _02770_, _02767_);
  or _24720_ (_02773_, _12671_, _06530_);
  and _24721_ (_02774_, _06828_, _06420_);
  or _24722_ (_02775_, _02774_, _06795_);
  or _24723_ (_02776_, _02775_, _02555_);
  or _24724_ (_02777_, _02776_, _02773_);
  and _24725_ (_02778_, _06755_, _06765_);
  and _24726_ (_02779_, _06547_, _06420_);
  or _24727_ (_02781_, _02779_, _02778_);
  or _24728_ (_02782_, _02781_, _01864_);
  and _24729_ (_02783_, _06828_, _06760_);
  and _24730_ (_02784_, _06564_, _06544_);
  or _24731_ (_02785_, _02784_, _02783_);
  or _24732_ (_02786_, _02785_, _02782_);
  or _24733_ (_02787_, _02786_, _02777_);
  or _24734_ (_02788_, _02553_, _01870_);
  and _24735_ (_02789_, _06755_, _06566_);
  or _24736_ (_02790_, _01379_, _06793_);
  or _24737_ (_02791_, _02790_, _02789_);
  or _24738_ (_02792_, _02791_, _06541_);
  or _24739_ (_02793_, _02792_, _02788_);
  or _24740_ (_02794_, _02793_, _02787_);
  or _24741_ (_02795_, _02794_, _02772_);
  and _24742_ (_02796_, _02795_, _06271_);
  and _24743_ (_02798_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _24744_ (_02799_, _06796_, _06821_);
  or _24745_ (_02800_, _02799_, _06813_);
  or _24746_ (_02801_, _02800_, _02798_);
  or _24747_ (_02802_, _02801_, _02796_);
  and _24748_ (_03195_, _02802_, _05141_);
  or _24749_ (_02803_, _01851_, _07037_);
  and _24750_ (_02805_, _02803_, _06531_);
  or _24751_ (_02807_, _02769_, _08332_);
  or _24752_ (_02808_, _02807_, _02805_);
  or _24753_ (_02809_, _12139_, _08334_);
  or _24754_ (_02810_, _02809_, _02781_);
  and _24755_ (_02811_, _07069_, _06528_);
  or _24756_ (_02812_, _11443_, _07042_);
  or _24757_ (_02813_, _02812_, _02811_);
  and _24758_ (_02814_, _06778_, _06528_);
  or _24759_ (_02815_, _02814_, _06781_);
  or _24760_ (_02816_, _07073_, _06793_);
  or _24761_ (_02817_, _02816_, _02815_);
  or _24762_ (_02818_, _02817_, _02813_);
  or _24763_ (_02819_, _02818_, _02810_);
  or _24764_ (_02820_, _02788_, _02777_);
  or _24765_ (_02821_, _02820_, _02819_);
  or _24766_ (_02822_, _02821_, _02808_);
  and _24767_ (_02823_, _02822_, _06271_);
  and _24768_ (_02825_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _24769_ (_02826_, _02825_, _02800_);
  or _24770_ (_02827_, _02826_, _02823_);
  and _24771_ (_03198_, _02827_, _05141_);
  and _24772_ (_02829_, _06154_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _24773_ (_02831_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _24774_ (_02833_, _02831_, _06156_);
  and _24775_ (_02834_, _05605_, _05291_);
  or _24776_ (_02835_, _02834_, _02833_);
  or _24777_ (_02836_, _02835_, _02829_);
  and _24778_ (_03300_, _02836_, _05141_);
  nor _24779_ (_02837_, _07259_, _06842_);
  and _24780_ (_02838_, _08171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _24781_ (_02839_, _02838_, _02837_);
  nor _24782_ (_02841_, _02839_, _06836_);
  not _24783_ (_02842_, _02841_);
  not _24784_ (_02843_, _08163_);
  nor _24785_ (_02844_, _08469_, _05339_);
  nor _24786_ (_02845_, _02844_, _10380_);
  or _24787_ (_02846_, _02845_, _02843_);
  nand _24788_ (_02847_, _07229_, _06836_);
  and _24789_ (_02848_, _02847_, _02846_);
  and _24790_ (_02849_, _02848_, _02842_);
  nor _24791_ (_03305_, _02849_, rst);
  and _24792_ (_02850_, _06293_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _24793_ (_02851_, _06570_, _06566_);
  or _24794_ (_02852_, _06767_, _06553_);
  or _24795_ (_02853_, _02852_, _02851_);
  and _24796_ (_02854_, _02853_, _06536_);
  or _24797_ (_02855_, _02854_, _00612_);
  or _24798_ (_02856_, _02789_, _11443_);
  or _24799_ (_02857_, _02856_, _06989_);
  or _24800_ (_02858_, _02857_, _07048_);
  or _24801_ (_02859_, _02858_, _02544_);
  nand _24802_ (_02860_, _06773_, _06566_);
  nand _24803_ (_02861_, _02860_, _07051_);
  and _24804_ (_02862_, _06570_, _06420_);
  or _24805_ (_02864_, _02862_, _06756_);
  or _24806_ (_02865_, _02539_, _06997_);
  or _24807_ (_02866_, _02865_, _02864_);
  or _24808_ (_02867_, _02866_, _02861_);
  or _24809_ (_02868_, _02867_, _06985_);
  or _24810_ (_02869_, _02868_, _02859_);
  or _24811_ (_02870_, _02869_, _02855_);
  and _24812_ (_02872_, _02870_, _06296_);
  or _24813_ (_03316_, _02872_, _02850_);
  and _24814_ (_02873_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _24815_ (_02874_, pc_log_change, _08551_);
  or _24816_ (_02875_, _02874_, _02873_);
  and _24817_ (_03319_, _02875_, _05141_);
  and _24818_ (_02877_, _06283_, _05617_);
  and _24819_ (_02878_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _24820_ (_02879_, _02878_, _02877_);
  and _24821_ (_03372_, _02879_, _05141_);
  nand _24822_ (_02880_, _08265_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or _24823_ (_02881_, _08265_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _24824_ (_02882_, _02881_, _05141_);
  nand _24825_ (_02883_, _02882_, _02880_);
  nor _24826_ (_03519_, _02883_, _08243_);
  and _24827_ (_02884_, _09451_, _08385_);
  and _24828_ (_02885_, _08388_, _09438_);
  and _24829_ (_02886_, _02885_, _09451_);
  nor _24830_ (_02887_, _08388_, _00625_);
  or _24831_ (_02889_, _02887_, _02886_);
  and _24832_ (_02890_, _02889_, _08246_);
  nand _24833_ (_02891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _24834_ (_02892_, _02891_, _08245_);
  or _24835_ (_02893_, _02892_, _02890_);
  and _24836_ (_02894_, _02893_, _09437_);
  or _24837_ (_02895_, _02894_, _02884_);
  nand _24838_ (_02896_, _02895_, _05141_);
  nor _24839_ (_03523_, _02896_, _08243_);
  or _24840_ (_02898_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand _24841_ (_02899_, pc_log_change, _02425_);
  and _24842_ (_02900_, _02899_, _05141_);
  and _24843_ (_03601_, _02900_, _02898_);
  and _24844_ (_02901_, _05615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _24845_ (_02902_, _05617_, _05561_);
  or _24846_ (_02903_, _02902_, _02901_);
  and _24847_ (_03623_, _02903_, _05141_);
  or _24848_ (_02904_, _12117_, _06996_);
  or _24849_ (_02905_, _02904_, _11429_);
  or _24850_ (_02906_, _02905_, _02553_);
  or _24851_ (_02907_, _02906_, _01866_);
  or _24852_ (_02908_, _02907_, _02792_);
  or _24853_ (_02909_, _01870_, _06979_);
  and _24854_ (_02910_, _02909_, _06449_);
  or _24855_ (_02911_, _02762_, _13288_);
  or _24856_ (_02912_, _02911_, _02862_);
  or _24857_ (_02913_, _02912_, _08336_);
  or _24858_ (_02914_, _01859_, _12131_);
  or _24859_ (_02916_, _02914_, _02913_);
  or _24860_ (_02917_, _02916_, _02910_);
  or _24861_ (_02918_, _02917_, _02908_);
  and _24862_ (_02919_, _02918_, _06296_);
  nor _24863_ (_02920_, _06821_, rst);
  and _24864_ (_02921_, _02920_, _06793_);
  and _24865_ (_02922_, _06293_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or _24866_ (_02923_, _02922_, _02921_);
  or _24867_ (_03634_, _02923_, _02919_);
  nor _24868_ (_02924_, _02773_, _01867_);
  nand _24869_ (_02926_, _02924_, _11445_);
  or _24870_ (_02927_, _06994_, _12927_);
  or _24871_ (_02928_, _02927_, _12112_);
  or _24872_ (_02929_, _02928_, _01381_);
  or _24873_ (_02930_, _02929_, _02926_);
  and _24874_ (_02931_, _06767_, _06535_);
  or _24875_ (_02932_, _02931_, _02774_);
  or _24876_ (_02933_, _02932_, _06780_);
  and _24877_ (_02934_, _06773_, _06564_);
  or _24878_ (_02936_, _02865_, _02781_);
  or _24879_ (_02937_, _02936_, _02934_);
  or _24880_ (_02938_, _02937_, _06764_);
  or _24881_ (_02939_, _02938_, _02933_);
  or _24882_ (_02940_, _02939_, _02930_);
  and _24883_ (_02941_, _02940_, _06271_);
  and _24884_ (_02942_, _06793_, _05143_);
  and _24885_ (_02943_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _24886_ (_02944_, _02943_, _02942_);
  or _24887_ (_02945_, _02944_, _02941_);
  and _24888_ (_03637_, _02945_, _05141_);
  and _24889_ (_02946_, _12261_, _12372_);
  and _24890_ (_02947_, _02946_, _01362_);
  and _24891_ (_02948_, _02947_, _06838_);
  nor _24892_ (_02949_, _02948_, _12697_);
  and _24893_ (_02950_, _01288_, _06703_);
  or _24894_ (_02951_, _02950_, _12610_);
  and _24895_ (_02952_, _01303_, _06179_);
  and _24896_ (_02953_, _01279_, _05561_);
  and _24897_ (_02954_, _01309_, _06290_);
  or _24898_ (_02955_, _02954_, _02953_);
  or _24899_ (_02956_, _02955_, _02952_);
  or _24900_ (_02957_, _02956_, _02951_);
  and _24901_ (_02958_, _01288_, _05522_);
  or _24902_ (_02959_, _02958_, _12608_);
  and _24903_ (_02960_, _01309_, _13031_);
  and _24904_ (_02961_, _01279_, _06283_);
  and _24905_ (_02962_, _01303_, _06004_);
  or _24906_ (_02963_, _02962_, _02961_);
  or _24907_ (_02964_, _02963_, _02960_);
  or _24908_ (_02965_, _02964_, _02959_);
  nand _24909_ (_02966_, _02965_, _02957_);
  nor _24910_ (_02967_, _02966_, _02949_);
  and _24911_ (_02968_, _12372_, _01280_);
  nand _24912_ (_02969_, _02968_, _12263_);
  or _24913_ (_02970_, _02969_, _01419_);
  nand _24914_ (_02971_, _02757_, _02756_);
  nand _24915_ (_02972_, _02971_, _08415_);
  or _24916_ (_02974_, _02971_, _08415_);
  nand _24917_ (_02975_, _02974_, _02972_);
  nand _24918_ (_02976_, _08187_, _08186_);
  nand _24919_ (_02977_, _08509_, _02976_);
  or _24920_ (_02978_, _08509_, _02976_);
  and _24921_ (_02979_, _02978_, _02977_);
  nand _24922_ (_02980_, _02979_, _02975_);
  or _24923_ (_02981_, _02979_, _02975_);
  nand _24924_ (_02982_, _02981_, _02980_);
  nand _24925_ (_02983_, _02748_, _08177_);
  or _24926_ (_02984_, _02748_, _08177_);
  and _24927_ (_02985_, _02984_, _02983_);
  nand _24928_ (_02986_, _02985_, _02982_);
  or _24929_ (_02988_, _02985_, _02982_);
  and _24930_ (_02989_, _02988_, _02986_);
  nand _24931_ (_02990_, _02849_, _06977_);
  or _24932_ (_02991_, _02849_, _06977_);
  and _24933_ (_02992_, _02991_, _02990_);
  nand _24934_ (_02993_, _02992_, _02989_);
  or _24935_ (_02994_, _02992_, _02989_);
  and _24936_ (_02995_, _02994_, _02993_);
  nand _24937_ (_02996_, _02995_, _12608_);
  or _24938_ (_02997_, _12608_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _24939_ (_02998_, _02997_, _01288_);
  and _24940_ (_03000_, _02998_, _02996_);
  and _24941_ (_03001_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _24942_ (_03002_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _24943_ (_03003_, _03002_, _03001_);
  and _24944_ (_03004_, _03003_, _12610_);
  and _24945_ (_03005_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _24946_ (_03007_, _12608_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _24947_ (_03008_, _03007_, _03005_);
  and _24948_ (_03009_, _03008_, _01279_);
  and _24949_ (_03010_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _24950_ (_03012_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _24951_ (_03013_, _03012_, _03010_);
  and _24952_ (_03014_, _03013_, _12608_);
  or _24953_ (_03015_, _03014_, _03009_);
  or _24954_ (_03016_, _03015_, _03004_);
  nor _24955_ (_03018_, _03016_, _03000_);
  nor _24956_ (_03019_, _03018_, _02970_);
  and _24957_ (_03020_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _24958_ (_03022_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _24959_ (_03023_, _03022_, _03020_);
  and _24960_ (_03024_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _24961_ (_03025_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _24962_ (_03026_, _03025_, _03024_);
  or _24963_ (_03027_, _03026_, _03023_);
  and _24964_ (_03028_, _03027_, _12608_);
  and _24965_ (_03029_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _24966_ (_03030_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _24967_ (_03032_, _03030_, _03029_);
  and _24968_ (_03034_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _24969_ (_03036_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _24970_ (_03038_, _03036_, _03034_);
  or _24971_ (_03040_, _03038_, _03032_);
  and _24972_ (_03041_, _03040_, _12610_);
  nor _24973_ (_03042_, _03041_, _03028_);
  nor _24974_ (_03043_, _03042_, _01318_);
  and _24975_ (_03044_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _24976_ (_03046_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _24977_ (_03047_, _03046_, _03044_);
  and _24978_ (_03048_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _24979_ (_03050_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _24980_ (_03051_, _03050_, _03048_);
  or _24981_ (_03052_, _03051_, _03047_);
  and _24982_ (_03053_, _03052_, _12608_);
  and _24983_ (_03054_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _24984_ (_03055_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _24985_ (_03056_, _03055_, _03054_);
  and _24986_ (_03057_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _24987_ (_03058_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _24988_ (_03059_, _03058_, _03057_);
  or _24989_ (_03060_, _03059_, _03056_);
  and _24990_ (_03061_, _03060_, _12610_);
  or _24991_ (_03062_, _03061_, _03053_);
  and _24992_ (_03063_, _03062_, _01283_);
  and _24993_ (_03064_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _24994_ (_03065_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _24995_ (_03066_, _03065_, _03064_);
  and _24996_ (_03068_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _24997_ (_03069_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _24998_ (_03070_, _03069_, _03068_);
  or _24999_ (_03071_, _03070_, _03066_);
  and _25000_ (_03072_, _03071_, _12608_);
  and _25001_ (_03073_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _25002_ (_03075_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _25003_ (_03076_, _03075_, _03073_);
  and _25004_ (_03077_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _25005_ (_03078_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _25006_ (_03079_, _03078_, _03077_);
  or _25007_ (_03081_, _03079_, _03076_);
  and _25008_ (_03082_, _03081_, _12610_);
  or _25009_ (_03083_, _03082_, _03072_);
  and _25010_ (_03084_, _03083_, _01343_);
  or _25011_ (_03085_, _03084_, _03063_);
  or _25012_ (_03086_, _03085_, _03043_);
  and _25013_ (_03088_, _03086_, _12374_);
  or _25014_ (_03089_, _01391_, p3_in[6]);
  or _25015_ (_03091_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _25016_ (_03092_, _03091_, _03089_);
  and _25017_ (_03093_, _03092_, _01279_);
  or _25018_ (_03094_, _03093_, _12608_);
  and _25019_ (_03095_, _01402_, _01309_);
  or _25020_ (_03096_, _01391_, p3_in[4]);
  or _25021_ (_03097_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _25022_ (_03099_, _03097_, _03096_);
  and _25023_ (_03100_, _03099_, _01288_);
  or _25024_ (_03101_, _01391_, p3_in[5]);
  or _25025_ (_03102_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _25026_ (_03103_, _03102_, _03101_);
  and _25027_ (_03104_, _03103_, _01303_);
  or _25028_ (_03105_, _03104_, _03100_);
  or _25029_ (_03106_, _03105_, _03095_);
  or _25030_ (_03107_, _03106_, _03094_);
  nor _25031_ (_03108_, _01391_, p3_in[0]);
  and _25032_ (_03109_, _01391_, _02024_);
  nor _25033_ (_03110_, _03109_, _03108_);
  and _25034_ (_03111_, _03110_, _01288_);
  or _25035_ (_03112_, _03111_, _12610_);
  or _25036_ (_03113_, _01391_, p3_in[3]);
  or _25037_ (_03114_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _25038_ (_03115_, _03114_, _03113_);
  and _25039_ (_03116_, _03115_, _01309_);
  or _25040_ (_03117_, _01391_, p3_in[2]);
  or _25041_ (_03118_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _25042_ (_03120_, _03118_, _03117_);
  and _25043_ (_03121_, _03120_, _01279_);
  or _25044_ (_03122_, _01391_, p3_in[1]);
  or _25045_ (_03124_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _25046_ (_03125_, _03124_, _03122_);
  and _25047_ (_03127_, _03125_, _01303_);
  or _25048_ (_03128_, _03127_, _03121_);
  or _25049_ (_03129_, _03128_, _03116_);
  or _25050_ (_03130_, _03129_, _03112_);
  and _25051_ (_03131_, _03130_, _03107_);
  or _25052_ (_03133_, _03131_, _12261_);
  or _25053_ (_03135_, _01317_, _12374_);
  or _25054_ (_03137_, _01391_, p2_in[4]);
  or _25055_ (_03138_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _25056_ (_03140_, _03138_, _03137_);
  and _25057_ (_03142_, _03140_, _01288_);
  or _25058_ (_03144_, _03142_, _12608_);
  or _25059_ (_03145_, _01391_, p2_in[6]);
  or _25060_ (_03146_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _25061_ (_03147_, _03146_, _03145_);
  and _25062_ (_03148_, _03147_, _01279_);
  or _25063_ (_03149_, _01391_, p2_in[5]);
  or _25064_ (_03151_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _25065_ (_03153_, _03151_, _03149_);
  and _25066_ (_03154_, _03153_, _01303_);
  and _25067_ (_03155_, _01397_, _01309_);
  or _25068_ (_03156_, _03155_, _03154_);
  or _25069_ (_03157_, _03156_, _03148_);
  or _25070_ (_03158_, _03157_, _03144_);
  or _25071_ (_03159_, _01391_, p2_in[1]);
  or _25072_ (_03161_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _25073_ (_03162_, _03161_, _03159_);
  and _25074_ (_03163_, _03162_, _01303_);
  or _25075_ (_03164_, _03163_, _12610_);
  or _25076_ (_03165_, _01391_, p2_in[2]);
  or _25077_ (_03166_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _25078_ (_03167_, _03166_, _03165_);
  and _25079_ (_03169_, _03167_, _01279_);
  nor _25080_ (_03171_, _01391_, p2_in[0]);
  and _25081_ (_03173_, _01391_, _02062_);
  nor _25082_ (_03174_, _03173_, _03171_);
  and _25083_ (_03176_, _03174_, _01288_);
  or _25084_ (_03177_, _01391_, p2_in[3]);
  or _25085_ (_03179_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _25086_ (_03181_, _03179_, _03177_);
  and _25087_ (_03182_, _03181_, _01309_);
  or _25088_ (_03184_, _03182_, _03176_);
  or _25089_ (_03185_, _03184_, _03169_);
  or _25090_ (_03186_, _03185_, _03164_);
  and _25091_ (_03187_, _03186_, _03158_);
  nor _25092_ (_03188_, _03187_, _12263_);
  nor _25093_ (_03189_, _03188_, _03135_);
  and _25094_ (_03190_, _03189_, _03133_);
  or _25095_ (_03191_, _01391_, p1_in[3]);
  or _25096_ (_03192_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25097_ (_03194_, _03192_, _03191_);
  and _25098_ (_03196_, _03194_, _01309_);
  or _25099_ (_03197_, _03196_, _12610_);
  or _25100_ (_03199_, _01391_, p1_in[1]);
  or _25101_ (_03200_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25102_ (_03201_, _03200_, _03199_);
  and _25103_ (_03202_, _03201_, _01303_);
  or _25104_ (_03203_, _01391_, p1_in[2]);
  or _25105_ (_03204_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _25106_ (_03205_, _03204_, _03203_);
  and _25107_ (_03206_, _03205_, _01279_);
  nor _25108_ (_03207_, _01391_, p1_in[0]);
  and _25109_ (_03208_, _01391_, _02233_);
  nor _25110_ (_03209_, _03208_, _03207_);
  and _25111_ (_03210_, _03209_, _01288_);
  or _25112_ (_03211_, _03210_, _03206_);
  or _25113_ (_03212_, _03211_, _03202_);
  or _25114_ (_03213_, _03212_, _03197_);
  and _25115_ (_03214_, _01343_, _12372_);
  and _25116_ (_03215_, _01412_, _01309_);
  or _25117_ (_03216_, _03215_, _12608_);
  or _25118_ (_03217_, _01391_, p1_in[5]);
  or _25119_ (_03218_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25120_ (_03219_, _03218_, _03217_);
  and _25121_ (_03220_, _03219_, _01303_);
  or _25122_ (_03221_, _01391_, p1_in[6]);
  or _25123_ (_03222_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _25124_ (_03223_, _03222_, _03221_);
  and _25125_ (_03224_, _03223_, _01279_);
  or _25126_ (_03225_, _01391_, p1_in[4]);
  or _25127_ (_03226_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _25128_ (_03227_, _03226_, _03225_);
  and _25129_ (_03228_, _03227_, _01288_);
  or _25130_ (_03229_, _03228_, _03224_);
  or _25131_ (_03230_, _03229_, _03220_);
  or _25132_ (_03231_, _03230_, _03216_);
  and _25133_ (_03232_, _03231_, _03214_);
  and _25134_ (_03233_, _03232_, _03213_);
  and _25135_ (_03234_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _25136_ (_03235_, _03234_, _12608_);
  and _25137_ (_03236_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _25138_ (_03237_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _25139_ (_03238_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _25140_ (_03239_, _03238_, _03237_);
  or _25141_ (_03240_, _03239_, _03236_);
  or _25142_ (_03241_, _03240_, _03235_);
  and _25143_ (_03242_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _25144_ (_03243_, _03242_, _12610_);
  and _25145_ (_03244_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _25146_ (_03245_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _25147_ (_03246_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _25148_ (_03247_, _03246_, _03245_);
  or _25149_ (_03248_, _03247_, _03244_);
  or _25150_ (_03249_, _03248_, _03243_);
  and _25151_ (_03250_, _03249_, _02947_);
  and _25152_ (_03251_, _03250_, _03241_);
  or _25153_ (_03252_, _03251_, _03233_);
  and _25154_ (_03253_, _12261_, _12374_);
  nand _25155_ (_03254_, _03253_, _01280_);
  or _25156_ (_03255_, _03254_, _01419_);
  and _25157_ (_03256_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _25158_ (_03257_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _25159_ (_03258_, _03257_, _03256_);
  and _25160_ (_03259_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _25161_ (_03260_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _25162_ (_03261_, _03260_, _03259_);
  or _25163_ (_03262_, _03261_, _03258_);
  and _25164_ (_03263_, _03262_, _12608_);
  and _25165_ (_03264_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25166_ (_03265_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _25167_ (_03266_, _03265_, _03264_);
  and _25168_ (_03267_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _25169_ (_03268_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _25170_ (_03269_, _03268_, _03267_);
  or _25171_ (_03270_, _03269_, _03266_);
  and _25172_ (_03271_, _03270_, _12610_);
  nor _25173_ (_03272_, _03271_, _03263_);
  nor _25174_ (_03273_, _03272_, _03255_);
  and _25175_ (_03274_, _01322_, _12374_);
  and _25176_ (_03275_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _25177_ (_03276_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _25178_ (_03277_, _03276_, _03275_);
  and _25179_ (_03278_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _25180_ (_03279_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _25181_ (_03280_, _03279_, _03278_);
  or _25182_ (_03281_, _03280_, _03277_);
  and _25183_ (_03282_, _03281_, _12608_);
  and _25184_ (_03283_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _25185_ (_03284_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _25186_ (_03285_, _03284_, _03283_);
  and _25187_ (_03286_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _25188_ (_03287_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _25189_ (_03288_, _03287_, _03286_);
  or _25190_ (_03289_, _03288_, _03285_);
  and _25191_ (_03290_, _03289_, _12610_);
  or _25192_ (_03291_, _03290_, _03282_);
  and _25193_ (_03292_, _03291_, _03274_);
  or _25194_ (_03293_, _03292_, _03273_);
  or _25195_ (_03294_, _03293_, _03252_);
  and _25196_ (_03295_, _12615_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  nand _25197_ (_03296_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _25198_ (_03297_, _03296_, _12610_);
  not _25199_ (_03298_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _25200_ (_03299_, _12557_, _12502_);
  or _25201_ (_03301_, _03299_, _03298_);
  nand _25202_ (_03302_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _25203_ (_03303_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _25204_ (_03304_, _03303_, _03302_);
  and _25205_ (_03306_, _03304_, _03301_);
  and _25206_ (_03307_, _03306_, _03297_);
  and _25207_ (_03308_, _12448_, _12313_);
  not _25208_ (_03309_, _03308_);
  or _25209_ (_03310_, _02969_, _03309_);
  nand _25210_ (_03311_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _25211_ (_03312_, _03311_, _12608_);
  nand _25212_ (_03313_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _25213_ (_03314_, _01303_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _25214_ (_03315_, _03299_, _00747_);
  and _25215_ (_03317_, _03315_, _03314_);
  and _25216_ (_03318_, _03317_, _03313_);
  and _25217_ (_03320_, _03318_, _03312_);
  or _25218_ (_03321_, _03320_, _03310_);
  nor _25219_ (_03322_, _03321_, _03307_);
  or _25220_ (_03323_, _03322_, _03295_);
  or _25221_ (_03324_, _01342_, _12374_);
  and _25222_ (_03325_, _03310_, _03135_);
  and _25223_ (_03326_, _03325_, _03324_);
  not _25224_ (_03327_, _02970_);
  nor _25225_ (_03328_, _03327_, _02947_);
  nand _25226_ (_03329_, _01281_, _12374_);
  and _25227_ (_03330_, _03329_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _25228_ (_03331_, _03330_, _03255_);
  and _25229_ (_03332_, _03331_, _03328_);
  and _25230_ (_03333_, _03332_, _03326_);
  or _25231_ (_03334_, _01391_, p0_in[4]);
  or _25232_ (_03335_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25233_ (_03336_, _03335_, _03334_);
  and _25234_ (_03337_, _03336_, _01288_);
  or _25235_ (_03338_, _03337_, _12608_);
  or _25236_ (_03339_, _01391_, p0_in[5]);
  or _25237_ (_03340_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25238_ (_03341_, _03340_, _03339_);
  and _25239_ (_03342_, _03341_, _01303_);
  and _25240_ (_03343_, _01408_, _01309_);
  or _25241_ (_03344_, _01391_, p0_in[6]);
  or _25242_ (_03345_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25243_ (_03346_, _03345_, _03344_);
  and _25244_ (_03347_, _03346_, _01279_);
  or _25245_ (_03348_, _03347_, _03343_);
  or _25246_ (_03349_, _03348_, _03342_);
  or _25247_ (_03350_, _03349_, _03338_);
  and _25248_ (_03351_, _01283_, _12372_);
  nor _25249_ (_03352_, _01391_, p0_in[0]);
  and _25250_ (_03353_, _01391_, _02094_);
  nor _25251_ (_03354_, _03353_, _03352_);
  and _25252_ (_03355_, _03354_, _01288_);
  or _25253_ (_03356_, _03355_, _12610_);
  or _25254_ (_03357_, _01391_, p0_in[2]);
  or _25255_ (_03358_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25256_ (_03359_, _03358_, _03357_);
  and _25257_ (_03360_, _03359_, _01279_);
  or _25258_ (_03361_, _01391_, p0_in[3]);
  or _25259_ (_03362_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _25260_ (_03363_, _03362_, _03361_);
  and _25261_ (_03364_, _03363_, _01309_);
  or _25262_ (_03365_, _01391_, p0_in[1]);
  or _25263_ (_03366_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _25264_ (_03367_, _03366_, _03365_);
  and _25265_ (_03368_, _03367_, _01303_);
  or _25266_ (_03369_, _03368_, _03364_);
  or _25267_ (_03370_, _03369_, _03360_);
  or _25268_ (_03371_, _03370_, _03356_);
  and _25269_ (_03373_, _03371_, _03351_);
  and _25270_ (_03374_, _03373_, _03350_);
  or _25271_ (_03375_, _03374_, _03333_);
  or _25272_ (_03376_, _03375_, _03323_);
  or _25273_ (_03377_, _03376_, _03294_);
  or _25274_ (_03378_, _03377_, _03190_);
  or _25275_ (_03379_, _03378_, _03088_);
  or _25276_ (_03380_, _03379_, _03019_);
  nand _25277_ (_03381_, _03295_, _05963_);
  and _25278_ (_03382_, _03381_, _02949_);
  and _25279_ (_03383_, _03382_, _03380_);
  or _25280_ (_03384_, _03383_, _02967_);
  and _25281_ (_03643_, _03384_, _05141_);
  nand _25282_ (_03385_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _25283_ (_03386_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _25284_ (_03387_, _03386_, _03385_);
  nand _25285_ (_03388_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _25286_ (_03389_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _25287_ (_03390_, _03389_, _03388_);
  and _25288_ (_03391_, _03390_, _03387_);
  nand _25289_ (_03392_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _25290_ (_03393_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _25291_ (_03394_, _03393_, _03392_);
  nand _25292_ (_03395_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _25293_ (_03396_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _25294_ (_03397_, _03396_, _03395_);
  and _25295_ (_03398_, _03397_, _03394_);
  and _25296_ (_03399_, _03398_, _03391_);
  nand _25297_ (_03400_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand _25298_ (_03401_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _25299_ (_03402_, _03401_, _03400_);
  nand _25300_ (_03403_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _25301_ (_03404_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _25302_ (_03405_, _03404_, _03403_);
  and _25303_ (_03406_, _03405_, _03402_);
  nand _25304_ (_03407_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _25305_ (_03408_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _25306_ (_03409_, _03408_, _03407_);
  nand _25307_ (_03410_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _25308_ (_03411_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and _25309_ (_03412_, _03411_, _03410_);
  and _25310_ (_03413_, _03412_, _03409_);
  and _25311_ (_03414_, _03413_, _03406_);
  and _25312_ (_03415_, _03414_, _03399_);
  nand _25313_ (_03416_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _25314_ (_03417_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _25315_ (_03418_, _03417_, _03416_);
  nand _25316_ (_03419_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not _25317_ (_03420_, _12463_);
  nand _25318_ (_03421_, _01368_, _03420_);
  and _25319_ (_03422_, _03421_, _03419_);
  and _25320_ (_03423_, _03422_, _03418_);
  nand _25321_ (_03424_, _03110_, _01399_);
  nand _25322_ (_03425_, _03174_, _01373_);
  and _25323_ (_03426_, _03425_, _03424_);
  nand _25324_ (_03427_, _03354_, _01405_);
  nand _25325_ (_03428_, _03209_, _01413_);
  and _25326_ (_03429_, _03428_, _03427_);
  and _25327_ (_03430_, _03429_, _03426_);
  and _25328_ (_03431_, _03430_, _03423_);
  not _25329_ (_03432_, _01422_);
  or _25330_ (_03433_, _02995_, _03432_);
  nand _25331_ (_03434_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _25332_ (_03435_, _03434_, _03433_);
  and _25333_ (_03436_, _03435_, _03431_);
  and _25334_ (_03437_, _03436_, _03415_);
  nor _25335_ (_03438_, _03437_, _01443_);
  not _25336_ (_03439_, _01287_);
  nand _25337_ (_03440_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _25338_ (_03441_, _03440_, _03439_);
  or _25339_ (_03442_, _03441_, _03438_);
  nand _25340_ (_03443_, _01287_, _07496_);
  and _25341_ (_03444_, _03443_, _05141_);
  and _25342_ (_03688_, _03444_, _03442_);
  or _25343_ (_03445_, _06979_, _06772_);
  or _25344_ (_03446_, _03445_, _06998_);
  or _25345_ (_03447_, _03446_, _06763_);
  or _25346_ (_03448_, _03447_, _00611_);
  or _25347_ (_03449_, _01869_, _01380_);
  or _25348_ (_03450_, _02934_, _02864_);
  or _25349_ (_03451_, _03450_, _03449_);
  or _25350_ (_03452_, _03451_, _02933_);
  or _25351_ (_03453_, _03452_, _03448_);
  and _25352_ (_03454_, _03453_, _06271_);
  and _25353_ (_03455_, _06795_, _05143_);
  and _25354_ (_03456_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25355_ (_03457_, _03456_, _03455_);
  or _25356_ (_03458_, _03457_, _03454_);
  and _25357_ (_03698_, _03458_, _05141_);
  or _25358_ (_03459_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _25359_ (_03460_, _01048_, rst);
  and _25360_ (_03700_, _03460_, _03459_);
  or _25361_ (_03461_, _01287_, rst);
  nor _25362_ (_03709_, _03461_, _01441_);
  nand _25363_ (_03462_, _02886_, _08245_);
  nand _25364_ (_03463_, _03462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _25365_ (_03464_, _03463_, _02884_);
  or _25366_ (_03465_, _03464_, _08243_);
  and _25367_ (_03713_, _03465_, _05141_);
  and _25368_ (_03466_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _25369_ (_03467_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _25370_ (_03468_, _03467_, _03466_);
  and _25371_ (_03469_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _25372_ (_03470_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _25373_ (_03471_, _03470_, _03469_);
  or _25374_ (_03472_, _03471_, _03468_);
  and _25375_ (_03473_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _25376_ (_03474_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _25377_ (_03475_, _03474_, _03473_);
  and _25378_ (_03476_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _25379_ (_03477_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _25380_ (_03478_, _03477_, _03476_);
  or _25381_ (_03479_, _03478_, _03475_);
  or _25382_ (_03480_, _03479_, _03472_);
  and _25383_ (_03481_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _25384_ (_03482_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _25385_ (_03483_, _03482_, _03481_);
  and _25386_ (_03484_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _25387_ (_03485_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _25388_ (_03486_, _03485_, _03484_);
  or _25389_ (_03487_, _03486_, _03483_);
  and _25390_ (_03488_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _25391_ (_03489_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _25392_ (_03490_, _03489_, _03488_);
  and _25393_ (_03491_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _25394_ (_03492_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _25395_ (_03493_, _03492_, _03491_);
  or _25396_ (_03494_, _03493_, _03490_);
  or _25397_ (_03495_, _03494_, _03487_);
  or _25398_ (_03496_, _03495_, _03480_);
  and _25399_ (_03497_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _25400_ (_03498_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _25401_ (_03499_, _03498_, _03497_);
  and _25402_ (_03500_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not _25403_ (_03501_, _12515_);
  and _25404_ (_03502_, _01368_, _03501_);
  or _25405_ (_03503_, _03502_, _03500_);
  or _25406_ (_03504_, _03503_, _03499_);
  and _25407_ (_03505_, _03162_, _01373_);
  and _25408_ (_03506_, _03125_, _01399_);
  or _25409_ (_03507_, _03506_, _03505_);
  and _25410_ (_03508_, _03367_, _01405_);
  and _25411_ (_03509_, _03201_, _01413_);
  or _25412_ (_03510_, _03509_, _03508_);
  or _25413_ (_03511_, _03510_, _03507_);
  or _25414_ (_03512_, _03511_, _03504_);
  and _25415_ (_03513_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _25416_ (_03514_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _25417_ (_03515_, _03514_, _03513_);
  or _25418_ (_03516_, _03515_, _03512_);
  or _25419_ (_03517_, _03516_, _03496_);
  and _25420_ (_03518_, _03517_, _01441_);
  and _25421_ (_03520_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or _25422_ (_03521_, _03520_, _03518_);
  or _25423_ (_03522_, _03521_, _01287_);
  nand _25424_ (_03524_, _01287_, _07434_);
  and _25425_ (_03525_, _03524_, _05141_);
  and _25426_ (_03716_, _03525_, _03522_);
  and _25427_ (_03526_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _25428_ (_03527_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _25429_ (_03528_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _25430_ (_03529_, _03528_, _03527_);
  and _25431_ (_03530_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _25432_ (_03531_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _25433_ (_03532_, _03531_, _03530_);
  or _25434_ (_03533_, _03532_, _03529_);
  and _25435_ (_03534_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _25436_ (_03535_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _25437_ (_03536_, _03535_, _03534_);
  and _25438_ (_03537_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _25439_ (_03538_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _25440_ (_03539_, _03538_, _03537_);
  or _25441_ (_03540_, _03539_, _03536_);
  or _25442_ (_03541_, _03540_, _03533_);
  and _25443_ (_03542_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _25444_ (_03543_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _25445_ (_03544_, _03543_, _03542_);
  and _25446_ (_03545_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _25447_ (_03546_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _25448_ (_03547_, _03546_, _03545_);
  or _25449_ (_03548_, _03547_, _03544_);
  and _25450_ (_03549_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _25451_ (_03550_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _25452_ (_03551_, _03550_, _03549_);
  and _25453_ (_03552_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _25454_ (_03553_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _25455_ (_03554_, _03553_, _03552_);
  or _25456_ (_03555_, _03554_, _03551_);
  or _25457_ (_03556_, _03555_, _03548_);
  or _25458_ (_03557_, _03556_, _03541_);
  and _25459_ (_03558_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _25460_ (_03559_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _25461_ (_03560_, _03559_, _03558_);
  and _25462_ (_03561_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _25463_ (_03562_, _12569_);
  and _25464_ (_03563_, _01368_, _03562_);
  or _25465_ (_03564_, _03563_, _03561_);
  or _25466_ (_03565_, _03564_, _03560_);
  and _25467_ (_03566_, _03120_, _01399_);
  and _25468_ (_03567_, _03167_, _01373_);
  or _25469_ (_03568_, _03567_, _03566_);
  and _25470_ (_03569_, _03359_, _01405_);
  and _25471_ (_03570_, _03205_, _01413_);
  or _25472_ (_03571_, _03570_, _03569_);
  or _25473_ (_03572_, _03571_, _03568_);
  or _25474_ (_03573_, _03572_, _03565_);
  and _25475_ (_03574_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _25476_ (_03575_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _25477_ (_03576_, _03575_, _03574_);
  or _25478_ (_03577_, _03576_, _03573_);
  or _25479_ (_03578_, _03577_, _03557_);
  and _25480_ (_03579_, _03578_, _01441_);
  or _25481_ (_03580_, _03579_, _01287_);
  or _25482_ (_03581_, _03580_, _03526_);
  nand _25483_ (_03582_, _01287_, _06617_);
  and _25484_ (_03583_, _03582_, _05141_);
  and _25485_ (_03728_, _03583_, _03581_);
  nor _25486_ (_03584_, _01048_, _01047_);
  or _25487_ (_03585_, _03584_, _01049_);
  and _25488_ (_03586_, _01051_, _05141_);
  and _25489_ (_03731_, _03586_, _03585_);
  or _25490_ (_03587_, _02459_, _06004_);
  or _25491_ (_03588_, _06678_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _25492_ (_03589_, _03588_, _05141_);
  and _25493_ (_03745_, _03589_, _03587_);
  not _25494_ (_03590_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _25495_ (_03591_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _25496_ (_03592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25497_ (_03593_, _05626_, _03592_);
  or _25498_ (_03594_, _03593_, _08654_);
  nor _25499_ (_03595_, _03594_, _03591_);
  nand _25500_ (_03596_, _03595_, _03590_);
  nor _25501_ (_03597_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor _25502_ (_03598_, _03597_, _03595_);
  nand _25503_ (_03599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _25504_ (_03600_, _03599_, _03598_);
  and _25505_ (_03602_, _03600_, _05141_);
  and _25506_ (_03777_, _03602_, _03596_);
  and _25507_ (_03604_, _06674_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nand _25508_ (_03605_, _05297_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _25509_ (_03606_, _03605_, _05278_);
  nor _25510_ (_03607_, _02459_, _06062_);
  or _25511_ (_03608_, _03607_, _03606_);
  or _25512_ (_03609_, _03608_, _03604_);
  and _25513_ (_03779_, _03609_, _05141_);
  and _25514_ (_03610_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _25515_ (_03611_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or _25516_ (_03612_, _03611_, _03610_);
  and _25517_ (_03795_, _03612_, _05141_);
  and _25518_ (_03613_, _06293_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _25519_ (_03614_, _06774_, _06560_);
  or _25520_ (_03615_, _03614_, _06990_);
  or _25521_ (_03616_, _12671_, _02778_);
  or _25522_ (_03617_, _03616_, _02862_);
  or _25523_ (_03618_, _03617_, _07107_);
  or _25524_ (_03619_, _03618_, _03615_);
  or _25525_ (_03620_, _03619_, _02855_);
  and _25526_ (_03621_, _03620_, _06296_);
  or _25527_ (_03806_, _03621_, _03613_);
  and _25528_ (_03816_, _03598_, _05141_);
  nor _25529_ (_03624_, _02621_, _08366_);
  and _25530_ (_03625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or _25531_ (_03626_, _03625_, rxd_i);
  or _25532_ (_03627_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _25533_ (_03628_, _03627_, _01801_);
  or _25534_ (_03629_, _03628_, _01789_);
  and _25535_ (_03630_, _03629_, _03626_);
  or _25536_ (_03631_, _03630_, _03624_);
  nand _25537_ (_03632_, _01789_, _02596_);
  and _25538_ (_03633_, _03632_, _06715_);
  and _25539_ (_03635_, _03633_, _03631_);
  and _25540_ (_03636_, _06713_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _25541_ (_03818_, _03636_, _03635_);
  nor _25542_ (_03835_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  nand _25543_ (_03638_, _06707_, _05604_);
  or _25544_ (_03639_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _25545_ (_03640_, _03639_, _05141_);
  and _25546_ (_03849_, _03640_, _03638_);
  or _25547_ (_03641_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nand _25548_ (_03642_, pc_log_change, _02403_);
  and _25549_ (_03644_, _03642_, _05141_);
  and _25550_ (_03854_, _03644_, _03641_);
  and _25551_ (_03645_, _02043_, _06008_);
  nand _25552_ (_03646_, _03645_, _05963_);
  or _25553_ (_03647_, _03645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _25554_ (_03648_, _03647_, _05647_);
  and _25555_ (_03649_, _03648_, _03646_);
  nand _25556_ (_03650_, _02049_, _05960_);
  or _25557_ (_03651_, _02049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _25558_ (_03652_, _03651_, _05925_);
  and _25559_ (_03653_, _03652_, _03650_);
  and _25560_ (_03654_, _00696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _25561_ (_03655_, _03654_, rst);
  or _25562_ (_03656_, _03655_, _03653_);
  or _25563_ (_03856_, _03656_, _03649_);
  or _25564_ (_03657_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand _25565_ (_03658_, _07619_, _06457_);
  and _25566_ (_03659_, _03658_, _05141_);
  and _25567_ (_03871_, _03659_, _03657_);
  and _25568_ (_03660_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _25569_ (_03661_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or _25570_ (_03662_, _03661_, _03660_);
  and _25571_ (_03876_, _03662_, _05141_);
  and _25572_ (_03663_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _25573_ (_03664_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  or _25574_ (_03665_, _03664_, _03663_);
  and _25575_ (_03882_, _03665_, _05141_);
  or _25576_ (_03666_, _07619_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand _25577_ (_03667_, _07619_, _06487_);
  and _25578_ (_03668_, _03667_, _05141_);
  and _25579_ (_03884_, _03668_, _03666_);
  and _25580_ (_03669_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _25581_ (_03670_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or _25582_ (_03671_, _03670_, _03669_);
  and _25583_ (_03886_, _03671_, _05141_);
  and _25584_ (_03672_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _25585_ (_03673_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or _25586_ (_03674_, _03673_, _03672_);
  and _25587_ (_03888_, _03674_, _05141_);
  and _25588_ (_03675_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _25589_ (_03890_, _03675_, _02614_);
  and _25590_ (_03676_, _06696_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _25591_ (_03677_, _03676_, _02594_);
  and _25592_ (_03894_, _03677_, _05141_);
  and _25593_ (_03678_, _01795_, _09587_);
  and _25594_ (_03679_, _03678_, _06697_);
  nand _25595_ (_03680_, _03679_, _02596_);
  or _25596_ (_03681_, _03679_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _25597_ (_03682_, _03681_, _05141_);
  and _25598_ (_03899_, _03682_, _03680_);
  and _25599_ (_03683_, _06715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _25600_ (_03904_, _03683_, _02675_);
  nor _25601_ (_03684_, _08440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor _25602_ (_03685_, _03684_, _02507_);
  and _25603_ (_03686_, _11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _25604_ (_03687_, _03686_, _08457_);
  or _25605_ (_03689_, _03687_, _03685_);
  and _25606_ (_03690_, _03689_, _08464_);
  nand _25607_ (_03691_, _08463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand _25608_ (_03692_, _03691_, _11727_);
  or _25609_ (_03693_, _03692_, _03690_);
  nand _25610_ (_03694_, _08471_, _06178_);
  or _25611_ (_03695_, _11789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _25612_ (_03696_, _03695_, _05141_);
  and _25613_ (_03697_, _03696_, _03694_);
  and _25614_ (_03908_, _03697_, _03693_);
  nand _25615_ (_03699_, _06707_, _06178_);
  or _25616_ (_03701_, _06707_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _25617_ (_03702_, _03701_, _05141_);
  and _25618_ (_03910_, _03702_, _03699_);
  and _25619_ (_03703_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _25620_ (_03704_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or _25621_ (_03705_, _03704_, _03703_);
  and _25622_ (_03912_, _03705_, _05141_);
  and _25623_ (_03706_, _08078_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _25624_ (_03707_, _06244_, _08078_);
  or _25625_ (_03708_, _03707_, _03706_);
  and _25626_ (_03920_, _03708_, _05141_);
  nand _25627_ (_03710_, _00698_, _06875_);
  or _25628_ (_03711_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25629_ (_03712_, _03711_, _05925_);
  and _25630_ (_03714_, _03712_, _03710_);
  nor _25631_ (_03715_, _05646_, _03298_);
  and _25632_ (_03717_, _00690_, _06008_);
  nand _25633_ (_03718_, _03717_, _05963_);
  or _25634_ (_03719_, _03717_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25635_ (_03720_, _03719_, _05647_);
  and _25636_ (_03721_, _03720_, _03718_);
  or _25637_ (_03722_, _03721_, _03715_);
  or _25638_ (_03723_, _03722_, _03714_);
  and _25639_ (_03923_, _03723_, _05141_);
  and _25640_ (_03724_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _25641_ (_03725_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or _25642_ (_03726_, _03725_, _03724_);
  and _25643_ (_03933_, _03726_, _05141_);
  and _25644_ (_03727_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _25645_ (_03729_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25646_ (_03730_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _25647_ (_03732_, _03730_, _03729_);
  and _25648_ (_03733_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _25649_ (_03734_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _25650_ (_03735_, _03734_, _03733_);
  or _25651_ (_03736_, _03735_, _03732_);
  and _25652_ (_03737_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _25653_ (_03738_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _25654_ (_03739_, _03738_, _03737_);
  and _25655_ (_03740_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _25656_ (_03741_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _25657_ (_03742_, _03741_, _03740_);
  or _25658_ (_03743_, _03742_, _03739_);
  or _25659_ (_03744_, _03743_, _03736_);
  and _25660_ (_03746_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _25661_ (_03747_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _25662_ (_03748_, _03747_, _03746_);
  and _25663_ (_03749_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _25664_ (_03750_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _25665_ (_03751_, _03750_, _03749_);
  or _25666_ (_03752_, _03751_, _03748_);
  and _25667_ (_03753_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _25668_ (_03754_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _25669_ (_03755_, _03754_, _03753_);
  and _25670_ (_03756_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _25671_ (_03757_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _25672_ (_03758_, _03757_, _03756_);
  or _25673_ (_03759_, _03758_, _03755_);
  or _25674_ (_03760_, _03759_, _03752_);
  or _25675_ (_03761_, _03760_, _03744_);
  and _25676_ (_03762_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _25677_ (_03763_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _25678_ (_03764_, _03763_, _03762_);
  and _25679_ (_03765_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _25680_ (_03766_, _01368_, _12257_);
  or _25681_ (_03767_, _03766_, _03765_);
  or _25682_ (_03768_, _03767_, _03764_);
  and _25683_ (_03769_, _03099_, _01399_);
  and _25684_ (_03770_, _03140_, _01373_);
  or _25685_ (_03771_, _03770_, _03769_);
  and _25686_ (_03772_, _03336_, _01405_);
  and _25687_ (_03773_, _03227_, _01413_);
  or _25688_ (_03774_, _03773_, _03772_);
  or _25689_ (_03775_, _03774_, _03771_);
  or _25690_ (_03776_, _03775_, _03768_);
  and _25691_ (_03778_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _25692_ (_03780_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _25693_ (_03781_, _03780_, _03778_);
  or _25694_ (_03782_, _03781_, _03776_);
  or _25695_ (_03783_, _03782_, _03761_);
  and _25696_ (_03784_, _03783_, _01441_);
  or _25697_ (_03785_, _03784_, _01287_);
  or _25698_ (_03786_, _03785_, _03727_);
  nand _25699_ (_03787_, _01287_, _07259_);
  and _25700_ (_03788_, _03787_, _05141_);
  and _25701_ (_03979_, _03788_, _03786_);
  and _25702_ (_03789_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _25703_ (_03790_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _25704_ (_03791_, _03790_, _03789_);
  and _25705_ (_03792_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _25706_ (_03793_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _25707_ (_03794_, _03793_, _03792_);
  or _25708_ (_03796_, _03794_, _03791_);
  and _25709_ (_03797_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _25710_ (_03798_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _25711_ (_03799_, _03798_, _03797_);
  and _25712_ (_03800_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _25713_ (_03801_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _25714_ (_03802_, _03801_, _03800_);
  or _25715_ (_03803_, _03802_, _03799_);
  or _25716_ (_03804_, _03803_, _03796_);
  and _25717_ (_03805_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _25718_ (_03807_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _25719_ (_03808_, _03807_, _03805_);
  and _25720_ (_03809_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _25721_ (_03810_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _25722_ (_03811_, _03810_, _03809_);
  or _25723_ (_03812_, _03811_, _03808_);
  and _25724_ (_03813_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _25725_ (_03814_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _25726_ (_03815_, _03814_, _03813_);
  and _25727_ (_03817_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _25728_ (_03819_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or _25729_ (_03820_, _03819_, _03817_);
  or _25730_ (_03821_, _03820_, _03815_);
  or _25731_ (_03822_, _03821_, _03812_);
  or _25732_ (_03823_, _03822_, _03804_);
  and _25733_ (_03824_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _25734_ (_03825_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _25735_ (_03826_, _03825_, _03824_);
  and _25736_ (_03827_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _25737_ (_03828_, _01368_, _12325_);
  or _25738_ (_03829_, _03828_, _03827_);
  or _25739_ (_03830_, _03829_, _03826_);
  and _25740_ (_03831_, _03181_, _01373_);
  and _25741_ (_03832_, _03115_, _01399_);
  or _25742_ (_03833_, _03832_, _03831_);
  and _25743_ (_03834_, _03363_, _01405_);
  and _25744_ (_03836_, _03194_, _01413_);
  or _25745_ (_03837_, _03836_, _03834_);
  or _25746_ (_03838_, _03837_, _03833_);
  or _25747_ (_03839_, _03838_, _03830_);
  and _25748_ (_03840_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _25749_ (_03841_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _25750_ (_03842_, _03841_, _03840_);
  or _25751_ (_03843_, _03842_, _03839_);
  or _25752_ (_03844_, _03843_, _03823_);
  and _25753_ (_03845_, _03844_, _01441_);
  and _25754_ (_03846_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or _25755_ (_03847_, _03846_, _03845_);
  or _25756_ (_03848_, _03847_, _01287_);
  nand _25757_ (_03850_, _01287_, _07350_);
  and _25758_ (_03851_, _03850_, _05141_);
  and _25759_ (_03983_, _03851_, _03848_);
  and _25760_ (_03852_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _25761_ (_03853_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _25762_ (_03855_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _25763_ (_03857_, _03855_, _03853_);
  and _25764_ (_03858_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _25765_ (_03859_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _25766_ (_03860_, _03859_, _03858_);
  or _25767_ (_03861_, _03860_, _03857_);
  and _25768_ (_03862_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _25769_ (_03863_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _25770_ (_03864_, _03863_, _03862_);
  and _25771_ (_03865_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _25772_ (_03866_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _25773_ (_03867_, _03866_, _03865_);
  or _25774_ (_03868_, _03867_, _03864_);
  or _25775_ (_03869_, _03868_, _03861_);
  and _25776_ (_03870_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _25777_ (_03872_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _25778_ (_03873_, _03872_, _03870_);
  and _25779_ (_03874_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _25780_ (_03875_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _25781_ (_03877_, _03875_, _03874_);
  or _25782_ (_03878_, _03877_, _03873_);
  and _25783_ (_03879_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _25784_ (_03880_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _25785_ (_03881_, _03880_, _03879_);
  and _25786_ (_03883_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _25787_ (_03885_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _25788_ (_03887_, _03885_, _03883_);
  or _25789_ (_03889_, _03887_, _03881_);
  or _25790_ (_03891_, _03889_, _03878_);
  or _25791_ (_03892_, _03891_, _03869_);
  and _25792_ (_03893_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _25793_ (_03895_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _25794_ (_03896_, _03895_, _03893_);
  and _25795_ (_03897_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _25796_ (_03898_, _01368_, _12409_);
  or _25797_ (_03900_, _03898_, _03897_);
  or _25798_ (_03901_, _03900_, _03896_);
  and _25799_ (_03902_, _03092_, _01399_);
  and _25800_ (_03903_, _03147_, _01373_);
  or _25801_ (_03905_, _03903_, _03902_);
  and _25802_ (_03906_, _03346_, _01405_);
  and _25803_ (_03907_, _03223_, _01413_);
  or _25804_ (_03909_, _03907_, _03906_);
  or _25805_ (_03911_, _03909_, _03905_);
  or _25806_ (_03913_, _03911_, _03901_);
  and _25807_ (_03914_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _25808_ (_03915_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _25809_ (_03916_, _03915_, _03914_);
  or _25810_ (_03917_, _03916_, _03913_);
  or _25811_ (_03918_, _03917_, _03892_);
  and _25812_ (_03919_, _03918_, _01441_);
  or _25813_ (_03921_, _03919_, _01287_);
  or _25814_ (_03922_, _03921_, _03852_);
  or _25815_ (_03924_, _03439_, _06669_);
  and _25816_ (_03925_, _03924_, _05141_);
  and _25817_ (_03989_, _03925_, _03922_);
  and _25818_ (_03926_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _25819_ (_03927_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _25820_ (_03928_, _03927_, _03926_);
  and _25821_ (_03929_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _25822_ (_03930_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _25823_ (_03931_, _03930_, _03929_);
  or _25824_ (_03932_, _03931_, _03928_);
  and _25825_ (_03934_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _25826_ (_03935_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _25827_ (_03937_, _03935_, _03934_);
  and _25828_ (_03938_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _25829_ (_03939_, _01325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _25830_ (_03940_, _03939_, _03938_);
  or _25831_ (_03941_, _03940_, _03937_);
  or _25832_ (_03942_, _03941_, _03932_);
  and _25833_ (_03943_, _01333_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _25834_ (_03944_, _01330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _25835_ (_03945_, _03944_, _03943_);
  and _25836_ (_03946_, _01336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _25837_ (_03947_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _25838_ (_03948_, _03947_, _03946_);
  or _25839_ (_03949_, _03948_, _03945_);
  and _25840_ (_03950_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _25841_ (_03951_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _25842_ (_03952_, _03951_, _03950_);
  and _25843_ (_03953_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _25844_ (_03954_, _01351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _25845_ (_03955_, _03954_, _03953_);
  or _25846_ (_03956_, _03955_, _03952_);
  or _25847_ (_03957_, _03956_, _03949_);
  or _25848_ (_03958_, _03957_, _03942_);
  and _25849_ (_03959_, _01286_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _25850_ (_03960_, _01359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _25851_ (_03961_, _03960_, _03959_);
  and _25852_ (_03962_, _01365_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not _25853_ (_03963_, _12304_);
  and _25854_ (_03964_, _01368_, _03963_);
  or _25855_ (_03965_, _03964_, _03962_);
  or _25856_ (_03966_, _03965_, _03961_);
  and _25857_ (_03967_, _03103_, _01399_);
  and _25858_ (_03968_, _03153_, _01373_);
  or _25859_ (_03969_, _03968_, _03967_);
  and _25860_ (_03970_, _03341_, _01405_);
  and _25861_ (_03971_, _03219_, _01413_);
  or _25862_ (_03972_, _03971_, _03970_);
  or _25863_ (_03973_, _03972_, _03969_);
  or _25864_ (_03974_, _03973_, _03966_);
  and _25865_ (_03975_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _25866_ (_03976_, _01425_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _25867_ (_03977_, _03976_, _03975_);
  or _25868_ (_03978_, _03977_, _03974_);
  or _25869_ (_03980_, _03978_, _03958_);
  and _25870_ (_03981_, _03980_, _01441_);
  and _25871_ (_03982_, _01474_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or _25872_ (_03984_, _03982_, _03981_);
  or _25873_ (_03985_, _03984_, _01287_);
  nand _25874_ (_03986_, _01287_, _07200_);
  and _25875_ (_03987_, _03986_, _05141_);
  and _25876_ (_03993_, _03987_, _03985_);
  nor _25877_ (_03988_, _05960_, _08078_);
  and _25878_ (_03990_, _08078_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _25879_ (_03991_, _03990_, _03988_);
  and _25880_ (_03995_, _03991_, _05141_);
  and _25881_ (_03992_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _25882_ (_03994_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or _25883_ (_03996_, _03994_, _03992_);
  and _25884_ (_03997_, _03996_, _05141_);
  and _25885_ (_03999_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _25886_ (_04000_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or _25887_ (_04001_, _04000_, _03999_);
  and _25888_ (_03998_, _04001_, _05141_);
  and _25889_ (_04002_, _07619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _25890_ (_04003_, _12951_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or _25891_ (_04004_, _04003_, _04002_);
  and _25892_ (_04059_, _04004_, _05141_);
  and _25893_ (_04005_, _13031_, _05523_);
  and _25894_ (_04006_, _01964_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or _25895_ (_04007_, _04006_, _04005_);
  and _25896_ (_04083_, _04007_, _05141_);
  and _25897_ (_04008_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _25898_ (_04009_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _25899_ (_04010_, pc_log_change, _04009_);
  or _25900_ (_04011_, _04010_, _04008_);
  and _25901_ (_04103_, _04011_, _05141_);
  and _25902_ (_04012_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _25903_ (_04013_, _04012_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _25904_ (_04014_, _04013_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and _25905_ (_04015_, _04014_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _25906_ (_04016_, _04015_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and _25907_ (_04017_, _04016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _25908_ (_04018_, _04017_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _25909_ (_04019_, _04018_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and _25910_ (_04020_, _04019_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _25911_ (_04021_, _04020_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _25912_ (_04022_, _04021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _25913_ (_04023_, _04022_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _25914_ (_04024_, _04022_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _25915_ (_04025_, _04024_, _04023_);
  nor _25916_ (_04026_, _04025_, cy_reg);
  and _25917_ (_04027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _25918_ (_04028_, _04027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  not _25919_ (_04029_, _04028_);
  or _25920_ (_04030_, _04027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25921_ (_04031_, _04030_, _04029_);
  not _25922_ (_04032_, _04031_);
  or _25923_ (_04033_, _04028_, _07607_);
  nand _25924_ (_04034_, _04028_, _07607_);
  and _25925_ (_04035_, _04034_, _04033_);
  nand _25926_ (_04036_, _04035_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _25927_ (_04038_, _04035_, _08192_);
  nand _25928_ (_04039_, _04038_, _04036_);
  nand _25929_ (_04040_, _04039_, _04032_);
  not _25930_ (_04041_, _04035_);
  or _25931_ (_04042_, _04041_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _25932_ (_04043_, _04035_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _25933_ (_04044_, _04043_, _04031_);
  nand _25934_ (_04045_, _04044_, _04042_);
  nand _25935_ (_04046_, _04045_, _04040_);
  nand _25936_ (_04047_, _04046_, _04027_);
  nor _25937_ (_04048_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nand _25938_ (_04049_, _04035_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _25939_ (_04050_, _04035_, _07661_);
  nand _25940_ (_04051_, _04050_, _04049_);
  nand _25941_ (_04052_, _04051_, _04032_);
  or _25942_ (_04053_, _04041_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _25943_ (_04054_, _04035_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _25944_ (_04055_, _04054_, _04031_);
  nand _25945_ (_04056_, _04055_, _04053_);
  nand _25946_ (_04057_, _04056_, _04052_);
  nand _25947_ (_04058_, _04057_, _04048_);
  and _25948_ (_04060_, _04058_, _04047_);
  and _25949_ (_04061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02390_);
  nand _25950_ (_04062_, _04035_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _25951_ (_04063_, _04035_, _07691_);
  and _25952_ (_04064_, _04063_, _04062_);
  or _25953_ (_04065_, _04064_, _04032_);
  or _25954_ (_04066_, _04035_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _25955_ (_04067_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _25956_ (_04068_, _04035_, _04067_);
  and _25957_ (_04069_, _04068_, _04066_);
  nand _25958_ (_04070_, _04069_, _04032_);
  nand _25959_ (_04071_, _04070_, _04065_);
  nand _25960_ (_04072_, _04071_, _04061_);
  and _25961_ (_04073_, _04009_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nand _25962_ (_04074_, _04035_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _25963_ (_04075_, _04035_, _08257_);
  nand _25964_ (_04076_, _04075_, _04074_);
  nand _25965_ (_04077_, _04076_, _04032_);
  or _25966_ (_04078_, _04035_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand _25967_ (_04079_, _04035_, _07652_);
  and _25968_ (_04080_, _04079_, _04031_);
  nand _25969_ (_04081_, _04080_, _04078_);
  nand _25970_ (_04082_, _04081_, _04077_);
  nand _25971_ (_04084_, _04082_, _04073_);
  and _25972_ (_04085_, _04084_, _04072_);
  and _25973_ (_04086_, _04085_, _04060_);
  and _25974_ (_04087_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _25975_ (_04088_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor _25976_ (_04089_, _04088_, _04087_);
  and _25977_ (_04090_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _25978_ (_04091_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _25979_ (_04092_, _04091_, _04090_);
  and _25980_ (_04093_, _04092_, _04089_);
  and _25981_ (_04094_, _04093_, _04032_);
  and _25982_ (_04095_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _25983_ (_04096_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nor _25984_ (_04097_, _04096_, _04095_);
  and _25985_ (_04098_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _25986_ (_04099_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _25987_ (_04100_, _04099_, _04098_);
  and _25988_ (_04101_, _04100_, _04097_);
  and _25989_ (_04102_, _04101_, _04031_);
  or _25990_ (_04104_, _04102_, _04041_);
  nor _25991_ (_04105_, _04104_, _04094_);
  and _25992_ (_04106_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _25993_ (_04107_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor _25994_ (_04108_, _04107_, _04106_);
  and _25995_ (_04109_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _25996_ (_04110_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _25997_ (_04111_, _04110_, _04109_);
  and _25998_ (_04112_, _04111_, _04108_);
  and _25999_ (_04113_, _04112_, _04032_);
  and _26000_ (_04114_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _26001_ (_04115_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor _26002_ (_04116_, _04115_, _04114_);
  and _26003_ (_04117_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _26004_ (_04118_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _26005_ (_04119_, _04118_, _04117_);
  and _26006_ (_04120_, _04119_, _04116_);
  and _26007_ (_04121_, _04120_, _04031_);
  or _26008_ (_04122_, _04121_, _04035_);
  nor _26009_ (_04123_, _04122_, _04113_);
  nor _26010_ (_04124_, _04123_, _04105_);
  nor _26011_ (_04125_, _04124_, _04086_);
  and _26012_ (_04126_, _04125_, _04025_);
  nor _26013_ (_04127_, _04125_, _04025_);
  nor _26014_ (_04128_, _04127_, _04126_);
  not _26015_ (_04129_, _04128_);
  nor _26016_ (_04130_, _04021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _26017_ (_04131_, _04130_, _04022_);
  and _26018_ (_04132_, _04131_, _04125_);
  not _26019_ (_04133_, _04132_);
  nor _26020_ (_04134_, _04020_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _26021_ (_04135_, _04134_, _04021_);
  and _26022_ (_04136_, _04135_, _04125_);
  nor _26023_ (_04137_, _04019_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _26024_ (_04138_, _04137_, _04020_);
  and _26025_ (_04139_, _04138_, _04125_);
  nor _26026_ (_04140_, _04139_, _04136_);
  nor _26027_ (_04142_, _04135_, _04125_);
  nor _26028_ (_04143_, _04142_, _04136_);
  not _26029_ (_04144_, _04143_);
  nor _26030_ (_04145_, _04138_, _04125_);
  nor _26031_ (_04146_, _04145_, _04139_);
  nor _26032_ (_04147_, _04018_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _26033_ (_04148_, _04147_, _04019_);
  and _26034_ (_04149_, _04148_, _04125_);
  nor _26035_ (_04150_, _04017_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _26036_ (_04151_, _04150_, _04018_);
  and _26037_ (_04152_, _04151_, _04125_);
  nor _26038_ (_04153_, _04152_, _04149_);
  nor _26039_ (_04154_, _04148_, _04125_);
  nor _26040_ (_04155_, _04154_, _04149_);
  not _26041_ (_04156_, _04155_);
  nor _26042_ (_04157_, _04016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _26043_ (_04158_, _04157_, _04017_);
  and _26044_ (_04159_, _04158_, _04125_);
  nor _26045_ (_04160_, _04158_, _04125_);
  nor _26046_ (_04161_, _04015_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _26047_ (_04162_, _04161_, _04016_);
  and _26048_ (_04163_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _26049_ (_04164_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _26050_ (_04165_, _04164_, _04163_);
  and _26051_ (_04166_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _26052_ (_04167_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _26053_ (_04168_, _04167_, _04166_);
  and _26054_ (_04169_, _04168_, _04165_);
  nor _26055_ (_04170_, _04169_, _04031_);
  and _26056_ (_04171_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _26057_ (_04172_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _26058_ (_04173_, _04172_, _04171_);
  and _26059_ (_04174_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _26060_ (_04175_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _26061_ (_04176_, _04175_, _04174_);
  and _26062_ (_04177_, _04176_, _04173_);
  nor _26063_ (_04178_, _04177_, _04032_);
  or _26064_ (_04179_, _04178_, _04170_);
  and _26065_ (_04180_, _04179_, _04035_);
  and _26066_ (_04181_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _26067_ (_04182_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _26068_ (_04183_, _04182_, _04181_);
  and _26069_ (_04184_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _26070_ (_04185_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _26071_ (_04186_, _04185_, _04184_);
  and _26072_ (_04187_, _04186_, _04183_);
  and _26073_ (_04188_, _04187_, _04032_);
  and _26074_ (_04189_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _26075_ (_04190_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _26076_ (_04191_, _04190_, _04189_);
  and _26077_ (_04192_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _26078_ (_04193_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _26079_ (_04194_, _04193_, _04192_);
  and _26080_ (_04195_, _04194_, _04191_);
  and _26081_ (_04196_, _04195_, _04031_);
  or _26082_ (_04197_, _04196_, _04035_);
  nor _26083_ (_04198_, _04197_, _04188_);
  nor _26084_ (_04199_, _04198_, _04180_);
  nor _26085_ (_04200_, _04199_, _04086_);
  and _26086_ (_04201_, _04200_, _04162_);
  nor _26087_ (_04202_, _04200_, _04162_);
  nor _26088_ (_04203_, _04202_, _04201_);
  and _26089_ (_04204_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _26090_ (_04205_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _26091_ (_04206_, _04205_, _04204_);
  and _26092_ (_04207_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _26093_ (_04208_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _26094_ (_04209_, _04208_, _04207_);
  and _26095_ (_04210_, _04209_, _04206_);
  nor _26096_ (_04211_, _04210_, _04031_);
  and _26097_ (_04212_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _26098_ (_04213_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _26099_ (_04214_, _04213_, _04212_);
  and _26100_ (_04215_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _26101_ (_04216_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _26102_ (_04217_, _04216_, _04215_);
  and _26103_ (_04218_, _04217_, _04214_);
  nor _26104_ (_04219_, _04218_, _04032_);
  or _26105_ (_04220_, _04219_, _04211_);
  and _26106_ (_04221_, _04220_, _04035_);
  and _26107_ (_04222_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _26108_ (_04223_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _26109_ (_04224_, _04223_, _04222_);
  and _26110_ (_04225_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _26111_ (_04226_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _26112_ (_04227_, _04226_, _04225_);
  and _26113_ (_04228_, _04227_, _04224_);
  nor _26114_ (_04229_, _04228_, _04031_);
  and _26115_ (_04230_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _26116_ (_04231_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _26117_ (_04232_, _04231_, _04230_);
  and _26118_ (_04233_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _26119_ (_04234_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _26120_ (_04235_, _04234_, _04233_);
  and _26121_ (_04236_, _04235_, _04232_);
  nor _26122_ (_04237_, _04236_, _04032_);
  or _26123_ (_04238_, _04237_, _04229_);
  and _26124_ (_04239_, _04238_, _04041_);
  nor _26125_ (_04240_, _04239_, _04221_);
  nor _26126_ (_04241_, _04240_, _04086_);
  nor _26127_ (_04242_, _04014_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _26128_ (_04243_, _04242_, _04015_);
  and _26129_ (_04244_, _04243_, _04241_);
  nor _26130_ (_04245_, _04243_, _04241_);
  nor _26131_ (_04246_, _04245_, _04244_);
  nor _26132_ (_04247_, _04013_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _26133_ (_04248_, _04247_, _04014_);
  and _26134_ (_04249_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _26135_ (_04250_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _26136_ (_04251_, _04250_, _04249_);
  and _26137_ (_04252_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _26138_ (_04253_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _26139_ (_04254_, _04253_, _04252_);
  and _26140_ (_04255_, _04254_, _04251_);
  and _26141_ (_04256_, _04255_, _04032_);
  and _26142_ (_04257_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _26143_ (_04258_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _26144_ (_04259_, _04258_, _04257_);
  and _26145_ (_04260_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _26146_ (_04261_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _26147_ (_04262_, _04261_, _04260_);
  and _26148_ (_04263_, _04262_, _04259_);
  and _26149_ (_04264_, _04263_, _04031_);
  or _26150_ (_04265_, _04264_, _04041_);
  nor _26151_ (_04266_, _04265_, _04256_);
  and _26152_ (_04267_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _26153_ (_04268_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _26154_ (_04269_, _04268_, _04267_);
  and _26155_ (_04270_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _26156_ (_04271_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _26157_ (_04272_, _04271_, _04270_);
  and _26158_ (_04273_, _04272_, _04269_);
  nor _26159_ (_04274_, _04273_, _04031_);
  and _26160_ (_04275_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _26161_ (_04276_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _26162_ (_04277_, _04276_, _04275_);
  and _26163_ (_04278_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _26164_ (_04279_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _26165_ (_04280_, _04279_, _04278_);
  and _26166_ (_04281_, _04280_, _04277_);
  nor _26167_ (_04282_, _04281_, _04032_);
  or _26168_ (_04283_, _04282_, _04274_);
  and _26169_ (_04284_, _04283_, _04041_);
  nor _26170_ (_04285_, _04284_, _04266_);
  nor _26171_ (_04286_, _04285_, _04086_);
  and _26172_ (_04287_, _04286_, _04248_);
  nor _26173_ (_04288_, _04012_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _26174_ (_04289_, _04288_, _04013_);
  and _26175_ (_04290_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _26176_ (_04291_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _26177_ (_04292_, _04291_, _04290_);
  and _26178_ (_04293_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _26179_ (_04294_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _26180_ (_04295_, _04294_, _04293_);
  and _26181_ (_04296_, _04295_, _04292_);
  and _26182_ (_04297_, _04296_, _04032_);
  and _26183_ (_04298_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _26184_ (_04299_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _26185_ (_04300_, _04299_, _04298_);
  and _26186_ (_04301_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _26187_ (_04302_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _26188_ (_04303_, _04302_, _04301_);
  and _26189_ (_04304_, _04303_, _04300_);
  and _26190_ (_04305_, _04304_, _04031_);
  or _26191_ (_04306_, _04305_, _04041_);
  nor _26192_ (_04307_, _04306_, _04297_);
  and _26193_ (_04308_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _26194_ (_04309_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _26195_ (_04310_, _04309_, _04308_);
  and _26196_ (_04311_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _26197_ (_04312_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _26198_ (_04313_, _04312_, _04311_);
  and _26199_ (_04314_, _04313_, _04310_);
  nor _26200_ (_04315_, _04314_, _04031_);
  and _26201_ (_04316_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _26202_ (_04317_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _26203_ (_04318_, _04317_, _04316_);
  and _26204_ (_04319_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _26205_ (_04320_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _26206_ (_04321_, _04320_, _04319_);
  and _26207_ (_04322_, _04321_, _04318_);
  nor _26208_ (_04323_, _04322_, _04032_);
  or _26209_ (_04324_, _04323_, _04315_);
  and _26210_ (_04325_, _04324_, _04041_);
  nor _26211_ (_04326_, _04325_, _04307_);
  nor _26212_ (_04327_, _04326_, _04086_);
  and _26213_ (_04328_, _04327_, _04289_);
  not _26214_ (_04329_, _04328_);
  nor _26215_ (_04330_, _04327_, _04289_);
  and _26216_ (_04331_, _02418_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _26217_ (_04332_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _02390_);
  nor _26218_ (_04333_, _04332_, _04331_);
  not _26219_ (_04334_, _04333_);
  not _26220_ (_04335_, _04086_);
  and _26221_ (_04336_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _26222_ (_04337_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _26223_ (_04338_, _04337_, _04336_);
  and _26224_ (_04339_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _26225_ (_04340_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _26226_ (_04341_, _04340_, _04339_);
  and _26227_ (_04342_, _04341_, _04338_);
  and _26228_ (_04343_, _04342_, _04032_);
  and _26229_ (_04344_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _26230_ (_04345_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _26231_ (_04346_, _04345_, _04344_);
  and _26232_ (_04347_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _26233_ (_04348_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _26234_ (_04349_, _04348_, _04347_);
  and _26235_ (_04350_, _04349_, _04346_);
  nand _26236_ (_04351_, _04350_, _04031_);
  nand _26237_ (_04352_, _04351_, _04041_);
  or _26238_ (_04353_, _04352_, _04343_);
  and _26239_ (_04354_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _26240_ (_04355_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _26241_ (_04356_, _04355_, _04354_);
  and _26242_ (_04357_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _26243_ (_04358_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _26244_ (_04359_, _04358_, _04357_);
  and _26245_ (_04360_, _04359_, _04356_);
  and _26246_ (_04361_, _04360_, _04031_);
  and _26247_ (_04362_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _26248_ (_04363_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _26249_ (_04364_, _04363_, _04362_);
  and _26250_ (_04365_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _26251_ (_04366_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _26252_ (_04367_, _04366_, _04365_);
  and _26253_ (_04368_, _04367_, _04364_);
  nand _26254_ (_04369_, _04368_, _04032_);
  nand _26255_ (_04370_, _04369_, _04035_);
  or _26256_ (_04371_, _04370_, _04361_);
  nand _26257_ (_04372_, _04371_, _04353_);
  and _26258_ (_04373_, _04372_, _04335_);
  nand _26259_ (_04374_, _04373_, _04334_);
  nand _26260_ (_04375_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nand _26261_ (_04376_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _26262_ (_04377_, _04376_, _04375_);
  nand _26263_ (_04378_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nand _26264_ (_04379_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _26265_ (_04380_, _04379_, _04378_);
  and _26266_ (_04381_, _04380_, _04377_);
  nand _26267_ (_04382_, _04381_, _04032_);
  nand _26268_ (_04383_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nand _26269_ (_04384_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _26270_ (_04385_, _04384_, _04383_);
  nand _26271_ (_04386_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nand _26272_ (_04387_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _26273_ (_04388_, _04387_, _04386_);
  and _26274_ (_04389_, _04388_, _04385_);
  nand _26275_ (_04390_, _04389_, _04031_);
  and _26276_ (_04391_, _04390_, _04041_);
  nand _26277_ (_04392_, _04391_, _04382_);
  nand _26278_ (_04393_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nand _26279_ (_04394_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _26280_ (_04395_, _04394_, _04393_);
  nand _26281_ (_04396_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nand _26282_ (_04397_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _26283_ (_04398_, _04397_, _04396_);
  and _26284_ (_04399_, _04398_, _04395_);
  nand _26285_ (_04400_, _04399_, _04032_);
  nand _26286_ (_04401_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nand _26287_ (_04402_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _26288_ (_04403_, _04402_, _04401_);
  nand _26289_ (_04404_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nand _26290_ (_04405_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _26291_ (_04406_, _04405_, _04404_);
  and _26292_ (_04407_, _04406_, _04403_);
  nand _26293_ (_04408_, _04407_, _04031_);
  and _26294_ (_04409_, _04408_, _04035_);
  nand _26295_ (_04410_, _04409_, _04400_);
  nand _26296_ (_04411_, _04410_, _04392_);
  and _26297_ (_04412_, _04411_, _04335_);
  nand _26298_ (_04413_, _04412_, _02390_);
  nand _26299_ (_04414_, _04073_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand _26300_ (_04415_, _04061_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _26301_ (_04416_, _04415_, _04414_);
  and _26302_ (_04417_, _04048_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _26303_ (_04418_, _04027_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _26304_ (_04419_, _04418_, _04417_);
  and _26305_ (_04420_, _04419_, _04416_);
  nand _26306_ (_04421_, _04420_, _04032_);
  nand _26307_ (_04422_, _04073_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand _26308_ (_04423_, _04027_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _26309_ (_04424_, _04423_, _04422_);
  nand _26310_ (_04425_, _04061_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand _26311_ (_04426_, _04048_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _26312_ (_04427_, _04426_, _04425_);
  and _26313_ (_04428_, _04427_, _04424_);
  nand _26314_ (_04429_, _04428_, _04031_);
  and _26315_ (_04430_, _04429_, _04035_);
  nand _26316_ (_04431_, _04430_, _04421_);
  and _26317_ (_04432_, _04061_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _26318_ (_04433_, _04027_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _26319_ (_04434_, _04433_, _04432_);
  and _26320_ (_04435_, _04073_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _26321_ (_04436_, _04048_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _26322_ (_04437_, _04436_, _04435_);
  and _26323_ (_04438_, _04437_, _04434_);
  nand _26324_ (_04439_, _04438_, _04032_);
  nand _26325_ (_04440_, _04073_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nand _26326_ (_04441_, _04048_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _26327_ (_04442_, _04441_, _04440_);
  nand _26328_ (_04443_, _04061_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nand _26329_ (_04444_, _04027_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _26330_ (_04445_, _04444_, _04443_);
  and _26331_ (_04446_, _04445_, _04442_);
  nand _26332_ (_04447_, _04446_, _04031_);
  and _26333_ (_04448_, _04447_, _04041_);
  nand _26334_ (_04449_, _04448_, _04439_);
  and _26335_ (_04450_, _04449_, _04431_);
  or _26336_ (_04451_, _04450_, _04086_);
  or _26337_ (_04452_, _04451_, _04009_);
  or _26338_ (_04453_, _04412_, _02390_);
  nand _26339_ (_04454_, _04453_, _04413_);
  or _26340_ (_04455_, _04454_, _04452_);
  and _26341_ (_04456_, _04455_, _04413_);
  not _26342_ (_04457_, _04456_);
  or _26343_ (_04458_, _04373_, _04334_);
  and _26344_ (_04459_, _04458_, _04374_);
  nand _26345_ (_04460_, _04459_, _04457_);
  and _26346_ (_04461_, _04460_, _04374_);
  or _26347_ (_04462_, _04461_, _04330_);
  nand _26348_ (_04463_, _04462_, _04329_);
  nor _26349_ (_04464_, _04286_, _04248_);
  nor _26350_ (_04465_, _04464_, _04287_);
  and _26351_ (_04466_, _04465_, _04463_);
  or _26352_ (_04467_, _04466_, _04287_);
  and _26353_ (_04468_, _04467_, _04246_);
  or _26354_ (_04469_, _04468_, _04244_);
  and _26355_ (_04470_, _04469_, _04203_);
  nor _26356_ (_04471_, _04470_, _04201_);
  nor _26357_ (_04472_, _04471_, _04160_);
  or _26358_ (_04473_, _04472_, _04159_);
  nor _26359_ (_04474_, _04151_, _04125_);
  nor _26360_ (_04475_, _04474_, _04152_);
  nand _26361_ (_04476_, _04475_, _04473_);
  or _26362_ (_04477_, _04476_, _04156_);
  nand _26363_ (_04478_, _04477_, _04153_);
  nand _26364_ (_04479_, _04478_, _04146_);
  or _26365_ (_04480_, _04479_, _04144_);
  nand _26366_ (_04481_, _04480_, _04140_);
  nor _26367_ (_04482_, _04131_, _04125_);
  nor _26368_ (_04483_, _04482_, _04132_);
  nand _26369_ (_04484_, _04483_, _04481_);
  nand _26370_ (_04485_, _04484_, _04133_);
  nor _26371_ (_04486_, _04485_, _04129_);
  and _26372_ (_04487_, _04485_, _04129_);
  nor _26373_ (_04488_, _04487_, _04486_);
  and _26374_ (_04489_, _04488_, cy_reg);
  nor _26375_ (_04490_, _04489_, _04026_);
  nor _26376_ (_04491_, _04490_, _01810_);
  and _26377_ (_04492_, _04490_, _01810_);
  nor _26378_ (_04493_, _04135_, cy_reg);
  and _26379_ (_04494_, _04478_, _04146_);
  nor _26380_ (_04495_, _04494_, _04139_);
  nand _26381_ (_04496_, _04495_, _04144_);
  or _26382_ (_04497_, _04495_, _04144_);
  nand _26383_ (_04498_, _04497_, _04496_);
  and _26384_ (_04499_, _04498_, cy_reg);
  or _26385_ (_04500_, _04499_, _04493_);
  nor _26386_ (_04501_, _04500_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _26387_ (_04502_, _04500_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not _26388_ (_04503_, cy_reg);
  and _26389_ (_04504_, _04148_, _04503_);
  and _26390_ (_04505_, _04475_, _04473_);
  nor _26391_ (_04506_, _04505_, _04152_);
  nand _26392_ (_04507_, _04506_, _04155_);
  or _26393_ (_04508_, _04506_, _04155_);
  nand _26394_ (_04509_, _04508_, _04507_);
  and _26395_ (_04510_, _04509_, cy_reg);
  nor _26396_ (_04511_, _04510_, _04504_);
  nor _26397_ (_04512_, _04511_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _26398_ (_04513_, _04511_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _26399_ (_04514_, _04151_, _04503_);
  or _26400_ (_04515_, _04475_, _04473_);
  and _26401_ (_04516_, _04515_, _04476_);
  and _26402_ (_04517_, _04516_, cy_reg);
  nor _26403_ (_04518_, _04517_, _04514_);
  nor _26404_ (_04519_, _04518_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _26405_ (_04520_, _04518_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _26406_ (_04521_, _04158_, cy_reg);
  nor _26407_ (_04522_, _04159_, _04160_);
  and _26408_ (_04523_, _04522_, _04471_);
  nor _26409_ (_04524_, _04522_, _04471_);
  nor _26410_ (_04525_, _04524_, _04523_);
  and _26411_ (_04526_, _04525_, cy_reg);
  nor _26412_ (_04527_, _04526_, _04521_);
  nor _26413_ (_04528_, _04527_, _02403_);
  and _26414_ (_04529_, _04527_, _02403_);
  and _26415_ (_04530_, _04162_, _04503_);
  nor _26416_ (_04531_, _04469_, _04203_);
  nor _26417_ (_04532_, _04531_, _04470_);
  and _26418_ (_04533_, _04532_, cy_reg);
  or _26419_ (_04534_, _04533_, _04530_);
  nor _26420_ (_04535_, _04534_, _08551_);
  and _26421_ (_04536_, _04534_, _08551_);
  and _26422_ (_04537_, _04243_, _04503_);
  nor _26423_ (_04538_, _04467_, _04246_);
  nor _26424_ (_04539_, _04538_, _04468_);
  and _26425_ (_04540_, _04539_, cy_reg);
  or _26426_ (_04541_, _04540_, _04537_);
  nor _26427_ (_04542_, _04541_, _01968_);
  and _26428_ (_04543_, _04541_, _01968_);
  and _26429_ (_04544_, _04248_, _04503_);
  nor _26430_ (_04545_, _04465_, _04463_);
  nor _26431_ (_04546_, _04545_, _04466_);
  and _26432_ (_04547_, _04546_, cy_reg);
  or _26433_ (_04548_, _04547_, _04544_);
  nor _26434_ (_04549_, _04548_, _02425_);
  and _26435_ (_04550_, _04548_, _02425_);
  nor _26436_ (_04551_, _04289_, cy_reg);
  nor _26437_ (_04552_, _04330_, _04328_);
  or _26438_ (_04553_, _04552_, _04461_);
  nand _26439_ (_04554_, _04552_, _04461_);
  and _26440_ (_04555_, _04554_, _04553_);
  and _26441_ (_04556_, _04555_, cy_reg);
  or _26442_ (_04557_, _04556_, _04551_);
  nor _26443_ (_04558_, _04557_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _26444_ (_04559_, _04557_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _26445_ (_04560_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _26446_ (_04561_, _04454_, _04452_);
  not _26447_ (_04562_, _04561_);
  and _26448_ (_04563_, _04455_, cy_reg);
  and _26449_ (_04564_, _04563_, _04562_);
  nor _26450_ (_04565_, _04564_, _04560_);
  nor _26451_ (_04566_, _04565_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _26452_ (_04567_, _04451_, _04503_);
  not _26453_ (_04568_, _04567_);
  nor _26454_ (_04569_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _26455_ (_04570_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _26456_ (_04571_, _04570_, _04569_);
  nor _26457_ (_04572_, _04571_, _04568_);
  and _26458_ (_04573_, _04571_, _04568_);
  or _26459_ (_04574_, _04573_, _04572_);
  and _26460_ (_04575_, _04565_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _26461_ (_04576_, _04575_, _04574_);
  or _26462_ (_04577_, _04576_, _04566_);
  nor _26463_ (_04578_, _04333_, cy_reg);
  or _26464_ (_04579_, _04459_, _04457_);
  and _26465_ (_04580_, _04579_, _04460_);
  and _26466_ (_04581_, _04580_, cy_reg);
  nor _26467_ (_04582_, _04581_, _04578_);
  nor _26468_ (_04583_, _04582_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26469_ (_04584_, _04582_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _26470_ (_04585_, _04584_, _04583_);
  or _26471_ (_04586_, _04585_, _04577_);
  or _26472_ (_04587_, _04586_, _04559_);
  or _26473_ (_04588_, _04587_, _04558_);
  or _26474_ (_04589_, _04588_, _04550_);
  or _26475_ (_04590_, _04589_, _04549_);
  or _26476_ (_04591_, _04590_, _04543_);
  or _26477_ (_04592_, _04591_, _04542_);
  or _26478_ (_04593_, _04592_, _04536_);
  or _26479_ (_04594_, _04593_, _04535_);
  or _26480_ (_04595_, _04594_, _04529_);
  or _26481_ (_04596_, _04595_, _04528_);
  or _26482_ (_04597_, _04596_, _04520_);
  or _26483_ (_04598_, _04597_, _04519_);
  or _26484_ (_04599_, _04598_, _04513_);
  or _26485_ (_04600_, _04599_, _04512_);
  and _26486_ (_04601_, _04138_, _04503_);
  or _26487_ (_04602_, _04478_, _04146_);
  and _26488_ (_04603_, _04602_, _04479_);
  and _26489_ (_04604_, _04603_, cy_reg);
  or _26490_ (_04605_, _04604_, _04601_);
  nor _26491_ (_04606_, _04605_, _02399_);
  and _26492_ (_04607_, _04605_, _02399_);
  or _26493_ (_04608_, _04607_, _04606_);
  or _26494_ (_04609_, _04608_, _04600_);
  or _26495_ (_04610_, _04609_, _04502_);
  or _26496_ (_04611_, _04610_, _04501_);
  and _26497_ (_04612_, _04131_, _04503_);
  or _26498_ (_04613_, _04483_, _04481_);
  and _26499_ (_04614_, _04613_, _04484_);
  and _26500_ (_04615_, _04614_, cy_reg);
  or _26501_ (_04616_, _04615_, _04612_);
  nor _26502_ (_04617_, _04616_, _13154_);
  and _26503_ (_04618_, _04616_, _13154_);
  or _26504_ (_04619_, _04618_, _04617_);
  or _26505_ (_04620_, _04619_, _04611_);
  or _26506_ (_04621_, _04620_, _04492_);
  or _26507_ (_04622_, _04621_, _04491_);
  and _26508_ (_04623_, _04023_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _26509_ (_04624_, _04023_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _26510_ (_04625_, _04624_, _04623_);
  and _26511_ (_04626_, _04625_, _04503_);
  or _26512_ (_04627_, _04484_, _04129_);
  and _26513_ (_04628_, _04132_, _13116_);
  nor _26514_ (_04629_, _04628_, _04126_);
  nand _26515_ (_04630_, _04629_, _04627_);
  and _26516_ (_04631_, _04625_, _04125_);
  nor _26517_ (_04632_, _04625_, _04125_);
  nor _26518_ (_04633_, _04632_, _04631_);
  nand _26519_ (_04634_, _04633_, _04630_);
  or _26520_ (_04635_, _04633_, _04630_);
  and _26521_ (_04636_, _04635_, _04634_);
  and _26522_ (_04637_, _04636_, cy_reg);
  nor _26523_ (_04638_, _04637_, _04626_);
  nor _26524_ (_04639_, _04638_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or _26525_ (_04640_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand _26526_ (_04641_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _26527_ (_04642_, _04641_, _04640_);
  or _26528_ (_04643_, _04642_, _04623_);
  nand _26529_ (_04644_, _04642_, _04623_);
  and _26530_ (_04645_, _04644_, _04643_);
  not _26531_ (_04646_, _04645_);
  and _26532_ (_04647_, _04630_, _04125_);
  not _26533_ (_04648_, _04625_);
  nor _26534_ (_04649_, _04630_, _04648_);
  or _26535_ (_04650_, _04632_, _04503_);
  or _26536_ (_04651_, _04650_, _04649_);
  or _26537_ (_04652_, _04651_, _04647_);
  nand _26538_ (_04653_, _04652_, _04646_);
  or _26539_ (_04654_, _04652_, _04646_);
  and _26540_ (_04655_, _04654_, _04653_);
  and _26541_ (_04656_, _04638_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or _26542_ (_04657_, _04656_, _04655_);
  or _26543_ (_04658_, _04657_, _04639_);
  or _26544_ (_04659_, _04658_, _04622_);
  nor _26545_ (_04660_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _26546_ (_04661_, _04660_, _13036_);
  nor _26547_ (_04662_, _04661_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _26548_ (_04663_, _04661_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _26549_ (_04664_, _04663_, _04662_);
  or _26550_ (_04665_, _00677_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _26551_ (_04666_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and _26552_ (_04667_, _04666_, _04665_);
  or _26553_ (_04668_, _04667_, _04664_);
  and _26554_ (_04669_, _04660_, _13036_);
  nor _26555_ (_04670_, _04669_, _04661_);
  not _26556_ (_04671_, _04670_);
  or _26557_ (_04672_, _00677_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _26558_ (_04673_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _26559_ (_04674_, _04673_, _04672_);
  nand _26560_ (_04675_, _04674_, _04664_);
  and _26561_ (_04676_, _04675_, _04671_);
  and _26562_ (_04677_, _04676_, _04668_);
  and _26563_ (_04678_, _04664_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _26564_ (_04679_, _02407_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _26565_ (_04680_, _04679_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _26566_ (_04681_, _04680_, _04678_);
  and _26567_ (_04682_, _04664_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _26568_ (_04683_, _02407_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _26569_ (_04684_, _04683_, _00677_);
  or _26570_ (_04685_, _04684_, _04682_);
  and _26571_ (_04686_, _04685_, _04670_);
  and _26572_ (_04687_, _04686_, _04681_);
  or _26573_ (_04688_, _04687_, _04677_);
  and _26574_ (_04689_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26575_ (_04690_, _04689_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _26576_ (_04691_, _04689_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _26577_ (_04692_, _04691_, _04690_);
  not _26578_ (_04693_, _04692_);
  nor _26579_ (_04694_, _04690_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _26580_ (_04695_, _04690_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _26581_ (_04696_, _04695_, _04694_);
  nand _26582_ (_04697_, _04696_, _07691_);
  or _26583_ (_04698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and _26584_ (_04699_, _04698_, _04697_);
  or _26585_ (_04700_, _04699_, _04693_);
  nor _26586_ (_04701_, _04696_, _04067_);
  and _26587_ (_04702_, _04696_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _26588_ (_04703_, _04702_, _04701_);
  or _26589_ (_04704_, _04703_, _04692_);
  and _26590_ (_04705_, _04704_, _04700_);
  or _26591_ (_04706_, _04705_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26592_ (_04707_, _04696_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _26593_ (_04708_, _04696_, _07686_);
  or _26594_ (_04709_, _04708_, _04707_);
  and _26595_ (_04710_, _04709_, _04693_);
  nand _26596_ (_04711_, _04696_, _07696_);
  or _26597_ (_04712_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and _26598_ (_04713_, _04712_, _04692_);
  and _26599_ (_04714_, _04713_, _04711_);
  or _26600_ (_04715_, _04714_, _00677_);
  or _26601_ (_04716_, _04715_, _04710_);
  and _26602_ (_04717_, _02407_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _26603_ (_04718_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [15]);
  or _26604_ (_04719_, _04718_, _04717_);
  and _26605_ (_04720_, _04719_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _26606_ (_04721_, _02407_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _26607_ (_04722_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and _26608_ (_04723_, _04722_, _13036_);
  and _26609_ (_04724_, _04723_, _04721_);
  or _26610_ (_04725_, _04724_, _04720_);
  and _26611_ (_04726_, _04725_, _04689_);
  and _26612_ (_04727_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _00677_);
  or _26613_ (_04728_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  or _26614_ (_04729_, _02407_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _26615_ (_04730_, _04729_, _04728_);
  or _26616_ (_04731_, _04730_, _13036_);
  or _26617_ (_04732_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _26618_ (_04733_, _02407_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _26619_ (_04734_, _04733_, _04732_);
  or _26620_ (_04735_, _04734_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26621_ (_04736_, _04735_, _04731_);
  and _26622_ (_04737_, _04736_, _04727_);
  or _26623_ (_04738_, _04737_, _04726_);
  and _26624_ (_04739_, _04725_, _00677_);
  and _26625_ (_04740_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26626_ (_04741_, _04740_, _04730_);
  or _26627_ (_04742_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _26628_ (_04743_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _26629_ (_04744_, _02407_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _26630_ (_04745_, _04744_, _04743_);
  and _26631_ (_04746_, _04745_, _04742_);
  or _26632_ (_04747_, _04746_, _04741_);
  or _26633_ (_04748_, _04747_, _04739_);
  and _26634_ (_04749_, _04748_, _04738_);
  and _26635_ (_04750_, _04749_, _04716_);
  and _26636_ (_04751_, _04750_, _04706_);
  and _26637_ (_04752_, _04751_, _04688_);
  and _26638_ (_04753_, _04664_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or _26639_ (_04754_, _04717_, _04671_);
  or _26640_ (_04755_, _04754_, _04753_);
  and _26641_ (_04756_, _04755_, _00677_);
  nand _26642_ (_04757_, _04664_, _08257_);
  or _26643_ (_04758_, _04664_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _26644_ (_04759_, _04758_, _04757_);
  or _26645_ (_04760_, _04759_, _04670_);
  and _26646_ (_04761_, _04760_, _04756_);
  or _26647_ (_04762_, _04761_, _04747_);
  and _26648_ (_04763_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _26649_ (_04764_, _02407_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _26650_ (_04765_, _04764_, _04763_);
  and _26651_ (_04766_, _04765_, _13036_);
  and _26652_ (_04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or _26653_ (_04768_, _04767_, _04679_);
  and _26654_ (_04769_, _04768_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _26655_ (_04770_, _04769_, _04766_);
  and _26656_ (_04771_, _04770_, _00677_);
  nand _26657_ (_04772_, _04696_, _07614_);
  and _26658_ (_04773_, _04728_, _04692_);
  and _26659_ (_04774_, _04773_, _04772_);
  nand _26660_ (_04775_, _04696_, _07661_);
  or _26661_ (_04776_, _04696_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _26662_ (_04777_, _04776_, _04693_);
  and _26663_ (_04778_, _04777_, _04775_);
  or _26664_ (_04779_, _04778_, _04774_);
  and _26665_ (_04780_, _04779_, _04771_);
  not _26666_ (_04781_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand _26667_ (_04782_, _04696_, _04781_);
  or _26668_ (_04783_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _26669_ (_04784_, _04783_, _04692_);
  and _26670_ (_04785_, _04784_, _04782_);
  or _26671_ (_04786_, _04696_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand _26672_ (_04787_, _04696_, _08257_);
  and _26673_ (_04788_, _04787_, _04693_);
  and _26674_ (_04789_, _04788_, _04786_);
  or _26675_ (_04790_, _04789_, _04785_);
  and _26676_ (_04791_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  or _26677_ (_04792_, _04683_, _13036_);
  or _26678_ (_04793_, _04792_, _04791_);
  or _26679_ (_04794_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _26680_ (_04795_, _02407_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _26681_ (_04796_, _04795_, _04794_);
  or _26682_ (_04797_, _04796_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26683_ (_04798_, _04797_, _04793_);
  and _26684_ (_04799_, _04798_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26685_ (_04800_, _04768_, _04740_);
  or _26686_ (_04801_, _02407_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _26687_ (_04802_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _26688_ (_04803_, _04802_, _04743_);
  and _26689_ (_04804_, _04803_, _04801_);
  or _26690_ (_04805_, _04804_, _04800_);
  and _26691_ (_04806_, _04805_, _04799_);
  and _26692_ (_04807_, _04806_, _04790_);
  or _26693_ (_04808_, _04807_, _04780_);
  or _26694_ (_04809_, _04805_, _04798_);
  and _26695_ (_04810_, _04809_, _02411_);
  and _26696_ (_04811_, _04810_, _04808_);
  and _26697_ (_04812_, _04811_, _04762_);
  or _26698_ (_04813_, _04812_, _04752_);
  nor _26699_ (_04814_, _04048_, _02418_);
  and _26700_ (_04815_, _04048_, _02418_);
  nor _26701_ (_04816_, _04815_, _04814_);
  nor _26702_ (_04817_, _04814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _26703_ (_04818_, _04814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _26704_ (_04819_, _04818_, _04817_);
  nand _26705_ (_04820_, _04819_, _07691_);
  or _26706_ (_04821_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and _26707_ (_04822_, _04821_, _04027_);
  and _26708_ (_04823_, _04822_, _04820_);
  nand _26709_ (_04824_, _04819_, _07696_);
  or _26710_ (_04825_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and _26711_ (_04826_, _04825_, _04061_);
  and _26712_ (_04827_, _04826_, _04824_);
  or _26713_ (_04828_, _04827_, _04823_);
  nand _26714_ (_04829_, _04819_, _04781_);
  or _26715_ (_04830_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _26716_ (_04831_, _04830_, _04048_);
  and _26717_ (_04832_, _04831_, _04829_);
  nand _26718_ (_04833_, _04819_, _07614_);
  or _26719_ (_04834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and _26720_ (_04835_, _04834_, _04073_);
  and _26721_ (_04836_, _04835_, _04833_);
  or _26722_ (_04837_, _04836_, _04832_);
  or _26723_ (_04838_, _04837_, _04828_);
  and _26724_ (_04839_, _04838_, _04816_);
  and _26725_ (_04840_, _04819_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _26726_ (_04841_, _04819_, _04067_);
  or _26727_ (_04842_, _04841_, _04840_);
  and _26728_ (_04843_, _04842_, _04027_);
  and _26729_ (_04844_, _04819_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _26730_ (_04845_, _04819_, _07686_);
  or _26731_ (_04846_, _04845_, _04844_);
  and _26732_ (_04847_, _04846_, _04061_);
  or _26733_ (_04848_, _04847_, _04843_);
  and _26734_ (_04849_, _04819_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _26735_ (_04850_, _04819_, _07645_);
  or _26736_ (_04851_, _04850_, _04849_);
  and _26737_ (_04852_, _04851_, _04048_);
  and _26738_ (_04853_, _04819_, \oc8051_symbolic_cxrom1.regvalid [9]);
  not _26739_ (_04854_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _26740_ (_04855_, _04819_, _04854_);
  or _26741_ (_04856_, _04855_, _04853_);
  and _26742_ (_04857_, _04856_, _04073_);
  or _26743_ (_04858_, _04857_, _04852_);
  nor _26744_ (_04859_, _04858_, _04848_);
  nor _26745_ (_04860_, _04859_, _04816_);
  or _26746_ (_04861_, _04860_, _04839_);
  or _26747_ (_04862_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand _26748_ (_04863_, _04862_, _04048_);
  and _26749_ (_04864_, _04863_, _02418_);
  or _26750_ (_04865_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand _26751_ (_04866_, _04865_, _04027_);
  or _26752_ (_04867_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand _26753_ (_04868_, _04867_, _04061_);
  and _26754_ (_04869_, _04868_, _04866_);
  or _26755_ (_04870_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand _26756_ (_04871_, _04870_, _04073_);
  or _26757_ (_04872_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nand _26758_ (_04873_, _04872_, _04048_);
  and _26759_ (_04874_, _04873_, _04871_);
  and _26760_ (_04875_, _04874_, _04869_);
  and _26761_ (_04876_, _04875_, _04864_);
  nand _26762_ (_04877_, _04061_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  or _26763_ (_04878_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nand _26764_ (_04879_, _04878_, _04073_);
  and _26765_ (_04880_, _04879_, _04877_);
  or _26766_ (_04881_, \oc8051_symbolic_cxrom1.regarray[3] [5], \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand _26767_ (_04882_, _04881_, _04027_);
  or _26768_ (_04883_, \oc8051_symbolic_cxrom1.regarray[1] [5], \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand _26769_ (_04884_, _04883_, _04061_);
  and _26770_ (_04885_, _04884_, _04882_);
  and _26771_ (_04886_, _04885_, _04880_);
  nand _26772_ (_04887_, _04073_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  or _26773_ (_04888_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand _26774_ (_04889_, _04888_, _04048_);
  and _26775_ (_04890_, _04889_, _04887_);
  nand _26776_ (_04891_, _04027_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _26777_ (_04892_, _04048_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _26778_ (_04893_, _04892_, _04891_);
  and _26779_ (_04894_, _04893_, _04890_);
  and _26780_ (_04895_, _04894_, _04886_);
  and _26781_ (_04896_, _04048_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _26782_ (_04897_, _04061_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or _26783_ (_04898_, _04897_, _04896_);
  and _26784_ (_04899_, _04073_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _26785_ (_04900_, _04027_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  or _26786_ (_04901_, _04900_, _04899_);
  or _26787_ (_04902_, _04901_, _04898_);
  or _26788_ (_04903_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand _26789_ (_04904_, _04903_, _04073_);
  or _26790_ (_04905_, \oc8051_symbolic_cxrom1.regarray[3] [1], \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand _26791_ (_04906_, _04905_, _04027_);
  or _26792_ (_04907_, \oc8051_symbolic_cxrom1.regarray[1] [1], \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand _26793_ (_04908_, _04907_, _04061_);
  and _26794_ (_04909_, _04908_, _04906_);
  and _26795_ (_04910_, _04909_, _04904_);
  and _26796_ (_04911_, _04910_, _04902_);
  and _26797_ (_04912_, _04911_, _04895_);
  and _26798_ (_04913_, _04912_, _04876_);
  or _26799_ (_04914_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nand _26800_ (_04915_, _04914_, _04073_);
  and _26801_ (_04916_, _04915_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _26802_ (_04917_, \oc8051_symbolic_cxrom1.regarray[7] [5], \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nand _26803_ (_04918_, _04917_, _04027_);
  or _26804_ (_04919_, \oc8051_symbolic_cxrom1.regarray[5] [5], \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nand _26805_ (_04920_, _04919_, _04061_);
  and _26806_ (_04921_, _04920_, _04918_);
  or _26807_ (_04922_, \oc8051_symbolic_cxrom1.regarray[7] [1], \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand _26808_ (_04923_, _04922_, _04027_);
  or _26809_ (_04924_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand _26810_ (_04925_, _04924_, _04073_);
  and _26811_ (_04926_, _04925_, _04923_);
  and _26812_ (_04927_, _04926_, _04921_);
  and _26813_ (_04928_, _04927_, _04916_);
  or _26814_ (_04929_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand _26815_ (_04930_, _04929_, _04048_);
  or _26816_ (_04931_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand _26817_ (_04932_, _04931_, _04073_);
  and _26818_ (_04933_, _04932_, _04930_);
  or _26819_ (_04934_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand _26820_ (_04935_, _04934_, _04027_);
  or _26821_ (_04936_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand _26822_ (_04937_, _04936_, _04061_);
  and _26823_ (_04938_, _04937_, _04935_);
  and _26824_ (_04939_, _04938_, _04933_);
  nand _26825_ (_04940_, _04073_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  or _26826_ (_04941_, \oc8051_symbolic_cxrom1.regarray[5] [1], \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand _26827_ (_04942_, _04941_, _04061_);
  and _26828_ (_04943_, _04942_, _04940_);
  nand _26829_ (_04944_, _04027_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _26830_ (_04945_, _04048_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _26831_ (_04946_, _04945_, _04944_);
  and _26832_ (_04947_, _04946_, _04943_);
  and _26833_ (_04948_, _04947_, _04939_);
  and _26834_ (_04949_, _04061_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _26835_ (_04950_, _04048_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or _26836_ (_04951_, _04950_, _04949_);
  and _26837_ (_04952_, _04027_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _26838_ (_04953_, _04073_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  or _26839_ (_04954_, _04953_, _04952_);
  or _26840_ (_04955_, _04954_, _04951_);
  or _26841_ (_04956_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand _26842_ (_04957_, _04956_, _04048_);
  nand _26843_ (_04958_, _04061_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  or _26844_ (_04959_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nand _26845_ (_04960_, _04959_, _04048_);
  and _26846_ (_04961_, _04960_, _04958_);
  and _26847_ (_04962_, _04961_, _04957_);
  and _26848_ (_04963_, _04962_, _04955_);
  and _26849_ (_04964_, _04963_, _04948_);
  and _26850_ (_04965_, _04964_, _04928_);
  or _26851_ (_04966_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _26852_ (_04967_, _04966_, _04913_);
  nor _26853_ (_04968_, _02383_, first_instr);
  and _26854_ (_04969_, _04968_, _04967_);
  nor _26855_ (_04970_, \oc8051_symbolic_cxrom1.regarray[13] [1], \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _26856_ (_04971_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand _26857_ (_04972_, _04971_, _04970_);
  nand _26858_ (_04973_, _04972_, _04061_);
  nor _26859_ (_04974_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _26860_ (_04975_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand _26861_ (_04976_, _04975_, _04974_);
  nand _26862_ (_04977_, _04976_, _04073_);
  not _26863_ (_04978_, _04027_);
  nor _26864_ (_04979_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _26865_ (_04980_, \oc8051_symbolic_cxrom1.regarray[15] [1], \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _26866_ (_04981_, _04980_, _04979_);
  or _26867_ (_04982_, _04981_, _04978_);
  and _26868_ (_04983_, _04982_, _04977_);
  and _26869_ (_04984_, _04983_, _04973_);
  nand _26870_ (_04985_, _04027_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _26871_ (_04986_, _04048_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _26872_ (_04987_, _04986_, _04985_);
  nand _26873_ (_04988_, _04061_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  or _26874_ (_04989_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nand _26875_ (_04990_, _04989_, _04073_);
  and _26876_ (_04991_, _04990_, _04988_);
  and _26877_ (_04992_, _04991_, _04987_);
  not _26878_ (_04993_, _04048_);
  nor _26879_ (_04994_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _26880_ (_04995_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _26881_ (_04996_, _04995_, _04994_);
  or _26882_ (_04997_, _04996_, _04993_);
  nand _26883_ (_04998_, _04073_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _26884_ (_04999_, _04998_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26885_ (_05000_, _04999_, _04997_);
  and _26886_ (_05001_, _05000_, _04992_);
  and _26887_ (_05002_, _04027_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _26888_ (_05003_, _04073_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or _26889_ (_05004_, _05003_, _05002_);
  and _26890_ (_05005_, _04061_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _26891_ (_05006_, _04048_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or _26892_ (_05007_, _05006_, _05005_);
  or _26893_ (_05008_, _05007_, _05004_);
  or _26894_ (_05009_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nand _26895_ (_05010_, _05009_, _04048_);
  or _26896_ (_05011_, \oc8051_symbolic_cxrom1.regarray[15] [5], \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nand _26897_ (_05012_, _05011_, _04027_);
  or _26898_ (_05013_, \oc8051_symbolic_cxrom1.regarray[13] [5], \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nand _26899_ (_05014_, _05013_, _04061_);
  and _26900_ (_05015_, _05014_, _05012_);
  and _26901_ (_05016_, _05015_, _05010_);
  and _26902_ (_05017_, _05016_, _05008_);
  and _26903_ (_05018_, _05017_, _05001_);
  and _26904_ (_05019_, _05018_, _04984_);
  nor _26905_ (_05020_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _26906_ (_05021_, \oc8051_symbolic_cxrom1.regarray[11] [1], \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _26907_ (_05022_, _05021_, _05020_);
  or _26908_ (_05023_, _05022_, _04978_);
  nor _26909_ (_05024_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _26910_ (_05025_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _26911_ (_05026_, _05025_, _05024_);
  or _26912_ (_05027_, _05026_, _04993_);
  nor _26913_ (_05028_, \oc8051_symbolic_cxrom1.regarray[9] [1], \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _26914_ (_05029_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand _26915_ (_05030_, _05029_, _05028_);
  nand _26916_ (_05031_, _05030_, _04061_);
  and _26917_ (_05032_, _05031_, _05027_);
  and _26918_ (_05033_, _05032_, _05023_);
  or _26919_ (_05034_, \oc8051_symbolic_cxrom1.regarray[9] [5], \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nand _26920_ (_05035_, _05034_, _04061_);
  or _26921_ (_05036_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nand _26922_ (_05037_, _05036_, _04073_);
  and _26923_ (_05038_, _05037_, _05035_);
  nand _26924_ (_05039_, _04073_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nand _26925_ (_05040_, _04073_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _26926_ (_05041_, _05040_, _05039_);
  and _26927_ (_05042_, _05041_, _05038_);
  or _26928_ (_05043_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand _26929_ (_05044_, _05043_, _04073_);
  and _26930_ (_05045_, _05044_, _02418_);
  or _26931_ (_05046_, \oc8051_symbolic_cxrom1.regarray[11] [5], \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nand _26932_ (_05047_, _05046_, _04027_);
  or _26933_ (_05048_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nand _26934_ (_05049_, _05048_, _04048_);
  and _26935_ (_05050_, _05049_, _05047_);
  and _26936_ (_05051_, _05050_, _05045_);
  and _26937_ (_05052_, _05051_, _05042_);
  nand _26938_ (_05053_, _04073_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _26939_ (_05054_, _04061_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _26940_ (_05055_, _05054_, _05053_);
  nand _26941_ (_05056_, _04027_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _26942_ (_05057_, _04048_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _26943_ (_05058_, _05057_, _05056_);
  and _26944_ (_05059_, _05058_, _05055_);
  and _26945_ (_05060_, _04027_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _26946_ (_05061_, _04073_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or _26947_ (_05062_, _05061_, _05060_);
  and _26948_ (_05063_, _04048_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _26949_ (_05064_, _04061_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or _26950_ (_05065_, _05064_, _05063_);
  or _26951_ (_05066_, _05065_, _05062_);
  and _26952_ (_05067_, _05066_, _05059_);
  and _26953_ (_05068_, _05067_, _05052_);
  and _26954_ (_05069_, _05068_, _05033_);
  or _26955_ (_05070_, _05069_, _07607_);
  or _26956_ (_05071_, _05070_, _05019_);
  or _26957_ (_05072_, _07607_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _26958_ (_05073_, _04821_, _05072_);
  or _26959_ (_05074_, _05073_, _02418_);
  or _26960_ (_05075_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _26961_ (_05076_, _07607_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _26962_ (_05077_, _05076_, _05075_);
  or _26963_ (_05078_, _05077_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26964_ (_05079_, _05078_, _05074_);
  and _26965_ (_05080_, _05079_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _26966_ (_05081_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _26967_ (_05082_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _26968_ (_05083_, _07607_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _26969_ (_05084_, _05083_, _05082_);
  and _26970_ (_05085_, _05084_, _05081_);
  or _26971_ (_05086_, _07607_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _26972_ (_05087_, _05086_, _04825_);
  and _26973_ (_05088_, _05087_, _04332_);
  or _26974_ (_05089_, _05088_, _05085_);
  or _26975_ (_05090_, _05089_, _05080_);
  and _26976_ (_05091_, _05079_, _02390_);
  and _26977_ (_05092_, _05087_, _04331_);
  or _26978_ (_05093_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or _26979_ (_05094_, _07607_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _26980_ (_05095_, _05094_, _04012_);
  and _26981_ (_05096_, _05095_, _05093_);
  or _26982_ (_05097_, _05096_, _05092_);
  or _26983_ (_05098_, _05097_, _05091_);
  and _26984_ (_05099_, _05098_, _04009_);
  and _26985_ (_05100_, _05099_, _05090_);
  or _26986_ (_05101_, _07607_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _26987_ (_05102_, _04830_, _05101_);
  or _26988_ (_05103_, _05102_, _02418_);
  or _26989_ (_05104_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or _26990_ (_05105_, _07607_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _26991_ (_05106_, _05105_, _05104_);
  or _26992_ (_05107_, _05106_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26993_ (_05108_, _05107_, _05103_);
  and _26994_ (_05109_, _05108_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _26995_ (_05110_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _26996_ (_05111_, _07607_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _26997_ (_05112_, _05111_, _05110_);
  and _26998_ (_05113_, _05112_, _05081_);
  or _26999_ (_05114_, _07607_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _27000_ (_05115_, _05114_, _04834_);
  and _27001_ (_05116_, _05115_, _04332_);
  or _27002_ (_05117_, _05116_, _05113_);
  or _27003_ (_05118_, _05117_, _05109_);
  and _27004_ (_05119_, _05108_, _02390_);
  and _27005_ (_05120_, _05115_, _04331_);
  or _27006_ (_05121_, _07607_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _27007_ (_05122_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27008_ (_05123_, _05122_, _04012_);
  and _27009_ (_05124_, _05123_, _05121_);
  or _27010_ (_05125_, _05124_, _05120_);
  or _27011_ (_05126_, _05125_, _05119_);
  and _27012_ (_05127_, _05126_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27013_ (_05128_, _05127_, _05118_);
  or _27014_ (_05129_, _05128_, _05100_);
  and _27015_ (_05130_, _05129_, _05071_);
  and _27016_ (_05131_, _05130_, _04969_);
  and _27017_ (_05133_, _05131_, _04861_);
  and _27018_ (_05134_, _05133_, _04335_);
  and _27019_ (_05135_, _05134_, _04813_);
  and _27020_ (property_invalid_jc, _05135_, _04659_);
  or _27021_ (_05136_, pc_log_change_r, _04503_);
  nand _27022_ (_05137_, pc_log_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand _27023_ (_00000_, _05137_, _05136_);
  and _27024_ (_05138_, _02383_, first_instr);
  or _27025_ (_00001_, _05138_, rst);
  dff _27026_ (cy_reg, _00000_, clk);
  dff _27027_ (pc_log_change_r, pc_log_change, clk);
  dff _27028_ (first_instr, _00001_, clk);
  dff _27029_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _08867_, clk);
  dff _27030_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _08870_, clk);
  dff _27031_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _08873_, clk);
  dff _27032_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _08877_, clk);
  dff _27033_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _08879_, clk);
  dff _27034_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _08882_, clk);
  dff _27035_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _08887_, clk);
  dff _27036_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _06058_, clk);
  dff _27037_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _08770_, clk);
  dff _27038_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _08775_, clk);
  dff _27039_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _08777_, clk);
  dff _27040_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _08781_, clk);
  dff _27041_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _08785_, clk);
  dff _27042_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _08788_, clk);
  dff _27043_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _08792_, clk);
  dff _27044_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _08796_, clk);
  dff _27045_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _13483_, clk);
  dff _27046_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _13484_, clk);
  dff _27047_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _13485_, clk);
  dff _27048_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _08679_, clk);
  dff _27049_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _13486_, clk);
  dff _27050_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _13487_, clk);
  dff _27051_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _13488_, clk);
  dff _27052_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _13489_, clk);
  dff _27053_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _13475_, clk);
  dff _27054_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _13476_, clk);
  dff _27055_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _13477_, clk);
  dff _27056_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _13478_, clk);
  dff _27057_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _13479_, clk);
  dff _27058_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _13480_, clk);
  dff _27059_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _13481_, clk);
  dff _27060_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _13482_, clk);
  dff _27061_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _08486_, clk);
  dff _27062_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _08490_, clk);
  dff _27063_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _08493_, clk);
  dff _27064_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _08495_, clk);
  dff _27065_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _08498_, clk);
  dff _27066_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _08502_, clk);
  dff _27067_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _08506_, clk);
  dff _27068_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _08510_, clk);
  dff _27069_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _08400_, clk);
  dff _27070_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _08403_, clk);
  dff _27071_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _08407_, clk);
  dff _27072_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _08410_, clk);
  dff _27073_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _08413_, clk);
  dff _27074_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _08416_, clk);
  dff _27075_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _08419_, clk);
  dff _27076_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _08421_, clk);
  dff _27077_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _08310_, clk);
  dff _27078_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _08314_, clk);
  dff _27079_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _08317_, clk);
  dff _27080_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _08321_, clk);
  dff _27081_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _08325_, clk);
  dff _27082_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _08329_, clk);
  dff _27083_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _08331_, clk);
  dff _27084_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _08335_, clk);
  dff _27085_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _13495_, clk);
  dff _27086_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _08219_, clk);
  dff _27087_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _08224_, clk);
  dff _27088_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _08229_, clk);
  dff _27089_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _08234_, clk);
  dff _27090_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _08236_, clk);
  dff _27091_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _08240_, clk);
  dff _27092_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _08244_, clk);
  dff _27093_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _08120_, clk);
  dff _27094_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _08123_, clk);
  dff _27095_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _13490_, clk);
  dff _27096_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _13491_, clk);
  dff _27097_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _13492_, clk);
  dff _27098_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _13493_, clk);
  dff _27099_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _13494_, clk);
  dff _27100_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _08141_, clk);
  dff _27101_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _08042_, clk);
  dff _27102_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _08045_, clk);
  dff _27103_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _08048_, clk);
  dff _27104_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _08051_, clk);
  dff _27105_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _08053_, clk);
  dff _27106_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _08056_, clk);
  dff _27107_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _08058_, clk);
  dff _27108_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _08060_, clk);
  dff _27109_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _07953_, clk);
  dff _27110_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _07957_, clk);
  dff _27111_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _07961_, clk);
  dff _27112_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _07965_, clk);
  dff _27113_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _07969_, clk);
  dff _27114_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _07971_, clk);
  dff _27115_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _07974_, clk);
  dff _27116_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _07976_, clk);
  dff _27117_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _07553_, clk);
  dff _27118_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _07558_, clk);
  dff _27119_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _07562_, clk);
  dff _27120_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _07565_, clk);
  dff _27121_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _07569_, clk);
  dff _27122_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _07573_, clk);
  dff _27123_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _07575_, clk);
  dff _27124_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _07578_, clk);
  dff _27125_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _07443_, clk);
  dff _27126_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _07449_, clk);
  dff _27127_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _07454_, clk);
  dff _27128_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _07460_, clk);
  dff _27129_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _07465_, clk);
  dff _27130_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _07470_, clk);
  dff _27131_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _07475_, clk);
  dff _27132_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _07477_, clk);
  dff _27133_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _07755_, clk);
  dff _27134_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _07760_, clk);
  dff _27135_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _07762_, clk);
  dff _27136_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _07764_, clk);
  dff _27137_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _07767_, clk);
  dff _27138_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _07770_, clk);
  dff _27139_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _07775_, clk);
  dff _27140_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _07778_, clk);
  dff _27141_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _07655_, clk);
  dff _27142_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _07660_, clk);
  dff _27143_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _07664_, clk);
  dff _27144_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _07667_, clk);
  dff _27145_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _07672_, clk);
  dff _27146_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _07677_, clk);
  dff _27147_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _07682_, clk);
  dff _27148_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _07687_, clk);
  dff _27149_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _07863_, clk);
  dff _27150_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _07866_, clk);
  dff _27151_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _07869_, clk);
  dff _27152_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _07873_, clk);
  dff _27153_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _07876_, clk);
  dff _27154_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _07879_, clk);
  dff _27155_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _07881_, clk);
  dff _27156_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _07885_, clk);
  dff _27157_ (\oc8051_symbolic_cxrom1.regvalid [0], _06079_, clk);
  dff _27158_ (\oc8051_symbolic_cxrom1.regvalid [1], _06108_, clk);
  dff _27159_ (\oc8051_symbolic_cxrom1.regvalid [2], _06149_, clk);
  dff _27160_ (\oc8051_symbolic_cxrom1.regvalid [3], _06196_, clk);
  dff _27161_ (\oc8051_symbolic_cxrom1.regvalid [4], _06252_, clk);
  dff _27162_ (\oc8051_symbolic_cxrom1.regvalid [5], _06294_, clk);
  dff _27163_ (\oc8051_symbolic_cxrom1.regvalid [6], _06359_, clk);
  dff _27164_ (\oc8051_symbolic_cxrom1.regvalid [7], _06435_, clk);
  dff _27165_ (\oc8051_symbolic_cxrom1.regvalid [8], _06513_, clk);
  dff _27166_ (\oc8051_symbolic_cxrom1.regvalid [9], _06609_, clk);
  dff _27167_ (\oc8051_symbolic_cxrom1.regvalid [10], _06704_, clk);
  dff _27168_ (\oc8051_symbolic_cxrom1.regvalid [11], _06794_, clk);
  dff _27169_ (\oc8051_symbolic_cxrom1.regvalid [12], _06887_, clk);
  dff _27170_ (\oc8051_symbolic_cxrom1.regvalid [13], _06971_, clk);
  dff _27171_ (\oc8051_symbolic_cxrom1.regvalid [14], _07082_, clk);
  dff _27172_ (\oc8051_symbolic_cxrom1.regvalid [15], _06029_, clk);
  dff _27173_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _05726_, clk);
  dff _27174_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _05729_, clk);
  dff _27175_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _05732_, clk);
  dff _27176_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _05735_, clk);
  dff _27177_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _05738_, clk);
  dff _27178_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _05741_, clk);
  dff _27179_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _05744_, clk);
  dff _27180_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _05596_, clk);
  dff _27181_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _10940_, clk);
  dff _27182_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _10986_, clk);
  dff _27183_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _12116_, clk);
  dff _27184_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _12113_, clk);
  dff _27185_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _12104_, clk);
  dff _27186_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _05756_, clk);
  dff _27187_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _12082_, clk);
  dff _27188_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _05599_, clk);
  dff _27189_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _05760_, clk);
  dff _27190_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _12791_, clk);
  dff _27191_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _05764_, clk);
  dff _27192_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _05767_, clk);
  dff _27193_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _05770_, clk);
  dff _27194_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _12656_, clk);
  dff _27195_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _12109_, clk);
  dff _27196_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _03035_, clk);
  dff _27197_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _11697_, clk);
  dff _27198_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _11719_, clk);
  dff _27199_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _06984_, clk);
  dff _27200_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _08889_, clk);
  dff _27201_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _05304_, clk);
  dff _27202_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _11658_, clk);
  dff _27203_ (\oc8051_top_1.oc8051_decoder1.state [0], _05369_, clk);
  dff _27204_ (\oc8051_top_1.oc8051_decoder1.state [1], _11638_, clk);
  dff _27205_ (\oc8051_top_1.oc8051_decoder1.op [0], _02768_, clk);
  dff _27206_ (\oc8051_top_1.oc8051_decoder1.op [1], _05558_, clk);
  dff _27207_ (\oc8051_top_1.oc8051_decoder1.op [2], _09689_, clk);
  dff _27208_ (\oc8051_top_1.oc8051_decoder1.op [3], _09833_, clk);
  dff _27209_ (\oc8051_top_1.oc8051_decoder1.op [4], _09859_, clk);
  dff _27210_ (\oc8051_top_1.oc8051_decoder1.op [5], _09855_, clk);
  dff _27211_ (\oc8051_top_1.oc8051_decoder1.op [6], _09862_, clk);
  dff _27212_ (\oc8051_top_1.oc8051_decoder1.op [7], _11677_, clk);
  dff _27213_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _00855_, clk);
  dff _27214_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03039_, clk);
  dff _27215_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _11679_, clk);
  dff _27216_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03080_, clk);
  dff _27217_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05235_, clk);
  dff _27218_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03150_, clk);
  dff _27219_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _03152_, clk);
  dff _27220_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05238_, clk);
  dff _27221_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _03195_, clk);
  dff _27222_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _03198_, clk);
  dff _27223_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05251_, clk);
  dff _27224_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03316_, clk);
  dff _27225_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05340_, clk);
  dff _27226_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _03634_, clk);
  dff _27227_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _03637_, clk);
  dff _27228_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _03698_, clk);
  dff _27229_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _01783_, clk);
  dff _27230_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _03806_, clk);
  dff _27231_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05502_, clk);
  dff _27232_ (\oc8051_top_1.oc8051_decoder1.wr , _05451_, clk);
  dff _27233_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03849_, clk);
  dff _27234_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _03910_, clk);
  dff _27235_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _13174_, clk);
  dff _27236_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _11890_, clk);
  dff _27237_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _05139_, clk);
  dff _27238_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _03936_, clk);
  dff _27239_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _00349_, clk);
  dff _27240_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _02876_, clk);
  dff _27241_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _08473_, clk);
  dff _27242_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _02698_, clk);
  dff _27243_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _02137_, clk);
  dff _27244_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _07122_, clk);
  dff _27245_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _04141_, clk);
  dff _27246_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _01027_, clk);
  dff _27247_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _03049_, clk);
  dff _27248_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _02871_, clk);
  dff _27249_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03622_, clk);
  dff _27250_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _02780_, clk);
  dff _27251_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _05140_, clk);
  dff _27252_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _03779_, clk);
  dff _27253_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _02888_, clk);
  dff _27254_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _03745_, clk);
  dff _27255_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _02194_, clk);
  dff _27256_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _02863_, clk);
  dff _27257_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _06673_, clk);
  dff _27258_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _06443_, clk);
  dff _27259_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _06424_, clk);
  dff _27260_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _06258_, clk);
  dff _27261_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _06405_, clk);
  dff _27262_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _06712_, clk);
  dff _27263_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _03920_, clk);
  dff _27264_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _03995_, clk);
  dff _27265_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _03300_, clk);
  dff _27266_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _08821_, clk);
  dff _27267_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _00486_, clk);
  dff _27268_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _02915_, clk);
  dff _27269_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _00457_, clk);
  dff _27270_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _05468_, clk);
  dff _27271_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _01578_, clk);
  dff _27272_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _02935_, clk);
  dff _27273_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _07680_, clk);
  dff _27274_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _12536_, clk);
  dff _27275_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _03623_, clk);
  dff _27276_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _11360_, clk);
  dff _27277_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _02660_, clk);
  dff _27278_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _07670_, clk);
  dff _27279_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _03372_, clk);
  dff _27280_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _02925_, clk);
  dff _27281_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _13260_, clk);
  dff _27282_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _07247_, clk);
  dff _27283_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _10437_, clk);
  dff _27284_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _01842_, clk);
  dff _27285_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _09109_, clk);
  dff _27286_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _07658_, clk);
  dff _27287_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _01927_, clk);
  dff _27288_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _04083_, clk);
  dff _27289_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _00002_, clk);
  dff _27290_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _01183_, clk);
  dff _27291_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _06783_, clk);
  dff _27292_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _00302_, clk);
  dff _27293_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _12994_, clk);
  dff _27294_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _12316_, clk);
  dff _27295_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _12641_, clk);
  dff _27296_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _12620_, clk);
  dff _27297_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _01890_, clk);
  dff _27298_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _01564_, clk);
  dff _27299_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _01467_, clk);
  dff _27300_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _01451_, clk);
  dff _27301_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _10557_, clk);
  dff _27302_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _02738_, clk);
  dff _27303_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _13067_, clk);
  dff _27304_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _10800_, clk);
  dff _27305_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _02734_, clk);
  dff _27306_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _02771_, clk);
  dff _27307_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _02067_, clk);
  dff _27308_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _03319_, clk);
  dff _27309_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _02730_, clk);
  dff _27310_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _01582_, clk);
  dff _27311_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02103_, clk);
  dff _27312_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _02726_, clk);
  dff _27313_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _02806_, clk);
  dff _27314_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _02701_, clk);
  dff _27315_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _01756_, clk);
  dff _27316_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _02723_, clk);
  dff _27317_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _13030_, clk);
  dff _27318_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _04103_, clk);
  dff _27319_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _02715_, clk);
  dff _27320_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _02760_, clk);
  dff _27321_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _05932_, clk);
  dff _27322_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _03601_, clk);
  dff _27323_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _02713_, clk);
  dff _27324_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _07446_, clk);
  dff _27325_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _03854_, clk);
  dff _27326_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _02710_, clk);
  dff _27327_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _02759_, clk);
  dff _27328_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _02797_, clk);
  dff _27329_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _02804_, clk);
  dff _27330_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _11239_, clk);
  dff _27331_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _11104_, clk);
  dff _27332_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _02705_, clk);
  dff _27333_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _13021_, clk);
  dff _27334_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _11979_, clk);
  dff _27335_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _10750_, clk);
  dff _27336_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _10890_, clk);
  dff _27337_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _01733_, clk);
  dff _27338_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _12623_, clk);
  dff _27339_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _03884_, clk);
  dff _27340_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _01824_, clk);
  dff _27341_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _11995_, clk);
  dff _27342_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _06232_, clk);
  dff _27343_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _08991_, clk);
  dff _27344_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _01626_, clk);
  dff _27345_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _07749_, clk);
  dff _27346_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _02840_, clk);
  dff _27347_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _11987_, clk);
  dff _27348_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _10747_, clk);
  dff _27349_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _03871_, clk);
  dff _27350_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _03888_, clk);
  dff _27351_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _03886_, clk);
  dff _27352_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _03882_, clk);
  dff _27353_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03876_, clk);
  dff _27354_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _12016_, clk);
  dff _27355_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _04059_, clk);
  dff _27356_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _03998_, clk);
  dff _27357_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _03997_, clk);
  dff _27358_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _03933_, clk);
  dff _27359_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _03912_, clk);
  dff _27360_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _12008_, clk);
  dff _27361_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _10742_, clk);
  dff _27362_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _10887_, clk);
  dff _27363_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _10943_, clk);
  dff _27364_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _03795_, clk);
  dff _27365_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03033_, clk);
  dff _27366_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _02832_, clk);
  dff _27367_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _02999_, clk);
  dff _27368_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _03045_, clk);
  dff _27369_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _03021_, clk);
  dff _27370_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _03011_, clk);
  dff _27371_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _03006_, clk);
  dff _27372_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _12076_, clk);
  dff _27373_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _03183_, clk);
  dff _27374_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _10555_, clk);
  dff _27375_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _03031_, clk);
  dff _27376_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _10656_, clk);
  dff _27377_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _10936_, clk);
  dff _27378_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _00706_, clk);
  dff _27379_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _00684_, clk);
  dff _27380_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _00670_, clk);
  dff _27381_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _00660_, clk);
  dff _27382_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _00657_, clk);
  dff _27383_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _12157_, clk);
  dff _27384_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _00826_, clk);
  dff _27385_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _00807_, clk);
  dff _27386_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _00788_, clk);
  dff _27387_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _00778_, clk);
  dff _27388_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _12146_, clk);
  dff _27389_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _10715_, clk);
  dff _27390_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _00387_, clk);
  dff _27391_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _00357_, clk);
  dff _27392_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _10647_, clk);
  dff _27393_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _12218_, clk);
  dff _27394_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _00147_, clk);
  dff _27395_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _00209_, clk);
  dff _27396_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _00172_, clk);
  dff _27397_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _00158_, clk);
  dff _27398_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _12212_, clk);
  dff _27399_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _10698_, clk);
  dff _27400_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _11034_, clk);
  dff _27401_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _11077_, clk);
  dff _27402_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _11068_, clk);
  dff _27403_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _11063_, clk);
  dff _27404_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _12227_, clk);
  dff _27405_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _13411_, clk);
  dff _27406_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _13436_, clk);
  dff _27407_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _13431_, clk);
  dff _27408_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _10640_, clk);
  dff _27409_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _02830_, clk);
  dff _27410_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _10388_, clk);
  dff _27411_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _10340_, clk);
  dff _27412_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _12738_, clk);
  dff _27413_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _12018_, clk);
  dff _27414_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _12013_, clk);
  dff _27415_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _11993_, clk);
  dff _27416_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _11975_, clk);
  dff _27417_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _11968_, clk);
  dff _27418_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _12734_, clk);
  dff _27419_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _10382_, clk);
  dff _27420_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _11632_, clk);
  dff _27421_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _11616_, clk);
  dff _27422_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _10377_, clk);
  dff _27423_ (\oc8051_top_1.oc8051_memory_interface1.reti , _10510_, clk);
  dff _27424_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11346_, clk);
  dff _27425_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _11335_, clk);
  dff _27426_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _11323_, clk);
  dff _27427_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _11319_, clk);
  dff _27428_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _12661_, clk);
  dff _27429_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _12648_, clk);
  dff _27430_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _12767_, clk);
  dff _27431_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _10503_, clk);
  dff _27432_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _10494_, clk);
  dff _27433_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _10476_, clk);
  dff _27434_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _11229_, clk);
  dff _27435_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _11523_, clk);
  dff _27436_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _11515_, clk);
  dff _27437_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _10458_, clk);
  dff _27438_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _11645_, clk);
  dff _27439_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _11641_, clk);
  dff _27440_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _11107_, clk);
  dff _27441_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _11221_, clk);
  dff _27442_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11263_, clk);
  dff _27443_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _11666_, clk);
  dff _27444_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _11664_, clk);
  dff _27445_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _11100_, clk);
  dff _27446_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _11675_, clk);
  dff _27447_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _11670_, clk);
  dff _27448_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _11098_, clk);
  dff _27449_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _11217_, clk);
  dff _27450_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _11688_, clk);
  dff _27451_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _11682_, clk);
  dff _27452_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _11703_, clk);
  dff _27453_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _11695_, clk);
  dff _27454_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _11094_, clk);
  dff _27455_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _11214_, clk);
  dff _27456_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _11259_, clk);
  dff _27457_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _11310_, clk);
  dff _27458_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11389_, clk);
  dff _27459_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _11376_, clk);
  dff _27460_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _11163_, clk);
  dff _27461_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11416_, clk);
  dff _27462_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _11409_, clk);
  dff _27463_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _11161_, clk);
  dff _27464_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11236_, clk);
  dff _27465_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _11363_, clk);
  dff _27466_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _11356_, clk);
  dff _27467_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _11166_, clk);
  dff _27468_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _11281_, clk);
  dff _27469_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _02828_, clk);
  dff _27470_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _10251_, clk);
  dff _27471_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _10245_, clk);
  dff _27472_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03037_, clk);
  dff _27473_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _11921_, clk);
  dff _27474_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _11030_, clk);
  dff _27475_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _11300_, clk);
  dff _27476_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _11947_, clk);
  dff _27477_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _10319_, clk);
  dff _27478_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _27479_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _27480_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _27481_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _27482_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _27483_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _27484_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _27485_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _27486_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _27487_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _27488_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _27489_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _27490_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _27491_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _27492_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _27493_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _27494_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _27495_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _27496_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _27497_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _27498_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _27499_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _27500_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _27501_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _27502_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _27503_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _27504_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _27505_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _27506_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _27507_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _27508_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _27509_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _27510_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _00911_, clk);
  dff _27511_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _03835_, clk);
  dff _27512_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _03700_, clk);
  dff _27513_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _03731_, clk);
  dff _27514_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _00666_, clk);
  dff _27515_ (\oc8051_top_1.oc8051_sfr1.bit_out , _03643_, clk);
  dff _27516_ (\oc8051_top_1.oc8051_sfr1.wait_data , _03709_, clk);
  dff _27517_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _03688_, clk);
  dff _27518_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _03716_, clk);
  dff _27519_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _03728_, clk);
  dff _27520_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _03983_, clk);
  dff _27521_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _03979_, clk);
  dff _27522_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _03993_, clk);
  dff _27523_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03989_, clk);
  dff _27524_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _01025_, clk);
  dff _27525_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _12630_, clk);
  dff _27526_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _07160_, clk);
  dff _27527_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _06507_, clk);
  dff _27528_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _03193_, clk);
  dff _27529_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _07061_, clk);
  dff _27530_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _03305_, clk);
  dff _27531_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _03180_, clk);
  dff _27532_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _06503_, clk);
  dff _27533_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _05329_, clk);
  dff _27534_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _13367_, clk);
  dff _27535_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _13352_, clk);
  dff _27536_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _02397_, clk);
  dff _27537_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _13387_, clk);
  dff _27538_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _13380_, clk);
  dff _27539_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _02394_, clk);
  dff _27540_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _13332_, clk);
  dff _27541_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03923_, clk);
  dff _27542_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _05720_, clk);
  dff _27543_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _05717_, clk);
  dff _27544_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _05714_, clk);
  dff _27545_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05707_, clk);
  dff _27546_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _05690_, clk);
  dff _27547_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05687_, clk);
  dff _27548_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _05698_, clk);
  dff _27549_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _02221_, clk);
  dff _27550_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _05790_, clk);
  dff _27551_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _05783_, clk);
  dff _27552_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _01188_, clk);
  dff _27553_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _10236_, clk);
  dff _27554_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _05793_, clk);
  dff _27555_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _05780_, clk);
  dff _27556_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _01207_, clk);
  dff _27557_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _01651_, clk);
  dff _27558_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _09119_, clk);
  dff _27559_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _01389_, clk);
  dff _27560_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _01479_, clk);
  dff _27561_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _01473_, clk);
  dff _27562_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00980_, clk);
  dff _27563_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _01500_, clk);
  dff _27564_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _01484_, clk);
  dff _27565_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00978_, clk);
  dff _27566_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _03087_, clk);
  dff _27567_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _01503_, clk);
  dff _27568_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _07816_, clk);
  dff _27569_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _10115_, clk);
  dff _27570_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _01392_, clk);
  dff _27571_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _01459_, clk);
  dff _27572_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _10191_, clk);
  dff _27573_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _01516_, clk);
  dff _27574_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _01511_, clk);
  dff _27575_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _07981_, clk);
  dff _27576_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _01523_, clk);
  dff _27577_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _01540_, clk);
  dff _27578_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _07616_, clk);
  dff _27579_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _08859_, clk);
  dff _27580_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _07277_, clk);
  dff _27581_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _07206_, clk);
  dff _27582_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _01005_, clk);
  dff _27583_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _01395_, clk);
  dff _27584_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _01465_, clk);
  dff _27585_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _10153_, clk);
  dff _27586_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _01545_, clk);
  dff _27587_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _01543_, clk);
  dff _27588_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00899_, clk);
  dff _27589_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _01553_, clk);
  dff _27590_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _01548_, clk);
  dff _27591_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00890_, clk);
  dff _27592_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _01032_, clk);
  dff _27593_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _10239_, clk);
  dff _27594_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _01758_, clk);
  dff _27595_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _01585_, clk);
  dff _27596_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00863_, clk);
  dff _27597_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _01764_, clk);
  dff _27598_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _01762_, clk);
  dff _27599_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00853_, clk);
  dff _27600_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _01030_, clk);
  dff _27601_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _07297_, clk);
  dff _27602_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02504_, clk);
  dff _27603_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02658_, clk);
  dff _27604_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _02526_, clk);
  dff _27605_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02502_, clk);
  dff _27606_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _02664_, clk);
  dff _27607_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02529_, clk);
  dff _27608_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _02661_, clk);
  dff _27609_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _02824_, clk);
  dff _27610_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02635_, clk);
  dff _27611_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _02523_, clk);
  dff _27612_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02499_, clk);
  dff _27613_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _02670_, clk);
  dff _27614_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _02525_, clk);
  dff _27615_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _02668_, clk);
  dff _27616_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02522_, clk);
  dff _27617_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _03856_, clk);
  dff _27618_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _02501_, clk);
  dff _27619_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02666_, clk);
  dff _27620_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _02634_, clk);
  dff _27621_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _02615_, clk);
  dff _27622_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _02613_, clk);
  dff _27623_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02519_, clk);
  dff _27624_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _02495_, clk);
  dff _27625_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _00987_, clk);
  dff _27626_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02493_, clk);
  dff _27627_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02672_, clk);
  dff _27628_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _02640_, clk);
  dff _27629_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02638_, clk);
  dff _27630_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _02679_, clk);
  dff _27631_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02517_, clk);
  dff _27632_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _02677_, clk);
  dff _27633_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _03119_, clk);
  dff _27634_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _09173_, clk);
  dff _27635_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _09170_, clk);
  dff _27636_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _01779_, clk);
  dff _27637_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _09564_, clk);
  dff _27638_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _09572_, clk);
  dff _27639_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _09569_, clk);
  dff _27640_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _03139_, clk);
  dff _27641_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _02431_, clk);
  dff _27642_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _12861_, clk);
  dff _27643_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _12858_, clk);
  dff _27644_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _12856_, clk);
  dff _27645_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _12854_, clk);
  dff _27646_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _02429_, clk);
  dff _27647_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _12788_, clk);
  dff _27648_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _13205_, clk);
  dff _27649_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _13207_, clk);
  dff _27650_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00366_, clk);
  dff _27651_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00370_, clk);
  dff _27652_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _12090_, clk);
  dff _27653_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _12098_, clk);
  dff _27654_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _12102_, clk);
  dff _27655_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _12073_, clk);
  dff _27656_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _12070_, clk);
  dff _27657_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _12067_, clk);
  dff _27658_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _12080_, clk);
  dff _27659_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _00379_, clk);
  dff _27660_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _12125_, clk);
  dff _27661_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _12119_, clk);
  dff _27662_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _12122_, clk);
  dff _27663_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _12143_, clk);
  dff _27664_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _12134_, clk);
  dff _27665_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _12140_, clk);
  dff _27666_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _12137_, clk);
  dff _27667_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _00374_, clk);
  dff _27668_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _00377_, clk);
  dff _27669_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _00376_, clk);
  dff _27670_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12160_, clk);
  dff _27671_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12154_, clk);
  dff _27672_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12180_, clk);
  dff _27673_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _12190_, clk);
  dff _27674_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12187_, clk);
  dff _27675_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _12246_, clk);
  dff _27676_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _12242_, clk);
  dff _27677_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _00341_, clk);
  dff _27678_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12328_, clk);
  dff _27679_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12324_, clk);
  dff _27680_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _12295_, clk);
  dff _27681_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _12298_, clk);
  dff _27682_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _12307_, clk);
  dff _27683_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _12311_, clk);
  dff _27684_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _12284_, clk);
  dff _27685_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _00345_, clk);
  dff _27686_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _00343_, clk);
  dff _27687_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12334_, clk);
  dff _27688_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12337_, clk);
  dff _27689_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _12348_, clk);
  dff _27690_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _12342_, clk);
  dff _27691_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _12345_, clk);
  dff _27692_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _12360_, clk);
  dff _27693_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _12353_, clk);
  dff _27694_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _00355_, clk);
  dff _27695_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01883_, clk);
  dff _27696_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01921_, clk);
  dff _27697_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01917_, clk);
  dff _27698_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01888_, clk);
  dff _27699_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _11180_, clk);
  dff _27700_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _05132_, clk);
  dff _27701_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _12210_, clk);
  dff _27702_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _12206_, clk);
  dff _27703_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _12203_, clk);
  dff _27704_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _12198_, clk);
  dff _27705_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _06991_, clk);
  dff _27706_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01886_, clk);
  dff _27707_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _12183_, clk);
  dff _27708_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _12163_, clk);
  dff _27709_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _12128_, clk);
  dff _27710_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _07075_, clk);
  dff _27711_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _01149_, clk);
  dff _27712_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _12058_, clk);
  dff _27713_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _07095_, clk);
  dff _27714_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01853_, clk);
  dff _27715_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01874_, clk);
  dff _27716_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _07098_, clk);
  dff _27717_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _03908_, clk);
  dff _27718_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _03017_, clk);
  dff _27719_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _10570_, clk);
  dff _27720_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _10610_, clk);
  dff _27721_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _10583_, clk);
  dff _27722_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _10575_, clk);
  dff _27723_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01871_, clk);
  dff _27724_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _10461_, clk);
  dff _27725_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _10499_, clk);
  dff _27726_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _10492_, clk);
  dff _27727_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _10489_, clk);
  dff _27728_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _11254_, clk);
  dff _27729_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _10529_, clk);
  dff _27730_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _10540_, clk);
  dff _27731_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01868_, clk);
  dff _27732_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01863_, clk);
  dff _27733_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _10347_, clk);
  dff _27734_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _10344_, clk);
  dff _27735_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _12002_, clk);
  dff _27736_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _10417_, clk);
  dff _27737_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _10412_, clk);
  dff _27738_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _10409_, clk);
  dff _27739_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _10406_, clk);
  dff _27740_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01860_, clk);
  dff _27741_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _03178_, clk);
  dff _27742_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _03175_, clk);
  dff _27743_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _03172_, clk);
  dff _27744_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _03170_, clk);
  dff _27745_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _03168_, clk);
  dff _27746_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _03143_, clk);
  dff _27747_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _03141_, clk);
  dff _27748_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _03136_, clk);
  dff _27749_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _03134_, clk);
  dff _27750_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _03132_, clk);
  dff _27751_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _03123_, clk);
  dff _27752_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _03818_, clk);
  dff _27753_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _07457_, clk);
  dff _27754_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _07493_, clk);
  dff _27755_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _10072_, clk);
  dff _27756_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _02973_, clk);
  dff _27757_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _01681_, clk);
  dff _27758_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _06960_, clk);
  dff _27759_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _03090_, clk);
  dff _27760_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _03899_, clk);
  dff _27761_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _08477_, clk);
  dff _27762_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _08312_, clk);
  dff _27763_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _03603_, clk);
  dff _27764_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _03894_, clk);
  dff _27765_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _09143_, clk);
  dff _27766_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _04037_, clk);
  dff _27767_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _03904_, clk);
  dff _27768_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _03098_, clk);
  dff _27769_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _03074_, clk);
  dff _27770_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _02987_, clk);
  dff _27771_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _02897_, clk);
  dff _27772_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _03890_, clk);
  dff _27773_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _03816_, clk);
  dff _27774_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _03777_, clk);
  dff _27775_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _03713_, clk);
  dff _27776_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _03523_, clk);
  dff _27777_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _06717_, clk);
  dff _27778_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _06903_, clk);
  dff _27779_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _06817_, clk);
  dff _27780_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _03519_, clk);
  dff _27781_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _08210_, clk);
  dff _27782_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _07165_, clk);
  dff _27783_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _07038_, clk);
  dff _27784_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _08682_, clk);
  dff _27785_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _08517_, clk);
  dff _27786_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _10068_, clk);
  dff _27787_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _08691_, clk);
  dff _27788_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _10792_, clk);
  dff _27789_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _10718_, clk);
  dff _27790_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _10871_, clk);
  dff _27791_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _03160_, clk);
  dff _27792_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _06966_, clk);
  dff _27793_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _11700_, clk);
  dff _27794_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _11526_, clk);
  dff _27795_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _12085_, clk);
  dff _27796_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _11717_, clk);
  dff _27797_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _06962_, clk);
  dff _27798_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _12406_, clk);
  dff _27799_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _03126_, clk);
  dff _27800_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _07027_, clk);
  dff _27801_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _12815_, clk);
  dff _27802_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _12722_, clk);
  dff _27803_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _06957_, clk);
  dff _27804_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _13390_, clk);
  dff _27805_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _12925_, clk);
  dff _27806_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _07024_, clk);
  dff _27807_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _03067_, clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [8], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [9], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [10], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [11], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [12], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [13], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [14], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [15], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [16], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [0], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [1], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [2], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [3], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [4], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [5], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [6], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [7], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [0], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [1], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [2], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [3], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [4], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [5], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [6], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [7], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.mulOv , ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [0], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [1], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [2], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [3], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [4], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [5], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [6], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [7], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_alu1.divOv , ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.ABINPUT000 [0], ABINPUT000[0]);
  buf(\oc8051_top_1.ABINPUT000 [1], ABINPUT000[1]);
  buf(\oc8051_top_1.ABINPUT000 [2], ABINPUT000[2]);
  buf(\oc8051_top_1.ABINPUT000 [3], ABINPUT000[3]);
  buf(\oc8051_top_1.ABINPUT000 [4], ABINPUT000[4]);
  buf(\oc8051_top_1.ABINPUT000 [5], ABINPUT000[5]);
  buf(\oc8051_top_1.ABINPUT000 [6], ABINPUT000[6]);
  buf(\oc8051_top_1.ABINPUT000 [7], ABINPUT000[7]);
  buf(\oc8051_top_1.ABINPUT000 [8], ABINPUT000[8]);
  buf(\oc8051_top_1.ABINPUT000 [9], ABINPUT000[9]);
  buf(\oc8051_top_1.ABINPUT000 [10], ABINPUT000[10]);
  buf(\oc8051_top_1.ABINPUT000 [11], ABINPUT000[11]);
  buf(\oc8051_top_1.ABINPUT000 [12], ABINPUT000[12]);
  buf(\oc8051_top_1.ABINPUT000 [13], ABINPUT000[13]);
  buf(\oc8051_top_1.ABINPUT000 [14], ABINPUT000[14]);
  buf(\oc8051_top_1.ABINPUT000 [15], ABINPUT000[15]);
  buf(\oc8051_top_1.ABINPUT000 [16], ABINPUT000[16]);
  buf(\oc8051_top_1.ABINPUT000000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.ABINPUT000000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.ABINPUT000000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.ABINPUT000000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.ABINPUT000000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.ABINPUT000000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.ABINPUT000000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.ABINPUT000000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.ABINPUT000000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.ABINPUT000000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.ABINPUT000000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.ABINPUT000000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.ABINPUT000000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.ABINPUT000000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.ABINPUT000000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.ABINPUT000000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.ABINPUT000000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
